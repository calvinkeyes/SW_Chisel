module SWCell(
  input  [1:0]  io_q,
  input  [1:0]  io_r,
  input  [15:0] io_e_i,
  input  [15:0] io_f_i,
  input  [15:0] io_ve_i,
  input  [15:0] io_vf_i,
  input  [15:0] io_vv_i,
  output [15:0] io_e_o,
  output [15:0] io_f_o,
  output [15:0] io_v_o
);
  wire [15:0] _T_2 = $signed(io_ve_i) - 16'sh2; // @[SWChisel.scala 78:17]
  wire [15:0] _T_5 = $signed(io_e_i) - 16'sh1; // @[SWChisel.scala 78:39]
  wire [15:0] e_max = $signed(_T_2) >= $signed(_T_5) ? $signed(_T_2) : $signed(_T_5); // @[SWChisel.scala 78:51 79:11 81:11]
  wire [15:0] _T_9 = $signed(io_vf_i) - 16'sh2; // @[SWChisel.scala 85:17]
  wire [15:0] _T_12 = $signed(io_f_i) - 16'sh1; // @[SWChisel.scala 85:38]
  wire [15:0] f_max = $signed(_T_9) > $signed(_T_12) ? $signed(_T_9) : $signed(_T_12); // @[SWChisel.scala 85:50 86:11 88:11]
  wire [15:0] ef_temp = $signed(e_max) > $signed(f_max) ? $signed(e_max) : $signed(f_max); // @[SWChisel.scala 92:24 93:13 95:13]
  wire [15:0] _v_temp_T_2 = $signed(io_vv_i) + 16'sh2; // @[SWChisel.scala 100:23]
  wire [15:0] _v_temp_T_5 = $signed(io_vv_i) - 16'sh2; // @[SWChisel.scala 102:23]
  wire [15:0] v_temp = io_q == io_r ? $signed(_v_temp_T_2) : $signed(_v_temp_T_5); // @[SWChisel.scala 100:12 102:12 99:24]
  assign io_e_o = $signed(_T_2) >= $signed(_T_5) ? $signed(_T_2) : $signed(_T_5); // @[SWChisel.scala 78:51 79:11 81:11]
  assign io_f_o = $signed(_T_9) > $signed(_T_12) ? $signed(_T_9) : $signed(_T_12); // @[SWChisel.scala 85:50 86:11 88:11]
  assign io_v_o = $signed(v_temp) > $signed(ef_temp) ? $signed(v_temp) : $signed(ef_temp); // @[SWChisel.scala 106:27 107:11 109:11]
endmodule
module MyCounter(
  input        clock,
  input        reset,
  input        io_en,
  output [8:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] _io_out_T_2 = io_out + 9'h1; // @[SWChisel.scala 155:55]
  reg [8:0] io_out_r; // @[Reg.scala 35:20]
  assign io_out = io_out_r; // @[SWChisel.scala 155:12]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      io_out_r <= 9'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_out < 9'h12c) begin // @[SWChisel.scala 155:28]
        io_out_r <= _io_out_T_2;
      end else begin
        io_out_r <= 9'h0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_out_r = _RAND_0[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MAX(
  input         clock,
  input         reset,
  input         io_start,
  input  [15:0] io_in,
  output        io_done,
  output [15:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] max; // @[SWChisel.scala 122:20]
  reg [8:0] counter; // @[SWChisel.scala 133:24]
  wire [8:0] _counter_T_1 = counter - 9'h1; // @[SWChisel.scala 135:24]
  assign io_done = counter == 9'h0; // @[SWChisel.scala 141:17]
  assign io_out = max; // @[SWChisel.scala 123:10]
  always @(posedge clock) begin
    if (reset) begin // @[SWChisel.scala 122:20]
      max <= 16'sh8000; // @[SWChisel.scala 122:20]
    end else if ($signed(io_in) > $signed(max)) begin // @[SWChisel.scala 126:22]
      max <= io_in; // @[SWChisel.scala 127:9]
    end
    if (reset) begin // @[SWChisel.scala 133:24]
      counter <= 9'h12d; // @[SWChisel.scala 133:24]
    end else if (counter == 9'h0) begin // @[SWChisel.scala 141:26]
      counter <= 9'h0; // @[SWChisel.scala 143:13]
    end else if (io_start) begin // @[SWChisel.scala 134:19]
      counter <= _counter_T_1; // @[SWChisel.scala 135:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  max = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  counter = _RAND_1[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SW(
  input         clock,
  input         reset,
  input  [1:0]  io_q_0_b,
  input  [1:0]  io_q_1_b,
  input  [1:0]  io_q_2_b,
  input  [1:0]  io_q_3_b,
  input  [1:0]  io_q_4_b,
  input  [1:0]  io_q_5_b,
  input  [1:0]  io_q_6_b,
  input  [1:0]  io_q_7_b,
  input  [1:0]  io_q_8_b,
  input  [1:0]  io_q_9_b,
  input  [1:0]  io_q_10_b,
  input  [1:0]  io_q_11_b,
  input  [1:0]  io_q_12_b,
  input  [1:0]  io_q_13_b,
  input  [1:0]  io_q_14_b,
  input  [1:0]  io_q_15_b,
  input  [1:0]  io_q_16_b,
  input  [1:0]  io_q_17_b,
  input  [1:0]  io_q_18_b,
  input  [1:0]  io_q_19_b,
  input  [1:0]  io_q_20_b,
  input  [1:0]  io_q_21_b,
  input  [1:0]  io_q_22_b,
  input  [1:0]  io_q_23_b,
  input  [1:0]  io_q_24_b,
  input  [1:0]  io_q_25_b,
  input  [1:0]  io_q_26_b,
  input  [1:0]  io_q_27_b,
  input  [1:0]  io_q_28_b,
  input  [1:0]  io_q_29_b,
  input  [1:0]  io_r_0_b,
  input  [1:0]  io_r_1_b,
  input  [1:0]  io_r_2_b,
  input  [1:0]  io_r_3_b,
  input  [1:0]  io_r_4_b,
  input  [1:0]  io_r_5_b,
  input  [1:0]  io_r_6_b,
  input  [1:0]  io_r_7_b,
  input  [1:0]  io_r_8_b,
  input  [1:0]  io_r_9_b,
  input  [1:0]  io_r_10_b,
  input  [1:0]  io_r_11_b,
  input  [1:0]  io_r_12_b,
  input  [1:0]  io_r_13_b,
  input  [1:0]  io_r_14_b,
  input  [1:0]  io_r_15_b,
  input  [1:0]  io_r_16_b,
  input  [1:0]  io_r_17_b,
  input  [1:0]  io_r_18_b,
  input  [1:0]  io_r_19_b,
  input  [1:0]  io_r_20_b,
  input  [1:0]  io_r_21_b,
  input  [1:0]  io_r_22_b,
  input  [1:0]  io_r_23_b,
  input  [1:0]  io_r_24_b,
  input  [1:0]  io_r_25_b,
  input  [1:0]  io_r_26_b,
  input  [1:0]  io_r_27_b,
  input  [1:0]  io_r_28_b,
  input  [1:0]  io_r_29_b,
  input  [1:0]  io_r_30_b,
  input  [1:0]  io_r_31_b,
  input  [1:0]  io_r_32_b,
  input  [1:0]  io_r_33_b,
  input  [1:0]  io_r_34_b,
  input  [1:0]  io_r_35_b,
  input  [1:0]  io_r_36_b,
  input  [1:0]  io_r_37_b,
  input  [1:0]  io_r_38_b,
  input  [1:0]  io_r_39_b,
  input  [1:0]  io_r_40_b,
  input  [1:0]  io_r_41_b,
  input  [1:0]  io_r_42_b,
  input  [1:0]  io_r_43_b,
  input  [1:0]  io_r_44_b,
  input  [1:0]  io_r_45_b,
  input  [1:0]  io_r_46_b,
  input  [1:0]  io_r_47_b,
  input  [1:0]  io_r_48_b,
  input  [1:0]  io_r_49_b,
  input  [1:0]  io_r_50_b,
  input  [1:0]  io_r_51_b,
  input  [1:0]  io_r_52_b,
  input  [1:0]  io_r_53_b,
  input  [1:0]  io_r_54_b,
  input  [1:0]  io_r_55_b,
  input  [1:0]  io_r_56_b,
  input  [1:0]  io_r_57_b,
  input  [1:0]  io_r_58_b,
  input  [1:0]  io_r_59_b,
  input  [1:0]  io_r_60_b,
  input  [1:0]  io_r_61_b,
  input  [1:0]  io_r_62_b,
  input  [1:0]  io_r_63_b,
  input  [1:0]  io_r_64_b,
  input  [1:0]  io_r_65_b,
  input  [1:0]  io_r_66_b,
  input  [1:0]  io_r_67_b,
  input  [1:0]  io_r_68_b,
  input  [1:0]  io_r_69_b,
  input  [1:0]  io_r_70_b,
  input  [1:0]  io_r_71_b,
  input  [1:0]  io_r_72_b,
  input  [1:0]  io_r_73_b,
  input  [1:0]  io_r_74_b,
  input  [1:0]  io_r_75_b,
  input  [1:0]  io_r_76_b,
  input  [1:0]  io_r_77_b,
  input  [1:0]  io_r_78_b,
  input  [1:0]  io_r_79_b,
  input  [1:0]  io_r_80_b,
  input  [1:0]  io_r_81_b,
  input  [1:0]  io_r_82_b,
  input  [1:0]  io_r_83_b,
  input  [1:0]  io_r_84_b,
  input  [1:0]  io_r_85_b,
  input  [1:0]  io_r_86_b,
  input  [1:0]  io_r_87_b,
  input  [1:0]  io_r_88_b,
  input  [1:0]  io_r_89_b,
  input  [1:0]  io_r_90_b,
  input  [1:0]  io_r_91_b,
  input  [1:0]  io_r_92_b,
  input  [1:0]  io_r_93_b,
  input  [1:0]  io_r_94_b,
  input  [1:0]  io_r_95_b,
  input  [1:0]  io_r_96_b,
  input  [1:0]  io_r_97_b,
  input  [1:0]  io_r_98_b,
  input  [1:0]  io_r_99_b,
  input  [1:0]  io_r_100_b,
  input  [1:0]  io_r_101_b,
  input  [1:0]  io_r_102_b,
  input  [1:0]  io_r_103_b,
  input  [1:0]  io_r_104_b,
  input  [1:0]  io_r_105_b,
  input  [1:0]  io_r_106_b,
  input  [1:0]  io_r_107_b,
  input  [1:0]  io_r_108_b,
  input  [1:0]  io_r_109_b,
  input  [1:0]  io_r_110_b,
  input  [1:0]  io_r_111_b,
  input  [1:0]  io_r_112_b,
  input  [1:0]  io_r_113_b,
  input  [1:0]  io_r_114_b,
  input  [1:0]  io_r_115_b,
  input  [1:0]  io_r_116_b,
  input  [1:0]  io_r_117_b,
  input  [1:0]  io_r_118_b,
  input  [1:0]  io_r_119_b,
  input  [1:0]  io_r_120_b,
  input  [1:0]  io_r_121_b,
  input  [1:0]  io_r_122_b,
  input  [1:0]  io_r_123_b,
  input  [1:0]  io_r_124_b,
  input  [1:0]  io_r_125_b,
  input  [1:0]  io_r_126_b,
  input  [1:0]  io_r_127_b,
  input  [1:0]  io_r_128_b,
  input  [1:0]  io_r_129_b,
  input  [1:0]  io_r_130_b,
  input  [1:0]  io_r_131_b,
  input  [1:0]  io_r_132_b,
  input  [1:0]  io_r_133_b,
  input  [1:0]  io_r_134_b,
  input  [1:0]  io_r_135_b,
  input  [1:0]  io_r_136_b,
  input  [1:0]  io_r_137_b,
  input  [1:0]  io_r_138_b,
  input  [1:0]  io_r_139_b,
  input  [1:0]  io_r_140_b,
  input  [1:0]  io_r_141_b,
  input  [1:0]  io_r_142_b,
  input  [1:0]  io_r_143_b,
  input  [1:0]  io_r_144_b,
  input  [1:0]  io_r_145_b,
  input  [1:0]  io_r_146_b,
  input  [1:0]  io_r_147_b,
  input  [1:0]  io_r_148_b,
  input  [1:0]  io_r_149_b,
  input  [1:0]  io_r_150_b,
  input  [1:0]  io_r_151_b,
  input  [1:0]  io_r_152_b,
  input  [1:0]  io_r_153_b,
  input  [1:0]  io_r_154_b,
  input  [1:0]  io_r_155_b,
  input  [1:0]  io_r_156_b,
  input  [1:0]  io_r_157_b,
  input  [1:0]  io_r_158_b,
  input  [1:0]  io_r_159_b,
  input  [1:0]  io_r_160_b,
  input  [1:0]  io_r_161_b,
  input  [1:0]  io_r_162_b,
  input  [1:0]  io_r_163_b,
  input  [1:0]  io_r_164_b,
  input  [1:0]  io_r_165_b,
  input  [1:0]  io_r_166_b,
  input  [1:0]  io_r_167_b,
  input  [1:0]  io_r_168_b,
  input  [1:0]  io_r_169_b,
  input  [1:0]  io_r_170_b,
  input  [1:0]  io_r_171_b,
  input  [1:0]  io_r_172_b,
  input  [1:0]  io_r_173_b,
  input  [1:0]  io_r_174_b,
  input  [1:0]  io_r_175_b,
  input  [1:0]  io_r_176_b,
  input  [1:0]  io_r_177_b,
  input  [1:0]  io_r_178_b,
  input  [1:0]  io_r_179_b,
  input  [1:0]  io_r_180_b,
  input  [1:0]  io_r_181_b,
  input  [1:0]  io_r_182_b,
  input  [1:0]  io_r_183_b,
  input  [1:0]  io_r_184_b,
  input  [1:0]  io_r_185_b,
  input  [1:0]  io_r_186_b,
  input  [1:0]  io_r_187_b,
  input  [1:0]  io_r_188_b,
  input  [1:0]  io_r_189_b,
  input  [1:0]  io_r_190_b,
  input  [1:0]  io_r_191_b,
  input  [1:0]  io_r_192_b,
  input  [1:0]  io_r_193_b,
  input  [1:0]  io_r_194_b,
  input  [1:0]  io_r_195_b,
  input  [1:0]  io_r_196_b,
  input  [1:0]  io_r_197_b,
  input  [1:0]  io_r_198_b,
  input  [1:0]  io_r_199_b,
  input  [1:0]  io_r_200_b,
  input  [1:0]  io_r_201_b,
  input  [1:0]  io_r_202_b,
  input  [1:0]  io_r_203_b,
  input  [1:0]  io_r_204_b,
  input  [1:0]  io_r_205_b,
  input  [1:0]  io_r_206_b,
  input  [1:0]  io_r_207_b,
  input  [1:0]  io_r_208_b,
  input  [1:0]  io_r_209_b,
  input  [1:0]  io_r_210_b,
  input  [1:0]  io_r_211_b,
  input  [1:0]  io_r_212_b,
  input  [1:0]  io_r_213_b,
  input  [1:0]  io_r_214_b,
  input  [1:0]  io_r_215_b,
  input  [1:0]  io_r_216_b,
  input  [1:0]  io_r_217_b,
  input  [1:0]  io_r_218_b,
  input  [1:0]  io_r_219_b,
  input  [1:0]  io_r_220_b,
  input  [1:0]  io_r_221_b,
  input  [1:0]  io_r_222_b,
  input  [1:0]  io_r_223_b,
  input  [1:0]  io_r_224_b,
  input  [1:0]  io_r_225_b,
  input  [1:0]  io_r_226_b,
  input  [1:0]  io_r_227_b,
  input  [1:0]  io_r_228_b,
  input  [1:0]  io_r_229_b,
  input  [1:0]  io_r_230_b,
  input  [1:0]  io_r_231_b,
  input  [1:0]  io_r_232_b,
  input  [1:0]  io_r_233_b,
  input  [1:0]  io_r_234_b,
  input  [1:0]  io_r_235_b,
  input  [1:0]  io_r_236_b,
  input  [1:0]  io_r_237_b,
  input  [1:0]  io_r_238_b,
  input  [1:0]  io_r_239_b,
  input  [1:0]  io_r_240_b,
  input  [1:0]  io_r_241_b,
  input  [1:0]  io_r_242_b,
  input  [1:0]  io_r_243_b,
  input  [1:0]  io_r_244_b,
  input  [1:0]  io_r_245_b,
  input  [1:0]  io_r_246_b,
  input  [1:0]  io_r_247_b,
  input  [1:0]  io_r_248_b,
  input  [1:0]  io_r_249_b,
  input  [1:0]  io_r_250_b,
  input  [1:0]  io_r_251_b,
  input  [1:0]  io_r_252_b,
  input  [1:0]  io_r_253_b,
  input  [1:0]  io_r_254_b,
  input  [1:0]  io_r_255_b,
  input  [1:0]  io_r_256_b,
  input  [1:0]  io_r_257_b,
  input  [1:0]  io_r_258_b,
  input  [1:0]  io_r_259_b,
  input  [1:0]  io_r_260_b,
  input  [1:0]  io_r_261_b,
  input  [1:0]  io_r_262_b,
  input  [1:0]  io_r_263_b,
  input  [1:0]  io_r_264_b,
  input  [1:0]  io_r_265_b,
  input  [1:0]  io_r_266_b,
  input  [1:0]  io_r_267_b,
  input  [1:0]  io_r_268_b,
  input  [1:0]  io_r_269_b,
  input  [1:0]  io_r_270_b,
  input  [1:0]  io_r_271_b,
  input  [1:0]  io_r_272_b,
  input  [1:0]  io_r_273_b,
  input  [1:0]  io_r_274_b,
  input  [1:0]  io_r_275_b,
  input  [1:0]  io_r_276_b,
  input  [1:0]  io_r_277_b,
  input  [1:0]  io_r_278_b,
  input  [1:0]  io_r_279_b,
  input  [1:0]  io_r_280_b,
  input  [1:0]  io_r_281_b,
  input  [1:0]  io_r_282_b,
  input  [1:0]  io_r_283_b,
  input  [1:0]  io_r_284_b,
  input  [1:0]  io_r_285_b,
  input  [1:0]  io_r_286_b,
  input  [1:0]  io_r_287_b,
  input  [1:0]  io_r_288_b,
  input  [1:0]  io_r_289_b,
  input  [1:0]  io_r_290_b,
  input  [1:0]  io_r_291_b,
  input  [1:0]  io_r_292_b,
  input  [1:0]  io_r_293_b,
  input  [1:0]  io_r_294_b,
  input  [1:0]  io_r_295_b,
  input  [1:0]  io_r_296_b,
  input  [1:0]  io_r_297_b,
  input  [1:0]  io_r_298_b,
  input  [1:0]  io_r_299_b,
  input         io_start,
  output [15:0] io_result,
  output        io_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
`endif // RANDOMIZE_REG_INIT
  wire [1:0] array_0_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_0_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_1_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_1_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_2_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_2_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_3_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_3_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_4_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_4_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_5_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_5_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_6_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_6_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_7_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_7_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_8_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_8_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_9_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_9_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_10_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_10_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_11_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_11_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_12_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_12_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_13_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_13_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_14_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_14_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_15_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_15_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_16_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_16_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_17_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_17_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_18_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_18_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_19_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_19_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_20_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_20_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_21_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_21_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_22_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_22_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_23_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_23_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_24_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_24_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_25_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_25_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_26_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_26_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_27_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_27_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_28_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_28_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_29_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_29_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_v_o; // @[SWChisel.scala 170:39]
  wire  r_count_0_clock; // @[SWChisel.scala 171:41]
  wire  r_count_0_reset; // @[SWChisel.scala 171:41]
  wire  r_count_0_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_0_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_1_clock; // @[SWChisel.scala 171:41]
  wire  r_count_1_reset; // @[SWChisel.scala 171:41]
  wire  r_count_1_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_1_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_2_clock; // @[SWChisel.scala 171:41]
  wire  r_count_2_reset; // @[SWChisel.scala 171:41]
  wire  r_count_2_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_2_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_3_clock; // @[SWChisel.scala 171:41]
  wire  r_count_3_reset; // @[SWChisel.scala 171:41]
  wire  r_count_3_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_3_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_4_clock; // @[SWChisel.scala 171:41]
  wire  r_count_4_reset; // @[SWChisel.scala 171:41]
  wire  r_count_4_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_4_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_5_clock; // @[SWChisel.scala 171:41]
  wire  r_count_5_reset; // @[SWChisel.scala 171:41]
  wire  r_count_5_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_5_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_6_clock; // @[SWChisel.scala 171:41]
  wire  r_count_6_reset; // @[SWChisel.scala 171:41]
  wire  r_count_6_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_6_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_7_clock; // @[SWChisel.scala 171:41]
  wire  r_count_7_reset; // @[SWChisel.scala 171:41]
  wire  r_count_7_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_7_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_8_clock; // @[SWChisel.scala 171:41]
  wire  r_count_8_reset; // @[SWChisel.scala 171:41]
  wire  r_count_8_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_8_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_9_clock; // @[SWChisel.scala 171:41]
  wire  r_count_9_reset; // @[SWChisel.scala 171:41]
  wire  r_count_9_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_9_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_10_clock; // @[SWChisel.scala 171:41]
  wire  r_count_10_reset; // @[SWChisel.scala 171:41]
  wire  r_count_10_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_10_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_11_clock; // @[SWChisel.scala 171:41]
  wire  r_count_11_reset; // @[SWChisel.scala 171:41]
  wire  r_count_11_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_11_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_12_clock; // @[SWChisel.scala 171:41]
  wire  r_count_12_reset; // @[SWChisel.scala 171:41]
  wire  r_count_12_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_12_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_13_clock; // @[SWChisel.scala 171:41]
  wire  r_count_13_reset; // @[SWChisel.scala 171:41]
  wire  r_count_13_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_13_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_14_clock; // @[SWChisel.scala 171:41]
  wire  r_count_14_reset; // @[SWChisel.scala 171:41]
  wire  r_count_14_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_14_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_15_clock; // @[SWChisel.scala 171:41]
  wire  r_count_15_reset; // @[SWChisel.scala 171:41]
  wire  r_count_15_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_15_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_16_clock; // @[SWChisel.scala 171:41]
  wire  r_count_16_reset; // @[SWChisel.scala 171:41]
  wire  r_count_16_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_16_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_17_clock; // @[SWChisel.scala 171:41]
  wire  r_count_17_reset; // @[SWChisel.scala 171:41]
  wire  r_count_17_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_17_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_18_clock; // @[SWChisel.scala 171:41]
  wire  r_count_18_reset; // @[SWChisel.scala 171:41]
  wire  r_count_18_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_18_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_19_clock; // @[SWChisel.scala 171:41]
  wire  r_count_19_reset; // @[SWChisel.scala 171:41]
  wire  r_count_19_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_19_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_20_clock; // @[SWChisel.scala 171:41]
  wire  r_count_20_reset; // @[SWChisel.scala 171:41]
  wire  r_count_20_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_20_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_21_clock; // @[SWChisel.scala 171:41]
  wire  r_count_21_reset; // @[SWChisel.scala 171:41]
  wire  r_count_21_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_21_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_22_clock; // @[SWChisel.scala 171:41]
  wire  r_count_22_reset; // @[SWChisel.scala 171:41]
  wire  r_count_22_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_22_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_23_clock; // @[SWChisel.scala 171:41]
  wire  r_count_23_reset; // @[SWChisel.scala 171:41]
  wire  r_count_23_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_23_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_24_clock; // @[SWChisel.scala 171:41]
  wire  r_count_24_reset; // @[SWChisel.scala 171:41]
  wire  r_count_24_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_24_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_25_clock; // @[SWChisel.scala 171:41]
  wire  r_count_25_reset; // @[SWChisel.scala 171:41]
  wire  r_count_25_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_25_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_26_clock; // @[SWChisel.scala 171:41]
  wire  r_count_26_reset; // @[SWChisel.scala 171:41]
  wire  r_count_26_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_26_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_27_clock; // @[SWChisel.scala 171:41]
  wire  r_count_27_reset; // @[SWChisel.scala 171:41]
  wire  r_count_27_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_27_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_28_clock; // @[SWChisel.scala 171:41]
  wire  r_count_28_reset; // @[SWChisel.scala 171:41]
  wire  r_count_28_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_28_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_29_clock; // @[SWChisel.scala 171:41]
  wire  r_count_29_reset; // @[SWChisel.scala 171:41]
  wire  r_count_29_io_en; // @[SWChisel.scala 171:41]
  wire [8:0] r_count_29_io_out; // @[SWChisel.scala 171:41]
  wire  max_clock; // @[SWChisel.scala 174:19]
  wire  max_reset; // @[SWChisel.scala 174:19]
  wire  max_io_start; // @[SWChisel.scala 174:19]
  wire [15:0] max_io_in; // @[SWChisel.scala 174:19]
  wire  max_io_done; // @[SWChisel.scala 174:19]
  wire [15:0] max_io_out; // @[SWChisel.scala 174:19]
  reg [15:0] E_0; // @[SWChisel.scala 162:18]
  reg [15:0] E_1; // @[SWChisel.scala 162:18]
  reg [15:0] E_2; // @[SWChisel.scala 162:18]
  reg [15:0] E_3; // @[SWChisel.scala 162:18]
  reg [15:0] E_4; // @[SWChisel.scala 162:18]
  reg [15:0] E_5; // @[SWChisel.scala 162:18]
  reg [15:0] E_6; // @[SWChisel.scala 162:18]
  reg [15:0] E_7; // @[SWChisel.scala 162:18]
  reg [15:0] E_8; // @[SWChisel.scala 162:18]
  reg [15:0] E_9; // @[SWChisel.scala 162:18]
  reg [15:0] E_10; // @[SWChisel.scala 162:18]
  reg [15:0] E_11; // @[SWChisel.scala 162:18]
  reg [15:0] E_12; // @[SWChisel.scala 162:18]
  reg [15:0] E_13; // @[SWChisel.scala 162:18]
  reg [15:0] E_14; // @[SWChisel.scala 162:18]
  reg [15:0] E_15; // @[SWChisel.scala 162:18]
  reg [15:0] E_16; // @[SWChisel.scala 162:18]
  reg [15:0] E_17; // @[SWChisel.scala 162:18]
  reg [15:0] E_18; // @[SWChisel.scala 162:18]
  reg [15:0] E_19; // @[SWChisel.scala 162:18]
  reg [15:0] E_20; // @[SWChisel.scala 162:18]
  reg [15:0] E_21; // @[SWChisel.scala 162:18]
  reg [15:0] E_22; // @[SWChisel.scala 162:18]
  reg [15:0] E_23; // @[SWChisel.scala 162:18]
  reg [15:0] E_24; // @[SWChisel.scala 162:18]
  reg [15:0] E_25; // @[SWChisel.scala 162:18]
  reg [15:0] E_26; // @[SWChisel.scala 162:18]
  reg [15:0] E_27; // @[SWChisel.scala 162:18]
  reg [15:0] E_28; // @[SWChisel.scala 162:18]
  reg [15:0] E_29; // @[SWChisel.scala 162:18]
  reg [15:0] F_1; // @[SWChisel.scala 163:18]
  reg [15:0] F_2; // @[SWChisel.scala 163:18]
  reg [15:0] F_3; // @[SWChisel.scala 163:18]
  reg [15:0] F_4; // @[SWChisel.scala 163:18]
  reg [15:0] F_5; // @[SWChisel.scala 163:18]
  reg [15:0] F_6; // @[SWChisel.scala 163:18]
  reg [15:0] F_7; // @[SWChisel.scala 163:18]
  reg [15:0] F_8; // @[SWChisel.scala 163:18]
  reg [15:0] F_9; // @[SWChisel.scala 163:18]
  reg [15:0] F_10; // @[SWChisel.scala 163:18]
  reg [15:0] F_11; // @[SWChisel.scala 163:18]
  reg [15:0] F_12; // @[SWChisel.scala 163:18]
  reg [15:0] F_13; // @[SWChisel.scala 163:18]
  reg [15:0] F_14; // @[SWChisel.scala 163:18]
  reg [15:0] F_15; // @[SWChisel.scala 163:18]
  reg [15:0] F_16; // @[SWChisel.scala 163:18]
  reg [15:0] F_17; // @[SWChisel.scala 163:18]
  reg [15:0] F_18; // @[SWChisel.scala 163:18]
  reg [15:0] F_19; // @[SWChisel.scala 163:18]
  reg [15:0] F_20; // @[SWChisel.scala 163:18]
  reg [15:0] F_21; // @[SWChisel.scala 163:18]
  reg [15:0] F_22; // @[SWChisel.scala 163:18]
  reg [15:0] F_23; // @[SWChisel.scala 163:18]
  reg [15:0] F_24; // @[SWChisel.scala 163:18]
  reg [15:0] F_25; // @[SWChisel.scala 163:18]
  reg [15:0] F_26; // @[SWChisel.scala 163:18]
  reg [15:0] F_27; // @[SWChisel.scala 163:18]
  reg [15:0] F_28; // @[SWChisel.scala 163:18]
  reg [15:0] F_29; // @[SWChisel.scala 163:18]
  reg [15:0] V1_0; // @[SWChisel.scala 164:19]
  reg [15:0] V1_1; // @[SWChisel.scala 164:19]
  reg [15:0] V1_2; // @[SWChisel.scala 164:19]
  reg [15:0] V1_3; // @[SWChisel.scala 164:19]
  reg [15:0] V1_4; // @[SWChisel.scala 164:19]
  reg [15:0] V1_5; // @[SWChisel.scala 164:19]
  reg [15:0] V1_6; // @[SWChisel.scala 164:19]
  reg [15:0] V1_7; // @[SWChisel.scala 164:19]
  reg [15:0] V1_8; // @[SWChisel.scala 164:19]
  reg [15:0] V1_9; // @[SWChisel.scala 164:19]
  reg [15:0] V1_10; // @[SWChisel.scala 164:19]
  reg [15:0] V1_11; // @[SWChisel.scala 164:19]
  reg [15:0] V1_12; // @[SWChisel.scala 164:19]
  reg [15:0] V1_13; // @[SWChisel.scala 164:19]
  reg [15:0] V1_14; // @[SWChisel.scala 164:19]
  reg [15:0] V1_15; // @[SWChisel.scala 164:19]
  reg [15:0] V1_16; // @[SWChisel.scala 164:19]
  reg [15:0] V1_17; // @[SWChisel.scala 164:19]
  reg [15:0] V1_18; // @[SWChisel.scala 164:19]
  reg [15:0] V1_19; // @[SWChisel.scala 164:19]
  reg [15:0] V1_20; // @[SWChisel.scala 164:19]
  reg [15:0] V1_21; // @[SWChisel.scala 164:19]
  reg [15:0] V1_22; // @[SWChisel.scala 164:19]
  reg [15:0] V1_23; // @[SWChisel.scala 164:19]
  reg [15:0] V1_24; // @[SWChisel.scala 164:19]
  reg [15:0] V1_25; // @[SWChisel.scala 164:19]
  reg [15:0] V1_26; // @[SWChisel.scala 164:19]
  reg [15:0] V1_27; // @[SWChisel.scala 164:19]
  reg [15:0] V1_28; // @[SWChisel.scala 164:19]
  reg [15:0] V1_29; // @[SWChisel.scala 164:19]
  reg [15:0] V1_30; // @[SWChisel.scala 164:19]
  reg [15:0] V2_0; // @[SWChisel.scala 166:19]
  reg [15:0] V2_1; // @[SWChisel.scala 166:19]
  reg [15:0] V2_2; // @[SWChisel.scala 166:19]
  reg [15:0] V2_3; // @[SWChisel.scala 166:19]
  reg [15:0] V2_4; // @[SWChisel.scala 166:19]
  reg [15:0] V2_5; // @[SWChisel.scala 166:19]
  reg [15:0] V2_6; // @[SWChisel.scala 166:19]
  reg [15:0] V2_7; // @[SWChisel.scala 166:19]
  reg [15:0] V2_8; // @[SWChisel.scala 166:19]
  reg [15:0] V2_9; // @[SWChisel.scala 166:19]
  reg [15:0] V2_10; // @[SWChisel.scala 166:19]
  reg [15:0] V2_11; // @[SWChisel.scala 166:19]
  reg [15:0] V2_12; // @[SWChisel.scala 166:19]
  reg [15:0] V2_13; // @[SWChisel.scala 166:19]
  reg [15:0] V2_14; // @[SWChisel.scala 166:19]
  reg [15:0] V2_15; // @[SWChisel.scala 166:19]
  reg [15:0] V2_16; // @[SWChisel.scala 166:19]
  reg [15:0] V2_17; // @[SWChisel.scala 166:19]
  reg [15:0] V2_18; // @[SWChisel.scala 166:19]
  reg [15:0] V2_19; // @[SWChisel.scala 166:19]
  reg [15:0] V2_20; // @[SWChisel.scala 166:19]
  reg [15:0] V2_21; // @[SWChisel.scala 166:19]
  reg [15:0] V2_22; // @[SWChisel.scala 166:19]
  reg [15:0] V2_23; // @[SWChisel.scala 166:19]
  reg [15:0] V2_24; // @[SWChisel.scala 166:19]
  reg [15:0] V2_25; // @[SWChisel.scala 166:19]
  reg [15:0] V2_26; // @[SWChisel.scala 166:19]
  reg [15:0] V2_27; // @[SWChisel.scala 166:19]
  reg [15:0] V2_28; // @[SWChisel.scala 166:19]
  reg [15:0] V2_29; // @[SWChisel.scala 166:19]
  reg  start_reg_0; // @[SWChisel.scala 167:26]
  reg  start_reg_1; // @[SWChisel.scala 167:26]
  reg  start_reg_2; // @[SWChisel.scala 167:26]
  reg  start_reg_3; // @[SWChisel.scala 167:26]
  reg  start_reg_4; // @[SWChisel.scala 167:26]
  reg  start_reg_5; // @[SWChisel.scala 167:26]
  reg  start_reg_6; // @[SWChisel.scala 167:26]
  reg  start_reg_7; // @[SWChisel.scala 167:26]
  reg  start_reg_8; // @[SWChisel.scala 167:26]
  reg  start_reg_9; // @[SWChisel.scala 167:26]
  reg  start_reg_10; // @[SWChisel.scala 167:26]
  reg  start_reg_11; // @[SWChisel.scala 167:26]
  reg  start_reg_12; // @[SWChisel.scala 167:26]
  reg  start_reg_13; // @[SWChisel.scala 167:26]
  reg  start_reg_14; // @[SWChisel.scala 167:26]
  reg  start_reg_15; // @[SWChisel.scala 167:26]
  reg  start_reg_16; // @[SWChisel.scala 167:26]
  reg  start_reg_17; // @[SWChisel.scala 167:26]
  reg  start_reg_18; // @[SWChisel.scala 167:26]
  reg  start_reg_19; // @[SWChisel.scala 167:26]
  reg  start_reg_20; // @[SWChisel.scala 167:26]
  reg  start_reg_21; // @[SWChisel.scala 167:26]
  reg  start_reg_22; // @[SWChisel.scala 167:26]
  reg  start_reg_23; // @[SWChisel.scala 167:26]
  reg  start_reg_24; // @[SWChisel.scala 167:26]
  reg  start_reg_25; // @[SWChisel.scala 167:26]
  reg  start_reg_26; // @[SWChisel.scala 167:26]
  reg  start_reg_27; // @[SWChisel.scala 167:26]
  reg  start_reg_28; // @[SWChisel.scala 167:26]
  reg  start_reg_29; // @[SWChisel.scala 167:26]
  wire [1:0] _GEN_91 = 9'h1 == r_count_0_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_92 = 9'h2 == r_count_0_io_out ? io_r_2_b : _GEN_91; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_93 = 9'h3 == r_count_0_io_out ? io_r_3_b : _GEN_92; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_94 = 9'h4 == r_count_0_io_out ? io_r_4_b : _GEN_93; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_95 = 9'h5 == r_count_0_io_out ? io_r_5_b : _GEN_94; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_96 = 9'h6 == r_count_0_io_out ? io_r_6_b : _GEN_95; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_97 = 9'h7 == r_count_0_io_out ? io_r_7_b : _GEN_96; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_98 = 9'h8 == r_count_0_io_out ? io_r_8_b : _GEN_97; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_99 = 9'h9 == r_count_0_io_out ? io_r_9_b : _GEN_98; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_100 = 9'ha == r_count_0_io_out ? io_r_10_b : _GEN_99; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_101 = 9'hb == r_count_0_io_out ? io_r_11_b : _GEN_100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_102 = 9'hc == r_count_0_io_out ? io_r_12_b : _GEN_101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_103 = 9'hd == r_count_0_io_out ? io_r_13_b : _GEN_102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_104 = 9'he == r_count_0_io_out ? io_r_14_b : _GEN_103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_105 = 9'hf == r_count_0_io_out ? io_r_15_b : _GEN_104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_106 = 9'h10 == r_count_0_io_out ? io_r_16_b : _GEN_105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_107 = 9'h11 == r_count_0_io_out ? io_r_17_b : _GEN_106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_108 = 9'h12 == r_count_0_io_out ? io_r_18_b : _GEN_107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_109 = 9'h13 == r_count_0_io_out ? io_r_19_b : _GEN_108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_110 = 9'h14 == r_count_0_io_out ? io_r_20_b : _GEN_109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_111 = 9'h15 == r_count_0_io_out ? io_r_21_b : _GEN_110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_112 = 9'h16 == r_count_0_io_out ? io_r_22_b : _GEN_111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_113 = 9'h17 == r_count_0_io_out ? io_r_23_b : _GEN_112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_114 = 9'h18 == r_count_0_io_out ? io_r_24_b : _GEN_113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_115 = 9'h19 == r_count_0_io_out ? io_r_25_b : _GEN_114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_116 = 9'h1a == r_count_0_io_out ? io_r_26_b : _GEN_115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_117 = 9'h1b == r_count_0_io_out ? io_r_27_b : _GEN_116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_118 = 9'h1c == r_count_0_io_out ? io_r_28_b : _GEN_117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_119 = 9'h1d == r_count_0_io_out ? io_r_29_b : _GEN_118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_120 = 9'h1e == r_count_0_io_out ? io_r_30_b : _GEN_119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_121 = 9'h1f == r_count_0_io_out ? io_r_31_b : _GEN_120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_122 = 9'h20 == r_count_0_io_out ? io_r_32_b : _GEN_121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_123 = 9'h21 == r_count_0_io_out ? io_r_33_b : _GEN_122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_124 = 9'h22 == r_count_0_io_out ? io_r_34_b : _GEN_123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_125 = 9'h23 == r_count_0_io_out ? io_r_35_b : _GEN_124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_126 = 9'h24 == r_count_0_io_out ? io_r_36_b : _GEN_125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_127 = 9'h25 == r_count_0_io_out ? io_r_37_b : _GEN_126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_128 = 9'h26 == r_count_0_io_out ? io_r_38_b : _GEN_127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_129 = 9'h27 == r_count_0_io_out ? io_r_39_b : _GEN_128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_130 = 9'h28 == r_count_0_io_out ? io_r_40_b : _GEN_129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_131 = 9'h29 == r_count_0_io_out ? io_r_41_b : _GEN_130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_132 = 9'h2a == r_count_0_io_out ? io_r_42_b : _GEN_131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_133 = 9'h2b == r_count_0_io_out ? io_r_43_b : _GEN_132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_134 = 9'h2c == r_count_0_io_out ? io_r_44_b : _GEN_133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_135 = 9'h2d == r_count_0_io_out ? io_r_45_b : _GEN_134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_136 = 9'h2e == r_count_0_io_out ? io_r_46_b : _GEN_135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_137 = 9'h2f == r_count_0_io_out ? io_r_47_b : _GEN_136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_138 = 9'h30 == r_count_0_io_out ? io_r_48_b : _GEN_137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_139 = 9'h31 == r_count_0_io_out ? io_r_49_b : _GEN_138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_140 = 9'h32 == r_count_0_io_out ? io_r_50_b : _GEN_139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_141 = 9'h33 == r_count_0_io_out ? io_r_51_b : _GEN_140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_142 = 9'h34 == r_count_0_io_out ? io_r_52_b : _GEN_141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_143 = 9'h35 == r_count_0_io_out ? io_r_53_b : _GEN_142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_144 = 9'h36 == r_count_0_io_out ? io_r_54_b : _GEN_143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_145 = 9'h37 == r_count_0_io_out ? io_r_55_b : _GEN_144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_146 = 9'h38 == r_count_0_io_out ? io_r_56_b : _GEN_145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_147 = 9'h39 == r_count_0_io_out ? io_r_57_b : _GEN_146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_148 = 9'h3a == r_count_0_io_out ? io_r_58_b : _GEN_147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_149 = 9'h3b == r_count_0_io_out ? io_r_59_b : _GEN_148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_150 = 9'h3c == r_count_0_io_out ? io_r_60_b : _GEN_149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_151 = 9'h3d == r_count_0_io_out ? io_r_61_b : _GEN_150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_152 = 9'h3e == r_count_0_io_out ? io_r_62_b : _GEN_151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_153 = 9'h3f == r_count_0_io_out ? io_r_63_b : _GEN_152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_154 = 9'h40 == r_count_0_io_out ? io_r_64_b : _GEN_153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_155 = 9'h41 == r_count_0_io_out ? io_r_65_b : _GEN_154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_156 = 9'h42 == r_count_0_io_out ? io_r_66_b : _GEN_155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_157 = 9'h43 == r_count_0_io_out ? io_r_67_b : _GEN_156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_158 = 9'h44 == r_count_0_io_out ? io_r_68_b : _GEN_157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_159 = 9'h45 == r_count_0_io_out ? io_r_69_b : _GEN_158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_160 = 9'h46 == r_count_0_io_out ? io_r_70_b : _GEN_159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_161 = 9'h47 == r_count_0_io_out ? io_r_71_b : _GEN_160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_162 = 9'h48 == r_count_0_io_out ? io_r_72_b : _GEN_161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_163 = 9'h49 == r_count_0_io_out ? io_r_73_b : _GEN_162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_164 = 9'h4a == r_count_0_io_out ? io_r_74_b : _GEN_163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_165 = 9'h4b == r_count_0_io_out ? io_r_75_b : _GEN_164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_166 = 9'h4c == r_count_0_io_out ? io_r_76_b : _GEN_165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_167 = 9'h4d == r_count_0_io_out ? io_r_77_b : _GEN_166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_168 = 9'h4e == r_count_0_io_out ? io_r_78_b : _GEN_167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_169 = 9'h4f == r_count_0_io_out ? io_r_79_b : _GEN_168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_170 = 9'h50 == r_count_0_io_out ? io_r_80_b : _GEN_169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_171 = 9'h51 == r_count_0_io_out ? io_r_81_b : _GEN_170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_172 = 9'h52 == r_count_0_io_out ? io_r_82_b : _GEN_171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_173 = 9'h53 == r_count_0_io_out ? io_r_83_b : _GEN_172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_174 = 9'h54 == r_count_0_io_out ? io_r_84_b : _GEN_173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_175 = 9'h55 == r_count_0_io_out ? io_r_85_b : _GEN_174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_176 = 9'h56 == r_count_0_io_out ? io_r_86_b : _GEN_175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_177 = 9'h57 == r_count_0_io_out ? io_r_87_b : _GEN_176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_178 = 9'h58 == r_count_0_io_out ? io_r_88_b : _GEN_177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_179 = 9'h59 == r_count_0_io_out ? io_r_89_b : _GEN_178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_180 = 9'h5a == r_count_0_io_out ? io_r_90_b : _GEN_179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_181 = 9'h5b == r_count_0_io_out ? io_r_91_b : _GEN_180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_182 = 9'h5c == r_count_0_io_out ? io_r_92_b : _GEN_181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_183 = 9'h5d == r_count_0_io_out ? io_r_93_b : _GEN_182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_184 = 9'h5e == r_count_0_io_out ? io_r_94_b : _GEN_183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_185 = 9'h5f == r_count_0_io_out ? io_r_95_b : _GEN_184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_186 = 9'h60 == r_count_0_io_out ? io_r_96_b : _GEN_185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_187 = 9'h61 == r_count_0_io_out ? io_r_97_b : _GEN_186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_188 = 9'h62 == r_count_0_io_out ? io_r_98_b : _GEN_187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_189 = 9'h63 == r_count_0_io_out ? io_r_99_b : _GEN_188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_190 = 9'h64 == r_count_0_io_out ? io_r_100_b : _GEN_189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_191 = 9'h65 == r_count_0_io_out ? io_r_101_b : _GEN_190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_192 = 9'h66 == r_count_0_io_out ? io_r_102_b : _GEN_191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_193 = 9'h67 == r_count_0_io_out ? io_r_103_b : _GEN_192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_194 = 9'h68 == r_count_0_io_out ? io_r_104_b : _GEN_193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_195 = 9'h69 == r_count_0_io_out ? io_r_105_b : _GEN_194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_196 = 9'h6a == r_count_0_io_out ? io_r_106_b : _GEN_195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_197 = 9'h6b == r_count_0_io_out ? io_r_107_b : _GEN_196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_198 = 9'h6c == r_count_0_io_out ? io_r_108_b : _GEN_197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_199 = 9'h6d == r_count_0_io_out ? io_r_109_b : _GEN_198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_200 = 9'h6e == r_count_0_io_out ? io_r_110_b : _GEN_199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_201 = 9'h6f == r_count_0_io_out ? io_r_111_b : _GEN_200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_202 = 9'h70 == r_count_0_io_out ? io_r_112_b : _GEN_201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_203 = 9'h71 == r_count_0_io_out ? io_r_113_b : _GEN_202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_204 = 9'h72 == r_count_0_io_out ? io_r_114_b : _GEN_203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_205 = 9'h73 == r_count_0_io_out ? io_r_115_b : _GEN_204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_206 = 9'h74 == r_count_0_io_out ? io_r_116_b : _GEN_205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_207 = 9'h75 == r_count_0_io_out ? io_r_117_b : _GEN_206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_208 = 9'h76 == r_count_0_io_out ? io_r_118_b : _GEN_207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_209 = 9'h77 == r_count_0_io_out ? io_r_119_b : _GEN_208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_210 = 9'h78 == r_count_0_io_out ? io_r_120_b : _GEN_209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_211 = 9'h79 == r_count_0_io_out ? io_r_121_b : _GEN_210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_212 = 9'h7a == r_count_0_io_out ? io_r_122_b : _GEN_211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_213 = 9'h7b == r_count_0_io_out ? io_r_123_b : _GEN_212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_214 = 9'h7c == r_count_0_io_out ? io_r_124_b : _GEN_213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_215 = 9'h7d == r_count_0_io_out ? io_r_125_b : _GEN_214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_216 = 9'h7e == r_count_0_io_out ? io_r_126_b : _GEN_215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_217 = 9'h7f == r_count_0_io_out ? io_r_127_b : _GEN_216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_218 = 9'h80 == r_count_0_io_out ? io_r_128_b : _GEN_217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_219 = 9'h81 == r_count_0_io_out ? io_r_129_b : _GEN_218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_220 = 9'h82 == r_count_0_io_out ? io_r_130_b : _GEN_219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_221 = 9'h83 == r_count_0_io_out ? io_r_131_b : _GEN_220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_222 = 9'h84 == r_count_0_io_out ? io_r_132_b : _GEN_221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_223 = 9'h85 == r_count_0_io_out ? io_r_133_b : _GEN_222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_224 = 9'h86 == r_count_0_io_out ? io_r_134_b : _GEN_223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_225 = 9'h87 == r_count_0_io_out ? io_r_135_b : _GEN_224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_226 = 9'h88 == r_count_0_io_out ? io_r_136_b : _GEN_225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_227 = 9'h89 == r_count_0_io_out ? io_r_137_b : _GEN_226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_228 = 9'h8a == r_count_0_io_out ? io_r_138_b : _GEN_227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_229 = 9'h8b == r_count_0_io_out ? io_r_139_b : _GEN_228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_230 = 9'h8c == r_count_0_io_out ? io_r_140_b : _GEN_229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_231 = 9'h8d == r_count_0_io_out ? io_r_141_b : _GEN_230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_232 = 9'h8e == r_count_0_io_out ? io_r_142_b : _GEN_231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_233 = 9'h8f == r_count_0_io_out ? io_r_143_b : _GEN_232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_234 = 9'h90 == r_count_0_io_out ? io_r_144_b : _GEN_233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_235 = 9'h91 == r_count_0_io_out ? io_r_145_b : _GEN_234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_236 = 9'h92 == r_count_0_io_out ? io_r_146_b : _GEN_235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_237 = 9'h93 == r_count_0_io_out ? io_r_147_b : _GEN_236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_238 = 9'h94 == r_count_0_io_out ? io_r_148_b : _GEN_237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_239 = 9'h95 == r_count_0_io_out ? io_r_149_b : _GEN_238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_240 = 9'h96 == r_count_0_io_out ? io_r_150_b : _GEN_239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_241 = 9'h97 == r_count_0_io_out ? io_r_151_b : _GEN_240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_242 = 9'h98 == r_count_0_io_out ? io_r_152_b : _GEN_241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_243 = 9'h99 == r_count_0_io_out ? io_r_153_b : _GEN_242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_244 = 9'h9a == r_count_0_io_out ? io_r_154_b : _GEN_243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_245 = 9'h9b == r_count_0_io_out ? io_r_155_b : _GEN_244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_246 = 9'h9c == r_count_0_io_out ? io_r_156_b : _GEN_245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_247 = 9'h9d == r_count_0_io_out ? io_r_157_b : _GEN_246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_248 = 9'h9e == r_count_0_io_out ? io_r_158_b : _GEN_247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_249 = 9'h9f == r_count_0_io_out ? io_r_159_b : _GEN_248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_250 = 9'ha0 == r_count_0_io_out ? io_r_160_b : _GEN_249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_251 = 9'ha1 == r_count_0_io_out ? io_r_161_b : _GEN_250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_252 = 9'ha2 == r_count_0_io_out ? io_r_162_b : _GEN_251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_253 = 9'ha3 == r_count_0_io_out ? io_r_163_b : _GEN_252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_254 = 9'ha4 == r_count_0_io_out ? io_r_164_b : _GEN_253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_255 = 9'ha5 == r_count_0_io_out ? io_r_165_b : _GEN_254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_256 = 9'ha6 == r_count_0_io_out ? io_r_166_b : _GEN_255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_257 = 9'ha7 == r_count_0_io_out ? io_r_167_b : _GEN_256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_258 = 9'ha8 == r_count_0_io_out ? io_r_168_b : _GEN_257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_259 = 9'ha9 == r_count_0_io_out ? io_r_169_b : _GEN_258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_260 = 9'haa == r_count_0_io_out ? io_r_170_b : _GEN_259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_261 = 9'hab == r_count_0_io_out ? io_r_171_b : _GEN_260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_262 = 9'hac == r_count_0_io_out ? io_r_172_b : _GEN_261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_263 = 9'had == r_count_0_io_out ? io_r_173_b : _GEN_262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_264 = 9'hae == r_count_0_io_out ? io_r_174_b : _GEN_263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_265 = 9'haf == r_count_0_io_out ? io_r_175_b : _GEN_264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_266 = 9'hb0 == r_count_0_io_out ? io_r_176_b : _GEN_265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_267 = 9'hb1 == r_count_0_io_out ? io_r_177_b : _GEN_266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_268 = 9'hb2 == r_count_0_io_out ? io_r_178_b : _GEN_267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_269 = 9'hb3 == r_count_0_io_out ? io_r_179_b : _GEN_268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_270 = 9'hb4 == r_count_0_io_out ? io_r_180_b : _GEN_269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_271 = 9'hb5 == r_count_0_io_out ? io_r_181_b : _GEN_270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_272 = 9'hb6 == r_count_0_io_out ? io_r_182_b : _GEN_271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_273 = 9'hb7 == r_count_0_io_out ? io_r_183_b : _GEN_272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_274 = 9'hb8 == r_count_0_io_out ? io_r_184_b : _GEN_273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_275 = 9'hb9 == r_count_0_io_out ? io_r_185_b : _GEN_274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_276 = 9'hba == r_count_0_io_out ? io_r_186_b : _GEN_275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_277 = 9'hbb == r_count_0_io_out ? io_r_187_b : _GEN_276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_278 = 9'hbc == r_count_0_io_out ? io_r_188_b : _GEN_277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_279 = 9'hbd == r_count_0_io_out ? io_r_189_b : _GEN_278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_280 = 9'hbe == r_count_0_io_out ? io_r_190_b : _GEN_279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_281 = 9'hbf == r_count_0_io_out ? io_r_191_b : _GEN_280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_282 = 9'hc0 == r_count_0_io_out ? io_r_192_b : _GEN_281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_283 = 9'hc1 == r_count_0_io_out ? io_r_193_b : _GEN_282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_284 = 9'hc2 == r_count_0_io_out ? io_r_194_b : _GEN_283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_285 = 9'hc3 == r_count_0_io_out ? io_r_195_b : _GEN_284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_286 = 9'hc4 == r_count_0_io_out ? io_r_196_b : _GEN_285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_287 = 9'hc5 == r_count_0_io_out ? io_r_197_b : _GEN_286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_288 = 9'hc6 == r_count_0_io_out ? io_r_198_b : _GEN_287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_289 = 9'hc7 == r_count_0_io_out ? io_r_199_b : _GEN_288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_290 = 9'hc8 == r_count_0_io_out ? io_r_200_b : _GEN_289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_291 = 9'hc9 == r_count_0_io_out ? io_r_201_b : _GEN_290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_292 = 9'hca == r_count_0_io_out ? io_r_202_b : _GEN_291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_293 = 9'hcb == r_count_0_io_out ? io_r_203_b : _GEN_292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_294 = 9'hcc == r_count_0_io_out ? io_r_204_b : _GEN_293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_295 = 9'hcd == r_count_0_io_out ? io_r_205_b : _GEN_294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_296 = 9'hce == r_count_0_io_out ? io_r_206_b : _GEN_295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_297 = 9'hcf == r_count_0_io_out ? io_r_207_b : _GEN_296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_298 = 9'hd0 == r_count_0_io_out ? io_r_208_b : _GEN_297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_299 = 9'hd1 == r_count_0_io_out ? io_r_209_b : _GEN_298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_300 = 9'hd2 == r_count_0_io_out ? io_r_210_b : _GEN_299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_301 = 9'hd3 == r_count_0_io_out ? io_r_211_b : _GEN_300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_302 = 9'hd4 == r_count_0_io_out ? io_r_212_b : _GEN_301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_303 = 9'hd5 == r_count_0_io_out ? io_r_213_b : _GEN_302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_304 = 9'hd6 == r_count_0_io_out ? io_r_214_b : _GEN_303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_305 = 9'hd7 == r_count_0_io_out ? io_r_215_b : _GEN_304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_306 = 9'hd8 == r_count_0_io_out ? io_r_216_b : _GEN_305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_307 = 9'hd9 == r_count_0_io_out ? io_r_217_b : _GEN_306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_308 = 9'hda == r_count_0_io_out ? io_r_218_b : _GEN_307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_309 = 9'hdb == r_count_0_io_out ? io_r_219_b : _GEN_308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_310 = 9'hdc == r_count_0_io_out ? io_r_220_b : _GEN_309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_311 = 9'hdd == r_count_0_io_out ? io_r_221_b : _GEN_310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_312 = 9'hde == r_count_0_io_out ? io_r_222_b : _GEN_311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_313 = 9'hdf == r_count_0_io_out ? io_r_223_b : _GEN_312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_314 = 9'he0 == r_count_0_io_out ? io_r_224_b : _GEN_313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_315 = 9'he1 == r_count_0_io_out ? io_r_225_b : _GEN_314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_316 = 9'he2 == r_count_0_io_out ? io_r_226_b : _GEN_315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_317 = 9'he3 == r_count_0_io_out ? io_r_227_b : _GEN_316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_318 = 9'he4 == r_count_0_io_out ? io_r_228_b : _GEN_317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_319 = 9'he5 == r_count_0_io_out ? io_r_229_b : _GEN_318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_320 = 9'he6 == r_count_0_io_out ? io_r_230_b : _GEN_319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_321 = 9'he7 == r_count_0_io_out ? io_r_231_b : _GEN_320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_322 = 9'he8 == r_count_0_io_out ? io_r_232_b : _GEN_321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_323 = 9'he9 == r_count_0_io_out ? io_r_233_b : _GEN_322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_324 = 9'hea == r_count_0_io_out ? io_r_234_b : _GEN_323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_325 = 9'heb == r_count_0_io_out ? io_r_235_b : _GEN_324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_326 = 9'hec == r_count_0_io_out ? io_r_236_b : _GEN_325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_327 = 9'hed == r_count_0_io_out ? io_r_237_b : _GEN_326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_328 = 9'hee == r_count_0_io_out ? io_r_238_b : _GEN_327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_329 = 9'hef == r_count_0_io_out ? io_r_239_b : _GEN_328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_330 = 9'hf0 == r_count_0_io_out ? io_r_240_b : _GEN_329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_331 = 9'hf1 == r_count_0_io_out ? io_r_241_b : _GEN_330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_332 = 9'hf2 == r_count_0_io_out ? io_r_242_b : _GEN_331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_333 = 9'hf3 == r_count_0_io_out ? io_r_243_b : _GEN_332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_334 = 9'hf4 == r_count_0_io_out ? io_r_244_b : _GEN_333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_335 = 9'hf5 == r_count_0_io_out ? io_r_245_b : _GEN_334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_336 = 9'hf6 == r_count_0_io_out ? io_r_246_b : _GEN_335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_337 = 9'hf7 == r_count_0_io_out ? io_r_247_b : _GEN_336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_338 = 9'hf8 == r_count_0_io_out ? io_r_248_b : _GEN_337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_339 = 9'hf9 == r_count_0_io_out ? io_r_249_b : _GEN_338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_340 = 9'hfa == r_count_0_io_out ? io_r_250_b : _GEN_339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_341 = 9'hfb == r_count_0_io_out ? io_r_251_b : _GEN_340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_342 = 9'hfc == r_count_0_io_out ? io_r_252_b : _GEN_341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_343 = 9'hfd == r_count_0_io_out ? io_r_253_b : _GEN_342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_344 = 9'hfe == r_count_0_io_out ? io_r_254_b : _GEN_343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_345 = 9'hff == r_count_0_io_out ? io_r_255_b : _GEN_344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_346 = 9'h100 == r_count_0_io_out ? io_r_256_b : _GEN_345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_347 = 9'h101 == r_count_0_io_out ? io_r_257_b : _GEN_346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_348 = 9'h102 == r_count_0_io_out ? io_r_258_b : _GEN_347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_349 = 9'h103 == r_count_0_io_out ? io_r_259_b : _GEN_348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_350 = 9'h104 == r_count_0_io_out ? io_r_260_b : _GEN_349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_351 = 9'h105 == r_count_0_io_out ? io_r_261_b : _GEN_350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_352 = 9'h106 == r_count_0_io_out ? io_r_262_b : _GEN_351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_353 = 9'h107 == r_count_0_io_out ? io_r_263_b : _GEN_352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_354 = 9'h108 == r_count_0_io_out ? io_r_264_b : _GEN_353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_355 = 9'h109 == r_count_0_io_out ? io_r_265_b : _GEN_354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_356 = 9'h10a == r_count_0_io_out ? io_r_266_b : _GEN_355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_357 = 9'h10b == r_count_0_io_out ? io_r_267_b : _GEN_356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_358 = 9'h10c == r_count_0_io_out ? io_r_268_b : _GEN_357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_359 = 9'h10d == r_count_0_io_out ? io_r_269_b : _GEN_358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_360 = 9'h10e == r_count_0_io_out ? io_r_270_b : _GEN_359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_361 = 9'h10f == r_count_0_io_out ? io_r_271_b : _GEN_360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_362 = 9'h110 == r_count_0_io_out ? io_r_272_b : _GEN_361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_363 = 9'h111 == r_count_0_io_out ? io_r_273_b : _GEN_362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_364 = 9'h112 == r_count_0_io_out ? io_r_274_b : _GEN_363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_365 = 9'h113 == r_count_0_io_out ? io_r_275_b : _GEN_364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_366 = 9'h114 == r_count_0_io_out ? io_r_276_b : _GEN_365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_367 = 9'h115 == r_count_0_io_out ? io_r_277_b : _GEN_366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_368 = 9'h116 == r_count_0_io_out ? io_r_278_b : _GEN_367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_369 = 9'h117 == r_count_0_io_out ? io_r_279_b : _GEN_368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_370 = 9'h118 == r_count_0_io_out ? io_r_280_b : _GEN_369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_371 = 9'h119 == r_count_0_io_out ? io_r_281_b : _GEN_370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_372 = 9'h11a == r_count_0_io_out ? io_r_282_b : _GEN_371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_373 = 9'h11b == r_count_0_io_out ? io_r_283_b : _GEN_372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_374 = 9'h11c == r_count_0_io_out ? io_r_284_b : _GEN_373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_375 = 9'h11d == r_count_0_io_out ? io_r_285_b : _GEN_374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_376 = 9'h11e == r_count_0_io_out ? io_r_286_b : _GEN_375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_377 = 9'h11f == r_count_0_io_out ? io_r_287_b : _GEN_376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_378 = 9'h120 == r_count_0_io_out ? io_r_288_b : _GEN_377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_379 = 9'h121 == r_count_0_io_out ? io_r_289_b : _GEN_378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_380 = 9'h122 == r_count_0_io_out ? io_r_290_b : _GEN_379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_381 = 9'h123 == r_count_0_io_out ? io_r_291_b : _GEN_380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_382 = 9'h124 == r_count_0_io_out ? io_r_292_b : _GEN_381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_383 = 9'h125 == r_count_0_io_out ? io_r_293_b : _GEN_382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_384 = 9'h126 == r_count_0_io_out ? io_r_294_b : _GEN_383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_385 = 9'h127 == r_count_0_io_out ? io_r_295_b : _GEN_384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_386 = 9'h128 == r_count_0_io_out ? io_r_296_b : _GEN_385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_387 = 9'h129 == r_count_0_io_out ? io_r_297_b : _GEN_386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_388 = 9'h12a == r_count_0_io_out ? io_r_298_b : _GEN_387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_391 = 9'h1 == r_count_1_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_392 = 9'h2 == r_count_1_io_out ? io_r_2_b : _GEN_391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_393 = 9'h3 == r_count_1_io_out ? io_r_3_b : _GEN_392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_394 = 9'h4 == r_count_1_io_out ? io_r_4_b : _GEN_393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_395 = 9'h5 == r_count_1_io_out ? io_r_5_b : _GEN_394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_396 = 9'h6 == r_count_1_io_out ? io_r_6_b : _GEN_395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_397 = 9'h7 == r_count_1_io_out ? io_r_7_b : _GEN_396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_398 = 9'h8 == r_count_1_io_out ? io_r_8_b : _GEN_397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_399 = 9'h9 == r_count_1_io_out ? io_r_9_b : _GEN_398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_400 = 9'ha == r_count_1_io_out ? io_r_10_b : _GEN_399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_401 = 9'hb == r_count_1_io_out ? io_r_11_b : _GEN_400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_402 = 9'hc == r_count_1_io_out ? io_r_12_b : _GEN_401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_403 = 9'hd == r_count_1_io_out ? io_r_13_b : _GEN_402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_404 = 9'he == r_count_1_io_out ? io_r_14_b : _GEN_403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_405 = 9'hf == r_count_1_io_out ? io_r_15_b : _GEN_404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_406 = 9'h10 == r_count_1_io_out ? io_r_16_b : _GEN_405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_407 = 9'h11 == r_count_1_io_out ? io_r_17_b : _GEN_406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_408 = 9'h12 == r_count_1_io_out ? io_r_18_b : _GEN_407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_409 = 9'h13 == r_count_1_io_out ? io_r_19_b : _GEN_408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_410 = 9'h14 == r_count_1_io_out ? io_r_20_b : _GEN_409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_411 = 9'h15 == r_count_1_io_out ? io_r_21_b : _GEN_410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_412 = 9'h16 == r_count_1_io_out ? io_r_22_b : _GEN_411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_413 = 9'h17 == r_count_1_io_out ? io_r_23_b : _GEN_412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_414 = 9'h18 == r_count_1_io_out ? io_r_24_b : _GEN_413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_415 = 9'h19 == r_count_1_io_out ? io_r_25_b : _GEN_414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_416 = 9'h1a == r_count_1_io_out ? io_r_26_b : _GEN_415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_417 = 9'h1b == r_count_1_io_out ? io_r_27_b : _GEN_416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_418 = 9'h1c == r_count_1_io_out ? io_r_28_b : _GEN_417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_419 = 9'h1d == r_count_1_io_out ? io_r_29_b : _GEN_418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_420 = 9'h1e == r_count_1_io_out ? io_r_30_b : _GEN_419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_421 = 9'h1f == r_count_1_io_out ? io_r_31_b : _GEN_420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_422 = 9'h20 == r_count_1_io_out ? io_r_32_b : _GEN_421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_423 = 9'h21 == r_count_1_io_out ? io_r_33_b : _GEN_422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_424 = 9'h22 == r_count_1_io_out ? io_r_34_b : _GEN_423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_425 = 9'h23 == r_count_1_io_out ? io_r_35_b : _GEN_424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_426 = 9'h24 == r_count_1_io_out ? io_r_36_b : _GEN_425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_427 = 9'h25 == r_count_1_io_out ? io_r_37_b : _GEN_426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_428 = 9'h26 == r_count_1_io_out ? io_r_38_b : _GEN_427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_429 = 9'h27 == r_count_1_io_out ? io_r_39_b : _GEN_428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_430 = 9'h28 == r_count_1_io_out ? io_r_40_b : _GEN_429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_431 = 9'h29 == r_count_1_io_out ? io_r_41_b : _GEN_430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_432 = 9'h2a == r_count_1_io_out ? io_r_42_b : _GEN_431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_433 = 9'h2b == r_count_1_io_out ? io_r_43_b : _GEN_432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_434 = 9'h2c == r_count_1_io_out ? io_r_44_b : _GEN_433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_435 = 9'h2d == r_count_1_io_out ? io_r_45_b : _GEN_434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_436 = 9'h2e == r_count_1_io_out ? io_r_46_b : _GEN_435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_437 = 9'h2f == r_count_1_io_out ? io_r_47_b : _GEN_436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_438 = 9'h30 == r_count_1_io_out ? io_r_48_b : _GEN_437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_439 = 9'h31 == r_count_1_io_out ? io_r_49_b : _GEN_438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_440 = 9'h32 == r_count_1_io_out ? io_r_50_b : _GEN_439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_441 = 9'h33 == r_count_1_io_out ? io_r_51_b : _GEN_440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_442 = 9'h34 == r_count_1_io_out ? io_r_52_b : _GEN_441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_443 = 9'h35 == r_count_1_io_out ? io_r_53_b : _GEN_442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_444 = 9'h36 == r_count_1_io_out ? io_r_54_b : _GEN_443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_445 = 9'h37 == r_count_1_io_out ? io_r_55_b : _GEN_444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_446 = 9'h38 == r_count_1_io_out ? io_r_56_b : _GEN_445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_447 = 9'h39 == r_count_1_io_out ? io_r_57_b : _GEN_446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_448 = 9'h3a == r_count_1_io_out ? io_r_58_b : _GEN_447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_449 = 9'h3b == r_count_1_io_out ? io_r_59_b : _GEN_448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_450 = 9'h3c == r_count_1_io_out ? io_r_60_b : _GEN_449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_451 = 9'h3d == r_count_1_io_out ? io_r_61_b : _GEN_450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_452 = 9'h3e == r_count_1_io_out ? io_r_62_b : _GEN_451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_453 = 9'h3f == r_count_1_io_out ? io_r_63_b : _GEN_452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_454 = 9'h40 == r_count_1_io_out ? io_r_64_b : _GEN_453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_455 = 9'h41 == r_count_1_io_out ? io_r_65_b : _GEN_454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_456 = 9'h42 == r_count_1_io_out ? io_r_66_b : _GEN_455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_457 = 9'h43 == r_count_1_io_out ? io_r_67_b : _GEN_456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_458 = 9'h44 == r_count_1_io_out ? io_r_68_b : _GEN_457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_459 = 9'h45 == r_count_1_io_out ? io_r_69_b : _GEN_458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_460 = 9'h46 == r_count_1_io_out ? io_r_70_b : _GEN_459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_461 = 9'h47 == r_count_1_io_out ? io_r_71_b : _GEN_460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_462 = 9'h48 == r_count_1_io_out ? io_r_72_b : _GEN_461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_463 = 9'h49 == r_count_1_io_out ? io_r_73_b : _GEN_462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_464 = 9'h4a == r_count_1_io_out ? io_r_74_b : _GEN_463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_465 = 9'h4b == r_count_1_io_out ? io_r_75_b : _GEN_464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_466 = 9'h4c == r_count_1_io_out ? io_r_76_b : _GEN_465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_467 = 9'h4d == r_count_1_io_out ? io_r_77_b : _GEN_466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_468 = 9'h4e == r_count_1_io_out ? io_r_78_b : _GEN_467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_469 = 9'h4f == r_count_1_io_out ? io_r_79_b : _GEN_468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_470 = 9'h50 == r_count_1_io_out ? io_r_80_b : _GEN_469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_471 = 9'h51 == r_count_1_io_out ? io_r_81_b : _GEN_470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_472 = 9'h52 == r_count_1_io_out ? io_r_82_b : _GEN_471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_473 = 9'h53 == r_count_1_io_out ? io_r_83_b : _GEN_472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_474 = 9'h54 == r_count_1_io_out ? io_r_84_b : _GEN_473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_475 = 9'h55 == r_count_1_io_out ? io_r_85_b : _GEN_474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_476 = 9'h56 == r_count_1_io_out ? io_r_86_b : _GEN_475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_477 = 9'h57 == r_count_1_io_out ? io_r_87_b : _GEN_476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_478 = 9'h58 == r_count_1_io_out ? io_r_88_b : _GEN_477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_479 = 9'h59 == r_count_1_io_out ? io_r_89_b : _GEN_478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_480 = 9'h5a == r_count_1_io_out ? io_r_90_b : _GEN_479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_481 = 9'h5b == r_count_1_io_out ? io_r_91_b : _GEN_480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_482 = 9'h5c == r_count_1_io_out ? io_r_92_b : _GEN_481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_483 = 9'h5d == r_count_1_io_out ? io_r_93_b : _GEN_482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_484 = 9'h5e == r_count_1_io_out ? io_r_94_b : _GEN_483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_485 = 9'h5f == r_count_1_io_out ? io_r_95_b : _GEN_484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_486 = 9'h60 == r_count_1_io_out ? io_r_96_b : _GEN_485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_487 = 9'h61 == r_count_1_io_out ? io_r_97_b : _GEN_486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_488 = 9'h62 == r_count_1_io_out ? io_r_98_b : _GEN_487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_489 = 9'h63 == r_count_1_io_out ? io_r_99_b : _GEN_488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_490 = 9'h64 == r_count_1_io_out ? io_r_100_b : _GEN_489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_491 = 9'h65 == r_count_1_io_out ? io_r_101_b : _GEN_490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_492 = 9'h66 == r_count_1_io_out ? io_r_102_b : _GEN_491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_493 = 9'h67 == r_count_1_io_out ? io_r_103_b : _GEN_492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_494 = 9'h68 == r_count_1_io_out ? io_r_104_b : _GEN_493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_495 = 9'h69 == r_count_1_io_out ? io_r_105_b : _GEN_494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_496 = 9'h6a == r_count_1_io_out ? io_r_106_b : _GEN_495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_497 = 9'h6b == r_count_1_io_out ? io_r_107_b : _GEN_496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_498 = 9'h6c == r_count_1_io_out ? io_r_108_b : _GEN_497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_499 = 9'h6d == r_count_1_io_out ? io_r_109_b : _GEN_498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_500 = 9'h6e == r_count_1_io_out ? io_r_110_b : _GEN_499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_501 = 9'h6f == r_count_1_io_out ? io_r_111_b : _GEN_500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_502 = 9'h70 == r_count_1_io_out ? io_r_112_b : _GEN_501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_503 = 9'h71 == r_count_1_io_out ? io_r_113_b : _GEN_502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_504 = 9'h72 == r_count_1_io_out ? io_r_114_b : _GEN_503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_505 = 9'h73 == r_count_1_io_out ? io_r_115_b : _GEN_504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_506 = 9'h74 == r_count_1_io_out ? io_r_116_b : _GEN_505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_507 = 9'h75 == r_count_1_io_out ? io_r_117_b : _GEN_506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_508 = 9'h76 == r_count_1_io_out ? io_r_118_b : _GEN_507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_509 = 9'h77 == r_count_1_io_out ? io_r_119_b : _GEN_508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_510 = 9'h78 == r_count_1_io_out ? io_r_120_b : _GEN_509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_511 = 9'h79 == r_count_1_io_out ? io_r_121_b : _GEN_510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_512 = 9'h7a == r_count_1_io_out ? io_r_122_b : _GEN_511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_513 = 9'h7b == r_count_1_io_out ? io_r_123_b : _GEN_512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_514 = 9'h7c == r_count_1_io_out ? io_r_124_b : _GEN_513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_515 = 9'h7d == r_count_1_io_out ? io_r_125_b : _GEN_514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_516 = 9'h7e == r_count_1_io_out ? io_r_126_b : _GEN_515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_517 = 9'h7f == r_count_1_io_out ? io_r_127_b : _GEN_516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_518 = 9'h80 == r_count_1_io_out ? io_r_128_b : _GEN_517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_519 = 9'h81 == r_count_1_io_out ? io_r_129_b : _GEN_518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_520 = 9'h82 == r_count_1_io_out ? io_r_130_b : _GEN_519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_521 = 9'h83 == r_count_1_io_out ? io_r_131_b : _GEN_520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_522 = 9'h84 == r_count_1_io_out ? io_r_132_b : _GEN_521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_523 = 9'h85 == r_count_1_io_out ? io_r_133_b : _GEN_522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_524 = 9'h86 == r_count_1_io_out ? io_r_134_b : _GEN_523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_525 = 9'h87 == r_count_1_io_out ? io_r_135_b : _GEN_524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_526 = 9'h88 == r_count_1_io_out ? io_r_136_b : _GEN_525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_527 = 9'h89 == r_count_1_io_out ? io_r_137_b : _GEN_526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_528 = 9'h8a == r_count_1_io_out ? io_r_138_b : _GEN_527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_529 = 9'h8b == r_count_1_io_out ? io_r_139_b : _GEN_528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_530 = 9'h8c == r_count_1_io_out ? io_r_140_b : _GEN_529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_531 = 9'h8d == r_count_1_io_out ? io_r_141_b : _GEN_530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_532 = 9'h8e == r_count_1_io_out ? io_r_142_b : _GEN_531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_533 = 9'h8f == r_count_1_io_out ? io_r_143_b : _GEN_532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_534 = 9'h90 == r_count_1_io_out ? io_r_144_b : _GEN_533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_535 = 9'h91 == r_count_1_io_out ? io_r_145_b : _GEN_534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_536 = 9'h92 == r_count_1_io_out ? io_r_146_b : _GEN_535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_537 = 9'h93 == r_count_1_io_out ? io_r_147_b : _GEN_536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_538 = 9'h94 == r_count_1_io_out ? io_r_148_b : _GEN_537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_539 = 9'h95 == r_count_1_io_out ? io_r_149_b : _GEN_538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_540 = 9'h96 == r_count_1_io_out ? io_r_150_b : _GEN_539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_541 = 9'h97 == r_count_1_io_out ? io_r_151_b : _GEN_540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_542 = 9'h98 == r_count_1_io_out ? io_r_152_b : _GEN_541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_543 = 9'h99 == r_count_1_io_out ? io_r_153_b : _GEN_542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_544 = 9'h9a == r_count_1_io_out ? io_r_154_b : _GEN_543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_545 = 9'h9b == r_count_1_io_out ? io_r_155_b : _GEN_544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_546 = 9'h9c == r_count_1_io_out ? io_r_156_b : _GEN_545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_547 = 9'h9d == r_count_1_io_out ? io_r_157_b : _GEN_546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_548 = 9'h9e == r_count_1_io_out ? io_r_158_b : _GEN_547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_549 = 9'h9f == r_count_1_io_out ? io_r_159_b : _GEN_548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_550 = 9'ha0 == r_count_1_io_out ? io_r_160_b : _GEN_549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_551 = 9'ha1 == r_count_1_io_out ? io_r_161_b : _GEN_550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_552 = 9'ha2 == r_count_1_io_out ? io_r_162_b : _GEN_551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_553 = 9'ha3 == r_count_1_io_out ? io_r_163_b : _GEN_552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_554 = 9'ha4 == r_count_1_io_out ? io_r_164_b : _GEN_553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_555 = 9'ha5 == r_count_1_io_out ? io_r_165_b : _GEN_554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_556 = 9'ha6 == r_count_1_io_out ? io_r_166_b : _GEN_555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_557 = 9'ha7 == r_count_1_io_out ? io_r_167_b : _GEN_556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_558 = 9'ha8 == r_count_1_io_out ? io_r_168_b : _GEN_557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_559 = 9'ha9 == r_count_1_io_out ? io_r_169_b : _GEN_558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_560 = 9'haa == r_count_1_io_out ? io_r_170_b : _GEN_559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_561 = 9'hab == r_count_1_io_out ? io_r_171_b : _GEN_560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_562 = 9'hac == r_count_1_io_out ? io_r_172_b : _GEN_561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_563 = 9'had == r_count_1_io_out ? io_r_173_b : _GEN_562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_564 = 9'hae == r_count_1_io_out ? io_r_174_b : _GEN_563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_565 = 9'haf == r_count_1_io_out ? io_r_175_b : _GEN_564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_566 = 9'hb0 == r_count_1_io_out ? io_r_176_b : _GEN_565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_567 = 9'hb1 == r_count_1_io_out ? io_r_177_b : _GEN_566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_568 = 9'hb2 == r_count_1_io_out ? io_r_178_b : _GEN_567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_569 = 9'hb3 == r_count_1_io_out ? io_r_179_b : _GEN_568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_570 = 9'hb4 == r_count_1_io_out ? io_r_180_b : _GEN_569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_571 = 9'hb5 == r_count_1_io_out ? io_r_181_b : _GEN_570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_572 = 9'hb6 == r_count_1_io_out ? io_r_182_b : _GEN_571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_573 = 9'hb7 == r_count_1_io_out ? io_r_183_b : _GEN_572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_574 = 9'hb8 == r_count_1_io_out ? io_r_184_b : _GEN_573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_575 = 9'hb9 == r_count_1_io_out ? io_r_185_b : _GEN_574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_576 = 9'hba == r_count_1_io_out ? io_r_186_b : _GEN_575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_577 = 9'hbb == r_count_1_io_out ? io_r_187_b : _GEN_576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_578 = 9'hbc == r_count_1_io_out ? io_r_188_b : _GEN_577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_579 = 9'hbd == r_count_1_io_out ? io_r_189_b : _GEN_578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_580 = 9'hbe == r_count_1_io_out ? io_r_190_b : _GEN_579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_581 = 9'hbf == r_count_1_io_out ? io_r_191_b : _GEN_580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_582 = 9'hc0 == r_count_1_io_out ? io_r_192_b : _GEN_581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_583 = 9'hc1 == r_count_1_io_out ? io_r_193_b : _GEN_582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_584 = 9'hc2 == r_count_1_io_out ? io_r_194_b : _GEN_583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_585 = 9'hc3 == r_count_1_io_out ? io_r_195_b : _GEN_584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_586 = 9'hc4 == r_count_1_io_out ? io_r_196_b : _GEN_585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_587 = 9'hc5 == r_count_1_io_out ? io_r_197_b : _GEN_586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_588 = 9'hc6 == r_count_1_io_out ? io_r_198_b : _GEN_587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_589 = 9'hc7 == r_count_1_io_out ? io_r_199_b : _GEN_588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_590 = 9'hc8 == r_count_1_io_out ? io_r_200_b : _GEN_589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_591 = 9'hc9 == r_count_1_io_out ? io_r_201_b : _GEN_590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_592 = 9'hca == r_count_1_io_out ? io_r_202_b : _GEN_591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_593 = 9'hcb == r_count_1_io_out ? io_r_203_b : _GEN_592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_594 = 9'hcc == r_count_1_io_out ? io_r_204_b : _GEN_593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_595 = 9'hcd == r_count_1_io_out ? io_r_205_b : _GEN_594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_596 = 9'hce == r_count_1_io_out ? io_r_206_b : _GEN_595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_597 = 9'hcf == r_count_1_io_out ? io_r_207_b : _GEN_596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_598 = 9'hd0 == r_count_1_io_out ? io_r_208_b : _GEN_597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_599 = 9'hd1 == r_count_1_io_out ? io_r_209_b : _GEN_598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_600 = 9'hd2 == r_count_1_io_out ? io_r_210_b : _GEN_599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_601 = 9'hd3 == r_count_1_io_out ? io_r_211_b : _GEN_600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_602 = 9'hd4 == r_count_1_io_out ? io_r_212_b : _GEN_601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_603 = 9'hd5 == r_count_1_io_out ? io_r_213_b : _GEN_602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_604 = 9'hd6 == r_count_1_io_out ? io_r_214_b : _GEN_603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_605 = 9'hd7 == r_count_1_io_out ? io_r_215_b : _GEN_604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_606 = 9'hd8 == r_count_1_io_out ? io_r_216_b : _GEN_605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_607 = 9'hd9 == r_count_1_io_out ? io_r_217_b : _GEN_606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_608 = 9'hda == r_count_1_io_out ? io_r_218_b : _GEN_607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_609 = 9'hdb == r_count_1_io_out ? io_r_219_b : _GEN_608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_610 = 9'hdc == r_count_1_io_out ? io_r_220_b : _GEN_609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_611 = 9'hdd == r_count_1_io_out ? io_r_221_b : _GEN_610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_612 = 9'hde == r_count_1_io_out ? io_r_222_b : _GEN_611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_613 = 9'hdf == r_count_1_io_out ? io_r_223_b : _GEN_612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_614 = 9'he0 == r_count_1_io_out ? io_r_224_b : _GEN_613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_615 = 9'he1 == r_count_1_io_out ? io_r_225_b : _GEN_614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_616 = 9'he2 == r_count_1_io_out ? io_r_226_b : _GEN_615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_617 = 9'he3 == r_count_1_io_out ? io_r_227_b : _GEN_616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_618 = 9'he4 == r_count_1_io_out ? io_r_228_b : _GEN_617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_619 = 9'he5 == r_count_1_io_out ? io_r_229_b : _GEN_618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_620 = 9'he6 == r_count_1_io_out ? io_r_230_b : _GEN_619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_621 = 9'he7 == r_count_1_io_out ? io_r_231_b : _GEN_620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_622 = 9'he8 == r_count_1_io_out ? io_r_232_b : _GEN_621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_623 = 9'he9 == r_count_1_io_out ? io_r_233_b : _GEN_622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_624 = 9'hea == r_count_1_io_out ? io_r_234_b : _GEN_623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_625 = 9'heb == r_count_1_io_out ? io_r_235_b : _GEN_624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_626 = 9'hec == r_count_1_io_out ? io_r_236_b : _GEN_625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_627 = 9'hed == r_count_1_io_out ? io_r_237_b : _GEN_626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_628 = 9'hee == r_count_1_io_out ? io_r_238_b : _GEN_627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_629 = 9'hef == r_count_1_io_out ? io_r_239_b : _GEN_628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_630 = 9'hf0 == r_count_1_io_out ? io_r_240_b : _GEN_629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_631 = 9'hf1 == r_count_1_io_out ? io_r_241_b : _GEN_630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_632 = 9'hf2 == r_count_1_io_out ? io_r_242_b : _GEN_631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_633 = 9'hf3 == r_count_1_io_out ? io_r_243_b : _GEN_632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_634 = 9'hf4 == r_count_1_io_out ? io_r_244_b : _GEN_633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_635 = 9'hf5 == r_count_1_io_out ? io_r_245_b : _GEN_634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_636 = 9'hf6 == r_count_1_io_out ? io_r_246_b : _GEN_635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_637 = 9'hf7 == r_count_1_io_out ? io_r_247_b : _GEN_636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_638 = 9'hf8 == r_count_1_io_out ? io_r_248_b : _GEN_637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_639 = 9'hf9 == r_count_1_io_out ? io_r_249_b : _GEN_638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_640 = 9'hfa == r_count_1_io_out ? io_r_250_b : _GEN_639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_641 = 9'hfb == r_count_1_io_out ? io_r_251_b : _GEN_640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_642 = 9'hfc == r_count_1_io_out ? io_r_252_b : _GEN_641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_643 = 9'hfd == r_count_1_io_out ? io_r_253_b : _GEN_642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_644 = 9'hfe == r_count_1_io_out ? io_r_254_b : _GEN_643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_645 = 9'hff == r_count_1_io_out ? io_r_255_b : _GEN_644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_646 = 9'h100 == r_count_1_io_out ? io_r_256_b : _GEN_645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_647 = 9'h101 == r_count_1_io_out ? io_r_257_b : _GEN_646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_648 = 9'h102 == r_count_1_io_out ? io_r_258_b : _GEN_647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_649 = 9'h103 == r_count_1_io_out ? io_r_259_b : _GEN_648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_650 = 9'h104 == r_count_1_io_out ? io_r_260_b : _GEN_649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_651 = 9'h105 == r_count_1_io_out ? io_r_261_b : _GEN_650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_652 = 9'h106 == r_count_1_io_out ? io_r_262_b : _GEN_651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_653 = 9'h107 == r_count_1_io_out ? io_r_263_b : _GEN_652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_654 = 9'h108 == r_count_1_io_out ? io_r_264_b : _GEN_653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_655 = 9'h109 == r_count_1_io_out ? io_r_265_b : _GEN_654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_656 = 9'h10a == r_count_1_io_out ? io_r_266_b : _GEN_655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_657 = 9'h10b == r_count_1_io_out ? io_r_267_b : _GEN_656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_658 = 9'h10c == r_count_1_io_out ? io_r_268_b : _GEN_657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_659 = 9'h10d == r_count_1_io_out ? io_r_269_b : _GEN_658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_660 = 9'h10e == r_count_1_io_out ? io_r_270_b : _GEN_659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_661 = 9'h10f == r_count_1_io_out ? io_r_271_b : _GEN_660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_662 = 9'h110 == r_count_1_io_out ? io_r_272_b : _GEN_661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_663 = 9'h111 == r_count_1_io_out ? io_r_273_b : _GEN_662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_664 = 9'h112 == r_count_1_io_out ? io_r_274_b : _GEN_663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_665 = 9'h113 == r_count_1_io_out ? io_r_275_b : _GEN_664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_666 = 9'h114 == r_count_1_io_out ? io_r_276_b : _GEN_665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_667 = 9'h115 == r_count_1_io_out ? io_r_277_b : _GEN_666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_668 = 9'h116 == r_count_1_io_out ? io_r_278_b : _GEN_667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_669 = 9'h117 == r_count_1_io_out ? io_r_279_b : _GEN_668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_670 = 9'h118 == r_count_1_io_out ? io_r_280_b : _GEN_669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_671 = 9'h119 == r_count_1_io_out ? io_r_281_b : _GEN_670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_672 = 9'h11a == r_count_1_io_out ? io_r_282_b : _GEN_671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_673 = 9'h11b == r_count_1_io_out ? io_r_283_b : _GEN_672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_674 = 9'h11c == r_count_1_io_out ? io_r_284_b : _GEN_673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_675 = 9'h11d == r_count_1_io_out ? io_r_285_b : _GEN_674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_676 = 9'h11e == r_count_1_io_out ? io_r_286_b : _GEN_675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_677 = 9'h11f == r_count_1_io_out ? io_r_287_b : _GEN_676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_678 = 9'h120 == r_count_1_io_out ? io_r_288_b : _GEN_677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_679 = 9'h121 == r_count_1_io_out ? io_r_289_b : _GEN_678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_680 = 9'h122 == r_count_1_io_out ? io_r_290_b : _GEN_679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_681 = 9'h123 == r_count_1_io_out ? io_r_291_b : _GEN_680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_682 = 9'h124 == r_count_1_io_out ? io_r_292_b : _GEN_681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_683 = 9'h125 == r_count_1_io_out ? io_r_293_b : _GEN_682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_684 = 9'h126 == r_count_1_io_out ? io_r_294_b : _GEN_683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_685 = 9'h127 == r_count_1_io_out ? io_r_295_b : _GEN_684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_686 = 9'h128 == r_count_1_io_out ? io_r_296_b : _GEN_685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_687 = 9'h129 == r_count_1_io_out ? io_r_297_b : _GEN_686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_688 = 9'h12a == r_count_1_io_out ? io_r_298_b : _GEN_687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_691 = 9'h1 == r_count_2_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_692 = 9'h2 == r_count_2_io_out ? io_r_2_b : _GEN_691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_693 = 9'h3 == r_count_2_io_out ? io_r_3_b : _GEN_692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_694 = 9'h4 == r_count_2_io_out ? io_r_4_b : _GEN_693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_695 = 9'h5 == r_count_2_io_out ? io_r_5_b : _GEN_694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_696 = 9'h6 == r_count_2_io_out ? io_r_6_b : _GEN_695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_697 = 9'h7 == r_count_2_io_out ? io_r_7_b : _GEN_696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_698 = 9'h8 == r_count_2_io_out ? io_r_8_b : _GEN_697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_699 = 9'h9 == r_count_2_io_out ? io_r_9_b : _GEN_698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_700 = 9'ha == r_count_2_io_out ? io_r_10_b : _GEN_699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_701 = 9'hb == r_count_2_io_out ? io_r_11_b : _GEN_700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_702 = 9'hc == r_count_2_io_out ? io_r_12_b : _GEN_701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_703 = 9'hd == r_count_2_io_out ? io_r_13_b : _GEN_702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_704 = 9'he == r_count_2_io_out ? io_r_14_b : _GEN_703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_705 = 9'hf == r_count_2_io_out ? io_r_15_b : _GEN_704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_706 = 9'h10 == r_count_2_io_out ? io_r_16_b : _GEN_705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_707 = 9'h11 == r_count_2_io_out ? io_r_17_b : _GEN_706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_708 = 9'h12 == r_count_2_io_out ? io_r_18_b : _GEN_707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_709 = 9'h13 == r_count_2_io_out ? io_r_19_b : _GEN_708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_710 = 9'h14 == r_count_2_io_out ? io_r_20_b : _GEN_709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_711 = 9'h15 == r_count_2_io_out ? io_r_21_b : _GEN_710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_712 = 9'h16 == r_count_2_io_out ? io_r_22_b : _GEN_711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_713 = 9'h17 == r_count_2_io_out ? io_r_23_b : _GEN_712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_714 = 9'h18 == r_count_2_io_out ? io_r_24_b : _GEN_713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_715 = 9'h19 == r_count_2_io_out ? io_r_25_b : _GEN_714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_716 = 9'h1a == r_count_2_io_out ? io_r_26_b : _GEN_715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_717 = 9'h1b == r_count_2_io_out ? io_r_27_b : _GEN_716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_718 = 9'h1c == r_count_2_io_out ? io_r_28_b : _GEN_717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_719 = 9'h1d == r_count_2_io_out ? io_r_29_b : _GEN_718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_720 = 9'h1e == r_count_2_io_out ? io_r_30_b : _GEN_719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_721 = 9'h1f == r_count_2_io_out ? io_r_31_b : _GEN_720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_722 = 9'h20 == r_count_2_io_out ? io_r_32_b : _GEN_721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_723 = 9'h21 == r_count_2_io_out ? io_r_33_b : _GEN_722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_724 = 9'h22 == r_count_2_io_out ? io_r_34_b : _GEN_723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_725 = 9'h23 == r_count_2_io_out ? io_r_35_b : _GEN_724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_726 = 9'h24 == r_count_2_io_out ? io_r_36_b : _GEN_725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_727 = 9'h25 == r_count_2_io_out ? io_r_37_b : _GEN_726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_728 = 9'h26 == r_count_2_io_out ? io_r_38_b : _GEN_727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_729 = 9'h27 == r_count_2_io_out ? io_r_39_b : _GEN_728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_730 = 9'h28 == r_count_2_io_out ? io_r_40_b : _GEN_729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_731 = 9'h29 == r_count_2_io_out ? io_r_41_b : _GEN_730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_732 = 9'h2a == r_count_2_io_out ? io_r_42_b : _GEN_731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_733 = 9'h2b == r_count_2_io_out ? io_r_43_b : _GEN_732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_734 = 9'h2c == r_count_2_io_out ? io_r_44_b : _GEN_733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_735 = 9'h2d == r_count_2_io_out ? io_r_45_b : _GEN_734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_736 = 9'h2e == r_count_2_io_out ? io_r_46_b : _GEN_735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_737 = 9'h2f == r_count_2_io_out ? io_r_47_b : _GEN_736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_738 = 9'h30 == r_count_2_io_out ? io_r_48_b : _GEN_737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_739 = 9'h31 == r_count_2_io_out ? io_r_49_b : _GEN_738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_740 = 9'h32 == r_count_2_io_out ? io_r_50_b : _GEN_739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_741 = 9'h33 == r_count_2_io_out ? io_r_51_b : _GEN_740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_742 = 9'h34 == r_count_2_io_out ? io_r_52_b : _GEN_741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_743 = 9'h35 == r_count_2_io_out ? io_r_53_b : _GEN_742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_744 = 9'h36 == r_count_2_io_out ? io_r_54_b : _GEN_743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_745 = 9'h37 == r_count_2_io_out ? io_r_55_b : _GEN_744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_746 = 9'h38 == r_count_2_io_out ? io_r_56_b : _GEN_745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_747 = 9'h39 == r_count_2_io_out ? io_r_57_b : _GEN_746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_748 = 9'h3a == r_count_2_io_out ? io_r_58_b : _GEN_747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_749 = 9'h3b == r_count_2_io_out ? io_r_59_b : _GEN_748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_750 = 9'h3c == r_count_2_io_out ? io_r_60_b : _GEN_749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_751 = 9'h3d == r_count_2_io_out ? io_r_61_b : _GEN_750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_752 = 9'h3e == r_count_2_io_out ? io_r_62_b : _GEN_751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_753 = 9'h3f == r_count_2_io_out ? io_r_63_b : _GEN_752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_754 = 9'h40 == r_count_2_io_out ? io_r_64_b : _GEN_753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_755 = 9'h41 == r_count_2_io_out ? io_r_65_b : _GEN_754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_756 = 9'h42 == r_count_2_io_out ? io_r_66_b : _GEN_755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_757 = 9'h43 == r_count_2_io_out ? io_r_67_b : _GEN_756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_758 = 9'h44 == r_count_2_io_out ? io_r_68_b : _GEN_757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_759 = 9'h45 == r_count_2_io_out ? io_r_69_b : _GEN_758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_760 = 9'h46 == r_count_2_io_out ? io_r_70_b : _GEN_759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_761 = 9'h47 == r_count_2_io_out ? io_r_71_b : _GEN_760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_762 = 9'h48 == r_count_2_io_out ? io_r_72_b : _GEN_761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_763 = 9'h49 == r_count_2_io_out ? io_r_73_b : _GEN_762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_764 = 9'h4a == r_count_2_io_out ? io_r_74_b : _GEN_763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_765 = 9'h4b == r_count_2_io_out ? io_r_75_b : _GEN_764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_766 = 9'h4c == r_count_2_io_out ? io_r_76_b : _GEN_765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_767 = 9'h4d == r_count_2_io_out ? io_r_77_b : _GEN_766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_768 = 9'h4e == r_count_2_io_out ? io_r_78_b : _GEN_767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_769 = 9'h4f == r_count_2_io_out ? io_r_79_b : _GEN_768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_770 = 9'h50 == r_count_2_io_out ? io_r_80_b : _GEN_769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_771 = 9'h51 == r_count_2_io_out ? io_r_81_b : _GEN_770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_772 = 9'h52 == r_count_2_io_out ? io_r_82_b : _GEN_771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_773 = 9'h53 == r_count_2_io_out ? io_r_83_b : _GEN_772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_774 = 9'h54 == r_count_2_io_out ? io_r_84_b : _GEN_773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_775 = 9'h55 == r_count_2_io_out ? io_r_85_b : _GEN_774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_776 = 9'h56 == r_count_2_io_out ? io_r_86_b : _GEN_775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_777 = 9'h57 == r_count_2_io_out ? io_r_87_b : _GEN_776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_778 = 9'h58 == r_count_2_io_out ? io_r_88_b : _GEN_777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_779 = 9'h59 == r_count_2_io_out ? io_r_89_b : _GEN_778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_780 = 9'h5a == r_count_2_io_out ? io_r_90_b : _GEN_779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_781 = 9'h5b == r_count_2_io_out ? io_r_91_b : _GEN_780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_782 = 9'h5c == r_count_2_io_out ? io_r_92_b : _GEN_781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_783 = 9'h5d == r_count_2_io_out ? io_r_93_b : _GEN_782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_784 = 9'h5e == r_count_2_io_out ? io_r_94_b : _GEN_783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_785 = 9'h5f == r_count_2_io_out ? io_r_95_b : _GEN_784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_786 = 9'h60 == r_count_2_io_out ? io_r_96_b : _GEN_785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_787 = 9'h61 == r_count_2_io_out ? io_r_97_b : _GEN_786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_788 = 9'h62 == r_count_2_io_out ? io_r_98_b : _GEN_787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_789 = 9'h63 == r_count_2_io_out ? io_r_99_b : _GEN_788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_790 = 9'h64 == r_count_2_io_out ? io_r_100_b : _GEN_789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_791 = 9'h65 == r_count_2_io_out ? io_r_101_b : _GEN_790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_792 = 9'h66 == r_count_2_io_out ? io_r_102_b : _GEN_791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_793 = 9'h67 == r_count_2_io_out ? io_r_103_b : _GEN_792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_794 = 9'h68 == r_count_2_io_out ? io_r_104_b : _GEN_793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_795 = 9'h69 == r_count_2_io_out ? io_r_105_b : _GEN_794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_796 = 9'h6a == r_count_2_io_out ? io_r_106_b : _GEN_795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_797 = 9'h6b == r_count_2_io_out ? io_r_107_b : _GEN_796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_798 = 9'h6c == r_count_2_io_out ? io_r_108_b : _GEN_797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_799 = 9'h6d == r_count_2_io_out ? io_r_109_b : _GEN_798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_800 = 9'h6e == r_count_2_io_out ? io_r_110_b : _GEN_799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_801 = 9'h6f == r_count_2_io_out ? io_r_111_b : _GEN_800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_802 = 9'h70 == r_count_2_io_out ? io_r_112_b : _GEN_801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_803 = 9'h71 == r_count_2_io_out ? io_r_113_b : _GEN_802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_804 = 9'h72 == r_count_2_io_out ? io_r_114_b : _GEN_803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_805 = 9'h73 == r_count_2_io_out ? io_r_115_b : _GEN_804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_806 = 9'h74 == r_count_2_io_out ? io_r_116_b : _GEN_805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_807 = 9'h75 == r_count_2_io_out ? io_r_117_b : _GEN_806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_808 = 9'h76 == r_count_2_io_out ? io_r_118_b : _GEN_807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_809 = 9'h77 == r_count_2_io_out ? io_r_119_b : _GEN_808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_810 = 9'h78 == r_count_2_io_out ? io_r_120_b : _GEN_809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_811 = 9'h79 == r_count_2_io_out ? io_r_121_b : _GEN_810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_812 = 9'h7a == r_count_2_io_out ? io_r_122_b : _GEN_811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_813 = 9'h7b == r_count_2_io_out ? io_r_123_b : _GEN_812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_814 = 9'h7c == r_count_2_io_out ? io_r_124_b : _GEN_813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_815 = 9'h7d == r_count_2_io_out ? io_r_125_b : _GEN_814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_816 = 9'h7e == r_count_2_io_out ? io_r_126_b : _GEN_815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_817 = 9'h7f == r_count_2_io_out ? io_r_127_b : _GEN_816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_818 = 9'h80 == r_count_2_io_out ? io_r_128_b : _GEN_817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_819 = 9'h81 == r_count_2_io_out ? io_r_129_b : _GEN_818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_820 = 9'h82 == r_count_2_io_out ? io_r_130_b : _GEN_819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_821 = 9'h83 == r_count_2_io_out ? io_r_131_b : _GEN_820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_822 = 9'h84 == r_count_2_io_out ? io_r_132_b : _GEN_821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_823 = 9'h85 == r_count_2_io_out ? io_r_133_b : _GEN_822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_824 = 9'h86 == r_count_2_io_out ? io_r_134_b : _GEN_823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_825 = 9'h87 == r_count_2_io_out ? io_r_135_b : _GEN_824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_826 = 9'h88 == r_count_2_io_out ? io_r_136_b : _GEN_825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_827 = 9'h89 == r_count_2_io_out ? io_r_137_b : _GEN_826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_828 = 9'h8a == r_count_2_io_out ? io_r_138_b : _GEN_827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_829 = 9'h8b == r_count_2_io_out ? io_r_139_b : _GEN_828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_830 = 9'h8c == r_count_2_io_out ? io_r_140_b : _GEN_829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_831 = 9'h8d == r_count_2_io_out ? io_r_141_b : _GEN_830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_832 = 9'h8e == r_count_2_io_out ? io_r_142_b : _GEN_831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_833 = 9'h8f == r_count_2_io_out ? io_r_143_b : _GEN_832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_834 = 9'h90 == r_count_2_io_out ? io_r_144_b : _GEN_833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_835 = 9'h91 == r_count_2_io_out ? io_r_145_b : _GEN_834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_836 = 9'h92 == r_count_2_io_out ? io_r_146_b : _GEN_835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_837 = 9'h93 == r_count_2_io_out ? io_r_147_b : _GEN_836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_838 = 9'h94 == r_count_2_io_out ? io_r_148_b : _GEN_837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_839 = 9'h95 == r_count_2_io_out ? io_r_149_b : _GEN_838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_840 = 9'h96 == r_count_2_io_out ? io_r_150_b : _GEN_839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_841 = 9'h97 == r_count_2_io_out ? io_r_151_b : _GEN_840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_842 = 9'h98 == r_count_2_io_out ? io_r_152_b : _GEN_841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_843 = 9'h99 == r_count_2_io_out ? io_r_153_b : _GEN_842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_844 = 9'h9a == r_count_2_io_out ? io_r_154_b : _GEN_843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_845 = 9'h9b == r_count_2_io_out ? io_r_155_b : _GEN_844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_846 = 9'h9c == r_count_2_io_out ? io_r_156_b : _GEN_845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_847 = 9'h9d == r_count_2_io_out ? io_r_157_b : _GEN_846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_848 = 9'h9e == r_count_2_io_out ? io_r_158_b : _GEN_847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_849 = 9'h9f == r_count_2_io_out ? io_r_159_b : _GEN_848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_850 = 9'ha0 == r_count_2_io_out ? io_r_160_b : _GEN_849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_851 = 9'ha1 == r_count_2_io_out ? io_r_161_b : _GEN_850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_852 = 9'ha2 == r_count_2_io_out ? io_r_162_b : _GEN_851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_853 = 9'ha3 == r_count_2_io_out ? io_r_163_b : _GEN_852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_854 = 9'ha4 == r_count_2_io_out ? io_r_164_b : _GEN_853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_855 = 9'ha5 == r_count_2_io_out ? io_r_165_b : _GEN_854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_856 = 9'ha6 == r_count_2_io_out ? io_r_166_b : _GEN_855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_857 = 9'ha7 == r_count_2_io_out ? io_r_167_b : _GEN_856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_858 = 9'ha8 == r_count_2_io_out ? io_r_168_b : _GEN_857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_859 = 9'ha9 == r_count_2_io_out ? io_r_169_b : _GEN_858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_860 = 9'haa == r_count_2_io_out ? io_r_170_b : _GEN_859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_861 = 9'hab == r_count_2_io_out ? io_r_171_b : _GEN_860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_862 = 9'hac == r_count_2_io_out ? io_r_172_b : _GEN_861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_863 = 9'had == r_count_2_io_out ? io_r_173_b : _GEN_862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_864 = 9'hae == r_count_2_io_out ? io_r_174_b : _GEN_863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_865 = 9'haf == r_count_2_io_out ? io_r_175_b : _GEN_864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_866 = 9'hb0 == r_count_2_io_out ? io_r_176_b : _GEN_865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_867 = 9'hb1 == r_count_2_io_out ? io_r_177_b : _GEN_866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_868 = 9'hb2 == r_count_2_io_out ? io_r_178_b : _GEN_867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_869 = 9'hb3 == r_count_2_io_out ? io_r_179_b : _GEN_868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_870 = 9'hb4 == r_count_2_io_out ? io_r_180_b : _GEN_869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_871 = 9'hb5 == r_count_2_io_out ? io_r_181_b : _GEN_870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_872 = 9'hb6 == r_count_2_io_out ? io_r_182_b : _GEN_871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_873 = 9'hb7 == r_count_2_io_out ? io_r_183_b : _GEN_872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_874 = 9'hb8 == r_count_2_io_out ? io_r_184_b : _GEN_873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_875 = 9'hb9 == r_count_2_io_out ? io_r_185_b : _GEN_874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_876 = 9'hba == r_count_2_io_out ? io_r_186_b : _GEN_875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_877 = 9'hbb == r_count_2_io_out ? io_r_187_b : _GEN_876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_878 = 9'hbc == r_count_2_io_out ? io_r_188_b : _GEN_877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_879 = 9'hbd == r_count_2_io_out ? io_r_189_b : _GEN_878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_880 = 9'hbe == r_count_2_io_out ? io_r_190_b : _GEN_879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_881 = 9'hbf == r_count_2_io_out ? io_r_191_b : _GEN_880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_882 = 9'hc0 == r_count_2_io_out ? io_r_192_b : _GEN_881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_883 = 9'hc1 == r_count_2_io_out ? io_r_193_b : _GEN_882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_884 = 9'hc2 == r_count_2_io_out ? io_r_194_b : _GEN_883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_885 = 9'hc3 == r_count_2_io_out ? io_r_195_b : _GEN_884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_886 = 9'hc4 == r_count_2_io_out ? io_r_196_b : _GEN_885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_887 = 9'hc5 == r_count_2_io_out ? io_r_197_b : _GEN_886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_888 = 9'hc6 == r_count_2_io_out ? io_r_198_b : _GEN_887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_889 = 9'hc7 == r_count_2_io_out ? io_r_199_b : _GEN_888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_890 = 9'hc8 == r_count_2_io_out ? io_r_200_b : _GEN_889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_891 = 9'hc9 == r_count_2_io_out ? io_r_201_b : _GEN_890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_892 = 9'hca == r_count_2_io_out ? io_r_202_b : _GEN_891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_893 = 9'hcb == r_count_2_io_out ? io_r_203_b : _GEN_892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_894 = 9'hcc == r_count_2_io_out ? io_r_204_b : _GEN_893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_895 = 9'hcd == r_count_2_io_out ? io_r_205_b : _GEN_894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_896 = 9'hce == r_count_2_io_out ? io_r_206_b : _GEN_895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_897 = 9'hcf == r_count_2_io_out ? io_r_207_b : _GEN_896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_898 = 9'hd0 == r_count_2_io_out ? io_r_208_b : _GEN_897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_899 = 9'hd1 == r_count_2_io_out ? io_r_209_b : _GEN_898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_900 = 9'hd2 == r_count_2_io_out ? io_r_210_b : _GEN_899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_901 = 9'hd3 == r_count_2_io_out ? io_r_211_b : _GEN_900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_902 = 9'hd4 == r_count_2_io_out ? io_r_212_b : _GEN_901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_903 = 9'hd5 == r_count_2_io_out ? io_r_213_b : _GEN_902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_904 = 9'hd6 == r_count_2_io_out ? io_r_214_b : _GEN_903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_905 = 9'hd7 == r_count_2_io_out ? io_r_215_b : _GEN_904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_906 = 9'hd8 == r_count_2_io_out ? io_r_216_b : _GEN_905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_907 = 9'hd9 == r_count_2_io_out ? io_r_217_b : _GEN_906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_908 = 9'hda == r_count_2_io_out ? io_r_218_b : _GEN_907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_909 = 9'hdb == r_count_2_io_out ? io_r_219_b : _GEN_908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_910 = 9'hdc == r_count_2_io_out ? io_r_220_b : _GEN_909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_911 = 9'hdd == r_count_2_io_out ? io_r_221_b : _GEN_910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_912 = 9'hde == r_count_2_io_out ? io_r_222_b : _GEN_911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_913 = 9'hdf == r_count_2_io_out ? io_r_223_b : _GEN_912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_914 = 9'he0 == r_count_2_io_out ? io_r_224_b : _GEN_913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_915 = 9'he1 == r_count_2_io_out ? io_r_225_b : _GEN_914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_916 = 9'he2 == r_count_2_io_out ? io_r_226_b : _GEN_915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_917 = 9'he3 == r_count_2_io_out ? io_r_227_b : _GEN_916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_918 = 9'he4 == r_count_2_io_out ? io_r_228_b : _GEN_917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_919 = 9'he5 == r_count_2_io_out ? io_r_229_b : _GEN_918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_920 = 9'he6 == r_count_2_io_out ? io_r_230_b : _GEN_919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_921 = 9'he7 == r_count_2_io_out ? io_r_231_b : _GEN_920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_922 = 9'he8 == r_count_2_io_out ? io_r_232_b : _GEN_921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_923 = 9'he9 == r_count_2_io_out ? io_r_233_b : _GEN_922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_924 = 9'hea == r_count_2_io_out ? io_r_234_b : _GEN_923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_925 = 9'heb == r_count_2_io_out ? io_r_235_b : _GEN_924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_926 = 9'hec == r_count_2_io_out ? io_r_236_b : _GEN_925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_927 = 9'hed == r_count_2_io_out ? io_r_237_b : _GEN_926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_928 = 9'hee == r_count_2_io_out ? io_r_238_b : _GEN_927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_929 = 9'hef == r_count_2_io_out ? io_r_239_b : _GEN_928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_930 = 9'hf0 == r_count_2_io_out ? io_r_240_b : _GEN_929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_931 = 9'hf1 == r_count_2_io_out ? io_r_241_b : _GEN_930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_932 = 9'hf2 == r_count_2_io_out ? io_r_242_b : _GEN_931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_933 = 9'hf3 == r_count_2_io_out ? io_r_243_b : _GEN_932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_934 = 9'hf4 == r_count_2_io_out ? io_r_244_b : _GEN_933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_935 = 9'hf5 == r_count_2_io_out ? io_r_245_b : _GEN_934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_936 = 9'hf6 == r_count_2_io_out ? io_r_246_b : _GEN_935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_937 = 9'hf7 == r_count_2_io_out ? io_r_247_b : _GEN_936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_938 = 9'hf8 == r_count_2_io_out ? io_r_248_b : _GEN_937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_939 = 9'hf9 == r_count_2_io_out ? io_r_249_b : _GEN_938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_940 = 9'hfa == r_count_2_io_out ? io_r_250_b : _GEN_939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_941 = 9'hfb == r_count_2_io_out ? io_r_251_b : _GEN_940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_942 = 9'hfc == r_count_2_io_out ? io_r_252_b : _GEN_941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_943 = 9'hfd == r_count_2_io_out ? io_r_253_b : _GEN_942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_944 = 9'hfe == r_count_2_io_out ? io_r_254_b : _GEN_943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_945 = 9'hff == r_count_2_io_out ? io_r_255_b : _GEN_944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_946 = 9'h100 == r_count_2_io_out ? io_r_256_b : _GEN_945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_947 = 9'h101 == r_count_2_io_out ? io_r_257_b : _GEN_946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_948 = 9'h102 == r_count_2_io_out ? io_r_258_b : _GEN_947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_949 = 9'h103 == r_count_2_io_out ? io_r_259_b : _GEN_948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_950 = 9'h104 == r_count_2_io_out ? io_r_260_b : _GEN_949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_951 = 9'h105 == r_count_2_io_out ? io_r_261_b : _GEN_950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_952 = 9'h106 == r_count_2_io_out ? io_r_262_b : _GEN_951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_953 = 9'h107 == r_count_2_io_out ? io_r_263_b : _GEN_952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_954 = 9'h108 == r_count_2_io_out ? io_r_264_b : _GEN_953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_955 = 9'h109 == r_count_2_io_out ? io_r_265_b : _GEN_954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_956 = 9'h10a == r_count_2_io_out ? io_r_266_b : _GEN_955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_957 = 9'h10b == r_count_2_io_out ? io_r_267_b : _GEN_956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_958 = 9'h10c == r_count_2_io_out ? io_r_268_b : _GEN_957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_959 = 9'h10d == r_count_2_io_out ? io_r_269_b : _GEN_958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_960 = 9'h10e == r_count_2_io_out ? io_r_270_b : _GEN_959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_961 = 9'h10f == r_count_2_io_out ? io_r_271_b : _GEN_960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_962 = 9'h110 == r_count_2_io_out ? io_r_272_b : _GEN_961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_963 = 9'h111 == r_count_2_io_out ? io_r_273_b : _GEN_962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_964 = 9'h112 == r_count_2_io_out ? io_r_274_b : _GEN_963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_965 = 9'h113 == r_count_2_io_out ? io_r_275_b : _GEN_964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_966 = 9'h114 == r_count_2_io_out ? io_r_276_b : _GEN_965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_967 = 9'h115 == r_count_2_io_out ? io_r_277_b : _GEN_966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_968 = 9'h116 == r_count_2_io_out ? io_r_278_b : _GEN_967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_969 = 9'h117 == r_count_2_io_out ? io_r_279_b : _GEN_968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_970 = 9'h118 == r_count_2_io_out ? io_r_280_b : _GEN_969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_971 = 9'h119 == r_count_2_io_out ? io_r_281_b : _GEN_970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_972 = 9'h11a == r_count_2_io_out ? io_r_282_b : _GEN_971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_973 = 9'h11b == r_count_2_io_out ? io_r_283_b : _GEN_972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_974 = 9'h11c == r_count_2_io_out ? io_r_284_b : _GEN_973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_975 = 9'h11d == r_count_2_io_out ? io_r_285_b : _GEN_974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_976 = 9'h11e == r_count_2_io_out ? io_r_286_b : _GEN_975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_977 = 9'h11f == r_count_2_io_out ? io_r_287_b : _GEN_976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_978 = 9'h120 == r_count_2_io_out ? io_r_288_b : _GEN_977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_979 = 9'h121 == r_count_2_io_out ? io_r_289_b : _GEN_978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_980 = 9'h122 == r_count_2_io_out ? io_r_290_b : _GEN_979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_981 = 9'h123 == r_count_2_io_out ? io_r_291_b : _GEN_980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_982 = 9'h124 == r_count_2_io_out ? io_r_292_b : _GEN_981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_983 = 9'h125 == r_count_2_io_out ? io_r_293_b : _GEN_982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_984 = 9'h126 == r_count_2_io_out ? io_r_294_b : _GEN_983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_985 = 9'h127 == r_count_2_io_out ? io_r_295_b : _GEN_984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_986 = 9'h128 == r_count_2_io_out ? io_r_296_b : _GEN_985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_987 = 9'h129 == r_count_2_io_out ? io_r_297_b : _GEN_986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_988 = 9'h12a == r_count_2_io_out ? io_r_298_b : _GEN_987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_991 = 9'h1 == r_count_3_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_992 = 9'h2 == r_count_3_io_out ? io_r_2_b : _GEN_991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_993 = 9'h3 == r_count_3_io_out ? io_r_3_b : _GEN_992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_994 = 9'h4 == r_count_3_io_out ? io_r_4_b : _GEN_993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_995 = 9'h5 == r_count_3_io_out ? io_r_5_b : _GEN_994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_996 = 9'h6 == r_count_3_io_out ? io_r_6_b : _GEN_995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_997 = 9'h7 == r_count_3_io_out ? io_r_7_b : _GEN_996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_998 = 9'h8 == r_count_3_io_out ? io_r_8_b : _GEN_997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_999 = 9'h9 == r_count_3_io_out ? io_r_9_b : _GEN_998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1000 = 9'ha == r_count_3_io_out ? io_r_10_b : _GEN_999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1001 = 9'hb == r_count_3_io_out ? io_r_11_b : _GEN_1000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1002 = 9'hc == r_count_3_io_out ? io_r_12_b : _GEN_1001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1003 = 9'hd == r_count_3_io_out ? io_r_13_b : _GEN_1002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1004 = 9'he == r_count_3_io_out ? io_r_14_b : _GEN_1003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1005 = 9'hf == r_count_3_io_out ? io_r_15_b : _GEN_1004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1006 = 9'h10 == r_count_3_io_out ? io_r_16_b : _GEN_1005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1007 = 9'h11 == r_count_3_io_out ? io_r_17_b : _GEN_1006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1008 = 9'h12 == r_count_3_io_out ? io_r_18_b : _GEN_1007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1009 = 9'h13 == r_count_3_io_out ? io_r_19_b : _GEN_1008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1010 = 9'h14 == r_count_3_io_out ? io_r_20_b : _GEN_1009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1011 = 9'h15 == r_count_3_io_out ? io_r_21_b : _GEN_1010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1012 = 9'h16 == r_count_3_io_out ? io_r_22_b : _GEN_1011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1013 = 9'h17 == r_count_3_io_out ? io_r_23_b : _GEN_1012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1014 = 9'h18 == r_count_3_io_out ? io_r_24_b : _GEN_1013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1015 = 9'h19 == r_count_3_io_out ? io_r_25_b : _GEN_1014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1016 = 9'h1a == r_count_3_io_out ? io_r_26_b : _GEN_1015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1017 = 9'h1b == r_count_3_io_out ? io_r_27_b : _GEN_1016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1018 = 9'h1c == r_count_3_io_out ? io_r_28_b : _GEN_1017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1019 = 9'h1d == r_count_3_io_out ? io_r_29_b : _GEN_1018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1020 = 9'h1e == r_count_3_io_out ? io_r_30_b : _GEN_1019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1021 = 9'h1f == r_count_3_io_out ? io_r_31_b : _GEN_1020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1022 = 9'h20 == r_count_3_io_out ? io_r_32_b : _GEN_1021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1023 = 9'h21 == r_count_3_io_out ? io_r_33_b : _GEN_1022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1024 = 9'h22 == r_count_3_io_out ? io_r_34_b : _GEN_1023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1025 = 9'h23 == r_count_3_io_out ? io_r_35_b : _GEN_1024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1026 = 9'h24 == r_count_3_io_out ? io_r_36_b : _GEN_1025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1027 = 9'h25 == r_count_3_io_out ? io_r_37_b : _GEN_1026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1028 = 9'h26 == r_count_3_io_out ? io_r_38_b : _GEN_1027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1029 = 9'h27 == r_count_3_io_out ? io_r_39_b : _GEN_1028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1030 = 9'h28 == r_count_3_io_out ? io_r_40_b : _GEN_1029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1031 = 9'h29 == r_count_3_io_out ? io_r_41_b : _GEN_1030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1032 = 9'h2a == r_count_3_io_out ? io_r_42_b : _GEN_1031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1033 = 9'h2b == r_count_3_io_out ? io_r_43_b : _GEN_1032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1034 = 9'h2c == r_count_3_io_out ? io_r_44_b : _GEN_1033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1035 = 9'h2d == r_count_3_io_out ? io_r_45_b : _GEN_1034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1036 = 9'h2e == r_count_3_io_out ? io_r_46_b : _GEN_1035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1037 = 9'h2f == r_count_3_io_out ? io_r_47_b : _GEN_1036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1038 = 9'h30 == r_count_3_io_out ? io_r_48_b : _GEN_1037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1039 = 9'h31 == r_count_3_io_out ? io_r_49_b : _GEN_1038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1040 = 9'h32 == r_count_3_io_out ? io_r_50_b : _GEN_1039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1041 = 9'h33 == r_count_3_io_out ? io_r_51_b : _GEN_1040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1042 = 9'h34 == r_count_3_io_out ? io_r_52_b : _GEN_1041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1043 = 9'h35 == r_count_3_io_out ? io_r_53_b : _GEN_1042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1044 = 9'h36 == r_count_3_io_out ? io_r_54_b : _GEN_1043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1045 = 9'h37 == r_count_3_io_out ? io_r_55_b : _GEN_1044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1046 = 9'h38 == r_count_3_io_out ? io_r_56_b : _GEN_1045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1047 = 9'h39 == r_count_3_io_out ? io_r_57_b : _GEN_1046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1048 = 9'h3a == r_count_3_io_out ? io_r_58_b : _GEN_1047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1049 = 9'h3b == r_count_3_io_out ? io_r_59_b : _GEN_1048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1050 = 9'h3c == r_count_3_io_out ? io_r_60_b : _GEN_1049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1051 = 9'h3d == r_count_3_io_out ? io_r_61_b : _GEN_1050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1052 = 9'h3e == r_count_3_io_out ? io_r_62_b : _GEN_1051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1053 = 9'h3f == r_count_3_io_out ? io_r_63_b : _GEN_1052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1054 = 9'h40 == r_count_3_io_out ? io_r_64_b : _GEN_1053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1055 = 9'h41 == r_count_3_io_out ? io_r_65_b : _GEN_1054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1056 = 9'h42 == r_count_3_io_out ? io_r_66_b : _GEN_1055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1057 = 9'h43 == r_count_3_io_out ? io_r_67_b : _GEN_1056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1058 = 9'h44 == r_count_3_io_out ? io_r_68_b : _GEN_1057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1059 = 9'h45 == r_count_3_io_out ? io_r_69_b : _GEN_1058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1060 = 9'h46 == r_count_3_io_out ? io_r_70_b : _GEN_1059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1061 = 9'h47 == r_count_3_io_out ? io_r_71_b : _GEN_1060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1062 = 9'h48 == r_count_3_io_out ? io_r_72_b : _GEN_1061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1063 = 9'h49 == r_count_3_io_out ? io_r_73_b : _GEN_1062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1064 = 9'h4a == r_count_3_io_out ? io_r_74_b : _GEN_1063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1065 = 9'h4b == r_count_3_io_out ? io_r_75_b : _GEN_1064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1066 = 9'h4c == r_count_3_io_out ? io_r_76_b : _GEN_1065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1067 = 9'h4d == r_count_3_io_out ? io_r_77_b : _GEN_1066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1068 = 9'h4e == r_count_3_io_out ? io_r_78_b : _GEN_1067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1069 = 9'h4f == r_count_3_io_out ? io_r_79_b : _GEN_1068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1070 = 9'h50 == r_count_3_io_out ? io_r_80_b : _GEN_1069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1071 = 9'h51 == r_count_3_io_out ? io_r_81_b : _GEN_1070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1072 = 9'h52 == r_count_3_io_out ? io_r_82_b : _GEN_1071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1073 = 9'h53 == r_count_3_io_out ? io_r_83_b : _GEN_1072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1074 = 9'h54 == r_count_3_io_out ? io_r_84_b : _GEN_1073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1075 = 9'h55 == r_count_3_io_out ? io_r_85_b : _GEN_1074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1076 = 9'h56 == r_count_3_io_out ? io_r_86_b : _GEN_1075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1077 = 9'h57 == r_count_3_io_out ? io_r_87_b : _GEN_1076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1078 = 9'h58 == r_count_3_io_out ? io_r_88_b : _GEN_1077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1079 = 9'h59 == r_count_3_io_out ? io_r_89_b : _GEN_1078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1080 = 9'h5a == r_count_3_io_out ? io_r_90_b : _GEN_1079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1081 = 9'h5b == r_count_3_io_out ? io_r_91_b : _GEN_1080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1082 = 9'h5c == r_count_3_io_out ? io_r_92_b : _GEN_1081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1083 = 9'h5d == r_count_3_io_out ? io_r_93_b : _GEN_1082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1084 = 9'h5e == r_count_3_io_out ? io_r_94_b : _GEN_1083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1085 = 9'h5f == r_count_3_io_out ? io_r_95_b : _GEN_1084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1086 = 9'h60 == r_count_3_io_out ? io_r_96_b : _GEN_1085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1087 = 9'h61 == r_count_3_io_out ? io_r_97_b : _GEN_1086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1088 = 9'h62 == r_count_3_io_out ? io_r_98_b : _GEN_1087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1089 = 9'h63 == r_count_3_io_out ? io_r_99_b : _GEN_1088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1090 = 9'h64 == r_count_3_io_out ? io_r_100_b : _GEN_1089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1091 = 9'h65 == r_count_3_io_out ? io_r_101_b : _GEN_1090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1092 = 9'h66 == r_count_3_io_out ? io_r_102_b : _GEN_1091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1093 = 9'h67 == r_count_3_io_out ? io_r_103_b : _GEN_1092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1094 = 9'h68 == r_count_3_io_out ? io_r_104_b : _GEN_1093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1095 = 9'h69 == r_count_3_io_out ? io_r_105_b : _GEN_1094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1096 = 9'h6a == r_count_3_io_out ? io_r_106_b : _GEN_1095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1097 = 9'h6b == r_count_3_io_out ? io_r_107_b : _GEN_1096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1098 = 9'h6c == r_count_3_io_out ? io_r_108_b : _GEN_1097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1099 = 9'h6d == r_count_3_io_out ? io_r_109_b : _GEN_1098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1100 = 9'h6e == r_count_3_io_out ? io_r_110_b : _GEN_1099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1101 = 9'h6f == r_count_3_io_out ? io_r_111_b : _GEN_1100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1102 = 9'h70 == r_count_3_io_out ? io_r_112_b : _GEN_1101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1103 = 9'h71 == r_count_3_io_out ? io_r_113_b : _GEN_1102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1104 = 9'h72 == r_count_3_io_out ? io_r_114_b : _GEN_1103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1105 = 9'h73 == r_count_3_io_out ? io_r_115_b : _GEN_1104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1106 = 9'h74 == r_count_3_io_out ? io_r_116_b : _GEN_1105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1107 = 9'h75 == r_count_3_io_out ? io_r_117_b : _GEN_1106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1108 = 9'h76 == r_count_3_io_out ? io_r_118_b : _GEN_1107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1109 = 9'h77 == r_count_3_io_out ? io_r_119_b : _GEN_1108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1110 = 9'h78 == r_count_3_io_out ? io_r_120_b : _GEN_1109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1111 = 9'h79 == r_count_3_io_out ? io_r_121_b : _GEN_1110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1112 = 9'h7a == r_count_3_io_out ? io_r_122_b : _GEN_1111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1113 = 9'h7b == r_count_3_io_out ? io_r_123_b : _GEN_1112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1114 = 9'h7c == r_count_3_io_out ? io_r_124_b : _GEN_1113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1115 = 9'h7d == r_count_3_io_out ? io_r_125_b : _GEN_1114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1116 = 9'h7e == r_count_3_io_out ? io_r_126_b : _GEN_1115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1117 = 9'h7f == r_count_3_io_out ? io_r_127_b : _GEN_1116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1118 = 9'h80 == r_count_3_io_out ? io_r_128_b : _GEN_1117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1119 = 9'h81 == r_count_3_io_out ? io_r_129_b : _GEN_1118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1120 = 9'h82 == r_count_3_io_out ? io_r_130_b : _GEN_1119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1121 = 9'h83 == r_count_3_io_out ? io_r_131_b : _GEN_1120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1122 = 9'h84 == r_count_3_io_out ? io_r_132_b : _GEN_1121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1123 = 9'h85 == r_count_3_io_out ? io_r_133_b : _GEN_1122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1124 = 9'h86 == r_count_3_io_out ? io_r_134_b : _GEN_1123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1125 = 9'h87 == r_count_3_io_out ? io_r_135_b : _GEN_1124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1126 = 9'h88 == r_count_3_io_out ? io_r_136_b : _GEN_1125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1127 = 9'h89 == r_count_3_io_out ? io_r_137_b : _GEN_1126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1128 = 9'h8a == r_count_3_io_out ? io_r_138_b : _GEN_1127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1129 = 9'h8b == r_count_3_io_out ? io_r_139_b : _GEN_1128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1130 = 9'h8c == r_count_3_io_out ? io_r_140_b : _GEN_1129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1131 = 9'h8d == r_count_3_io_out ? io_r_141_b : _GEN_1130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1132 = 9'h8e == r_count_3_io_out ? io_r_142_b : _GEN_1131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1133 = 9'h8f == r_count_3_io_out ? io_r_143_b : _GEN_1132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1134 = 9'h90 == r_count_3_io_out ? io_r_144_b : _GEN_1133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1135 = 9'h91 == r_count_3_io_out ? io_r_145_b : _GEN_1134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1136 = 9'h92 == r_count_3_io_out ? io_r_146_b : _GEN_1135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1137 = 9'h93 == r_count_3_io_out ? io_r_147_b : _GEN_1136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1138 = 9'h94 == r_count_3_io_out ? io_r_148_b : _GEN_1137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1139 = 9'h95 == r_count_3_io_out ? io_r_149_b : _GEN_1138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1140 = 9'h96 == r_count_3_io_out ? io_r_150_b : _GEN_1139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1141 = 9'h97 == r_count_3_io_out ? io_r_151_b : _GEN_1140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1142 = 9'h98 == r_count_3_io_out ? io_r_152_b : _GEN_1141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1143 = 9'h99 == r_count_3_io_out ? io_r_153_b : _GEN_1142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1144 = 9'h9a == r_count_3_io_out ? io_r_154_b : _GEN_1143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1145 = 9'h9b == r_count_3_io_out ? io_r_155_b : _GEN_1144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1146 = 9'h9c == r_count_3_io_out ? io_r_156_b : _GEN_1145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1147 = 9'h9d == r_count_3_io_out ? io_r_157_b : _GEN_1146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1148 = 9'h9e == r_count_3_io_out ? io_r_158_b : _GEN_1147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1149 = 9'h9f == r_count_3_io_out ? io_r_159_b : _GEN_1148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1150 = 9'ha0 == r_count_3_io_out ? io_r_160_b : _GEN_1149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1151 = 9'ha1 == r_count_3_io_out ? io_r_161_b : _GEN_1150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1152 = 9'ha2 == r_count_3_io_out ? io_r_162_b : _GEN_1151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1153 = 9'ha3 == r_count_3_io_out ? io_r_163_b : _GEN_1152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1154 = 9'ha4 == r_count_3_io_out ? io_r_164_b : _GEN_1153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1155 = 9'ha5 == r_count_3_io_out ? io_r_165_b : _GEN_1154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1156 = 9'ha6 == r_count_3_io_out ? io_r_166_b : _GEN_1155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1157 = 9'ha7 == r_count_3_io_out ? io_r_167_b : _GEN_1156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1158 = 9'ha8 == r_count_3_io_out ? io_r_168_b : _GEN_1157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1159 = 9'ha9 == r_count_3_io_out ? io_r_169_b : _GEN_1158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1160 = 9'haa == r_count_3_io_out ? io_r_170_b : _GEN_1159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1161 = 9'hab == r_count_3_io_out ? io_r_171_b : _GEN_1160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1162 = 9'hac == r_count_3_io_out ? io_r_172_b : _GEN_1161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1163 = 9'had == r_count_3_io_out ? io_r_173_b : _GEN_1162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1164 = 9'hae == r_count_3_io_out ? io_r_174_b : _GEN_1163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1165 = 9'haf == r_count_3_io_out ? io_r_175_b : _GEN_1164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1166 = 9'hb0 == r_count_3_io_out ? io_r_176_b : _GEN_1165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1167 = 9'hb1 == r_count_3_io_out ? io_r_177_b : _GEN_1166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1168 = 9'hb2 == r_count_3_io_out ? io_r_178_b : _GEN_1167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1169 = 9'hb3 == r_count_3_io_out ? io_r_179_b : _GEN_1168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1170 = 9'hb4 == r_count_3_io_out ? io_r_180_b : _GEN_1169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1171 = 9'hb5 == r_count_3_io_out ? io_r_181_b : _GEN_1170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1172 = 9'hb6 == r_count_3_io_out ? io_r_182_b : _GEN_1171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1173 = 9'hb7 == r_count_3_io_out ? io_r_183_b : _GEN_1172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1174 = 9'hb8 == r_count_3_io_out ? io_r_184_b : _GEN_1173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1175 = 9'hb9 == r_count_3_io_out ? io_r_185_b : _GEN_1174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1176 = 9'hba == r_count_3_io_out ? io_r_186_b : _GEN_1175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1177 = 9'hbb == r_count_3_io_out ? io_r_187_b : _GEN_1176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1178 = 9'hbc == r_count_3_io_out ? io_r_188_b : _GEN_1177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1179 = 9'hbd == r_count_3_io_out ? io_r_189_b : _GEN_1178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1180 = 9'hbe == r_count_3_io_out ? io_r_190_b : _GEN_1179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1181 = 9'hbf == r_count_3_io_out ? io_r_191_b : _GEN_1180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1182 = 9'hc0 == r_count_3_io_out ? io_r_192_b : _GEN_1181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1183 = 9'hc1 == r_count_3_io_out ? io_r_193_b : _GEN_1182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1184 = 9'hc2 == r_count_3_io_out ? io_r_194_b : _GEN_1183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1185 = 9'hc3 == r_count_3_io_out ? io_r_195_b : _GEN_1184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1186 = 9'hc4 == r_count_3_io_out ? io_r_196_b : _GEN_1185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1187 = 9'hc5 == r_count_3_io_out ? io_r_197_b : _GEN_1186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1188 = 9'hc6 == r_count_3_io_out ? io_r_198_b : _GEN_1187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1189 = 9'hc7 == r_count_3_io_out ? io_r_199_b : _GEN_1188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1190 = 9'hc8 == r_count_3_io_out ? io_r_200_b : _GEN_1189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1191 = 9'hc9 == r_count_3_io_out ? io_r_201_b : _GEN_1190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1192 = 9'hca == r_count_3_io_out ? io_r_202_b : _GEN_1191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1193 = 9'hcb == r_count_3_io_out ? io_r_203_b : _GEN_1192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1194 = 9'hcc == r_count_3_io_out ? io_r_204_b : _GEN_1193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1195 = 9'hcd == r_count_3_io_out ? io_r_205_b : _GEN_1194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1196 = 9'hce == r_count_3_io_out ? io_r_206_b : _GEN_1195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1197 = 9'hcf == r_count_3_io_out ? io_r_207_b : _GEN_1196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1198 = 9'hd0 == r_count_3_io_out ? io_r_208_b : _GEN_1197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1199 = 9'hd1 == r_count_3_io_out ? io_r_209_b : _GEN_1198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1200 = 9'hd2 == r_count_3_io_out ? io_r_210_b : _GEN_1199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1201 = 9'hd3 == r_count_3_io_out ? io_r_211_b : _GEN_1200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1202 = 9'hd4 == r_count_3_io_out ? io_r_212_b : _GEN_1201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1203 = 9'hd5 == r_count_3_io_out ? io_r_213_b : _GEN_1202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1204 = 9'hd6 == r_count_3_io_out ? io_r_214_b : _GEN_1203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1205 = 9'hd7 == r_count_3_io_out ? io_r_215_b : _GEN_1204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1206 = 9'hd8 == r_count_3_io_out ? io_r_216_b : _GEN_1205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1207 = 9'hd9 == r_count_3_io_out ? io_r_217_b : _GEN_1206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1208 = 9'hda == r_count_3_io_out ? io_r_218_b : _GEN_1207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1209 = 9'hdb == r_count_3_io_out ? io_r_219_b : _GEN_1208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1210 = 9'hdc == r_count_3_io_out ? io_r_220_b : _GEN_1209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1211 = 9'hdd == r_count_3_io_out ? io_r_221_b : _GEN_1210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1212 = 9'hde == r_count_3_io_out ? io_r_222_b : _GEN_1211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1213 = 9'hdf == r_count_3_io_out ? io_r_223_b : _GEN_1212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1214 = 9'he0 == r_count_3_io_out ? io_r_224_b : _GEN_1213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1215 = 9'he1 == r_count_3_io_out ? io_r_225_b : _GEN_1214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1216 = 9'he2 == r_count_3_io_out ? io_r_226_b : _GEN_1215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1217 = 9'he3 == r_count_3_io_out ? io_r_227_b : _GEN_1216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1218 = 9'he4 == r_count_3_io_out ? io_r_228_b : _GEN_1217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1219 = 9'he5 == r_count_3_io_out ? io_r_229_b : _GEN_1218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1220 = 9'he6 == r_count_3_io_out ? io_r_230_b : _GEN_1219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1221 = 9'he7 == r_count_3_io_out ? io_r_231_b : _GEN_1220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1222 = 9'he8 == r_count_3_io_out ? io_r_232_b : _GEN_1221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1223 = 9'he9 == r_count_3_io_out ? io_r_233_b : _GEN_1222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1224 = 9'hea == r_count_3_io_out ? io_r_234_b : _GEN_1223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1225 = 9'heb == r_count_3_io_out ? io_r_235_b : _GEN_1224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1226 = 9'hec == r_count_3_io_out ? io_r_236_b : _GEN_1225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1227 = 9'hed == r_count_3_io_out ? io_r_237_b : _GEN_1226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1228 = 9'hee == r_count_3_io_out ? io_r_238_b : _GEN_1227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1229 = 9'hef == r_count_3_io_out ? io_r_239_b : _GEN_1228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1230 = 9'hf0 == r_count_3_io_out ? io_r_240_b : _GEN_1229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1231 = 9'hf1 == r_count_3_io_out ? io_r_241_b : _GEN_1230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1232 = 9'hf2 == r_count_3_io_out ? io_r_242_b : _GEN_1231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1233 = 9'hf3 == r_count_3_io_out ? io_r_243_b : _GEN_1232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1234 = 9'hf4 == r_count_3_io_out ? io_r_244_b : _GEN_1233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1235 = 9'hf5 == r_count_3_io_out ? io_r_245_b : _GEN_1234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1236 = 9'hf6 == r_count_3_io_out ? io_r_246_b : _GEN_1235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1237 = 9'hf7 == r_count_3_io_out ? io_r_247_b : _GEN_1236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1238 = 9'hf8 == r_count_3_io_out ? io_r_248_b : _GEN_1237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1239 = 9'hf9 == r_count_3_io_out ? io_r_249_b : _GEN_1238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1240 = 9'hfa == r_count_3_io_out ? io_r_250_b : _GEN_1239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1241 = 9'hfb == r_count_3_io_out ? io_r_251_b : _GEN_1240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1242 = 9'hfc == r_count_3_io_out ? io_r_252_b : _GEN_1241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1243 = 9'hfd == r_count_3_io_out ? io_r_253_b : _GEN_1242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1244 = 9'hfe == r_count_3_io_out ? io_r_254_b : _GEN_1243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1245 = 9'hff == r_count_3_io_out ? io_r_255_b : _GEN_1244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1246 = 9'h100 == r_count_3_io_out ? io_r_256_b : _GEN_1245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1247 = 9'h101 == r_count_3_io_out ? io_r_257_b : _GEN_1246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1248 = 9'h102 == r_count_3_io_out ? io_r_258_b : _GEN_1247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1249 = 9'h103 == r_count_3_io_out ? io_r_259_b : _GEN_1248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1250 = 9'h104 == r_count_3_io_out ? io_r_260_b : _GEN_1249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1251 = 9'h105 == r_count_3_io_out ? io_r_261_b : _GEN_1250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1252 = 9'h106 == r_count_3_io_out ? io_r_262_b : _GEN_1251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1253 = 9'h107 == r_count_3_io_out ? io_r_263_b : _GEN_1252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1254 = 9'h108 == r_count_3_io_out ? io_r_264_b : _GEN_1253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1255 = 9'h109 == r_count_3_io_out ? io_r_265_b : _GEN_1254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1256 = 9'h10a == r_count_3_io_out ? io_r_266_b : _GEN_1255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1257 = 9'h10b == r_count_3_io_out ? io_r_267_b : _GEN_1256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1258 = 9'h10c == r_count_3_io_out ? io_r_268_b : _GEN_1257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1259 = 9'h10d == r_count_3_io_out ? io_r_269_b : _GEN_1258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1260 = 9'h10e == r_count_3_io_out ? io_r_270_b : _GEN_1259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1261 = 9'h10f == r_count_3_io_out ? io_r_271_b : _GEN_1260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1262 = 9'h110 == r_count_3_io_out ? io_r_272_b : _GEN_1261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1263 = 9'h111 == r_count_3_io_out ? io_r_273_b : _GEN_1262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1264 = 9'h112 == r_count_3_io_out ? io_r_274_b : _GEN_1263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1265 = 9'h113 == r_count_3_io_out ? io_r_275_b : _GEN_1264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1266 = 9'h114 == r_count_3_io_out ? io_r_276_b : _GEN_1265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1267 = 9'h115 == r_count_3_io_out ? io_r_277_b : _GEN_1266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1268 = 9'h116 == r_count_3_io_out ? io_r_278_b : _GEN_1267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1269 = 9'h117 == r_count_3_io_out ? io_r_279_b : _GEN_1268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1270 = 9'h118 == r_count_3_io_out ? io_r_280_b : _GEN_1269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1271 = 9'h119 == r_count_3_io_out ? io_r_281_b : _GEN_1270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1272 = 9'h11a == r_count_3_io_out ? io_r_282_b : _GEN_1271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1273 = 9'h11b == r_count_3_io_out ? io_r_283_b : _GEN_1272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1274 = 9'h11c == r_count_3_io_out ? io_r_284_b : _GEN_1273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1275 = 9'h11d == r_count_3_io_out ? io_r_285_b : _GEN_1274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1276 = 9'h11e == r_count_3_io_out ? io_r_286_b : _GEN_1275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1277 = 9'h11f == r_count_3_io_out ? io_r_287_b : _GEN_1276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1278 = 9'h120 == r_count_3_io_out ? io_r_288_b : _GEN_1277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1279 = 9'h121 == r_count_3_io_out ? io_r_289_b : _GEN_1278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1280 = 9'h122 == r_count_3_io_out ? io_r_290_b : _GEN_1279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1281 = 9'h123 == r_count_3_io_out ? io_r_291_b : _GEN_1280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1282 = 9'h124 == r_count_3_io_out ? io_r_292_b : _GEN_1281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1283 = 9'h125 == r_count_3_io_out ? io_r_293_b : _GEN_1282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1284 = 9'h126 == r_count_3_io_out ? io_r_294_b : _GEN_1283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1285 = 9'h127 == r_count_3_io_out ? io_r_295_b : _GEN_1284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1286 = 9'h128 == r_count_3_io_out ? io_r_296_b : _GEN_1285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1287 = 9'h129 == r_count_3_io_out ? io_r_297_b : _GEN_1286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1288 = 9'h12a == r_count_3_io_out ? io_r_298_b : _GEN_1287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1291 = 9'h1 == r_count_4_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1292 = 9'h2 == r_count_4_io_out ? io_r_2_b : _GEN_1291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1293 = 9'h3 == r_count_4_io_out ? io_r_3_b : _GEN_1292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1294 = 9'h4 == r_count_4_io_out ? io_r_4_b : _GEN_1293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1295 = 9'h5 == r_count_4_io_out ? io_r_5_b : _GEN_1294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1296 = 9'h6 == r_count_4_io_out ? io_r_6_b : _GEN_1295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1297 = 9'h7 == r_count_4_io_out ? io_r_7_b : _GEN_1296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1298 = 9'h8 == r_count_4_io_out ? io_r_8_b : _GEN_1297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1299 = 9'h9 == r_count_4_io_out ? io_r_9_b : _GEN_1298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1300 = 9'ha == r_count_4_io_out ? io_r_10_b : _GEN_1299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1301 = 9'hb == r_count_4_io_out ? io_r_11_b : _GEN_1300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1302 = 9'hc == r_count_4_io_out ? io_r_12_b : _GEN_1301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1303 = 9'hd == r_count_4_io_out ? io_r_13_b : _GEN_1302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1304 = 9'he == r_count_4_io_out ? io_r_14_b : _GEN_1303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1305 = 9'hf == r_count_4_io_out ? io_r_15_b : _GEN_1304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1306 = 9'h10 == r_count_4_io_out ? io_r_16_b : _GEN_1305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1307 = 9'h11 == r_count_4_io_out ? io_r_17_b : _GEN_1306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1308 = 9'h12 == r_count_4_io_out ? io_r_18_b : _GEN_1307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1309 = 9'h13 == r_count_4_io_out ? io_r_19_b : _GEN_1308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1310 = 9'h14 == r_count_4_io_out ? io_r_20_b : _GEN_1309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1311 = 9'h15 == r_count_4_io_out ? io_r_21_b : _GEN_1310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1312 = 9'h16 == r_count_4_io_out ? io_r_22_b : _GEN_1311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1313 = 9'h17 == r_count_4_io_out ? io_r_23_b : _GEN_1312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1314 = 9'h18 == r_count_4_io_out ? io_r_24_b : _GEN_1313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1315 = 9'h19 == r_count_4_io_out ? io_r_25_b : _GEN_1314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1316 = 9'h1a == r_count_4_io_out ? io_r_26_b : _GEN_1315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1317 = 9'h1b == r_count_4_io_out ? io_r_27_b : _GEN_1316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1318 = 9'h1c == r_count_4_io_out ? io_r_28_b : _GEN_1317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1319 = 9'h1d == r_count_4_io_out ? io_r_29_b : _GEN_1318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1320 = 9'h1e == r_count_4_io_out ? io_r_30_b : _GEN_1319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1321 = 9'h1f == r_count_4_io_out ? io_r_31_b : _GEN_1320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1322 = 9'h20 == r_count_4_io_out ? io_r_32_b : _GEN_1321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1323 = 9'h21 == r_count_4_io_out ? io_r_33_b : _GEN_1322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1324 = 9'h22 == r_count_4_io_out ? io_r_34_b : _GEN_1323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1325 = 9'h23 == r_count_4_io_out ? io_r_35_b : _GEN_1324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1326 = 9'h24 == r_count_4_io_out ? io_r_36_b : _GEN_1325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1327 = 9'h25 == r_count_4_io_out ? io_r_37_b : _GEN_1326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1328 = 9'h26 == r_count_4_io_out ? io_r_38_b : _GEN_1327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1329 = 9'h27 == r_count_4_io_out ? io_r_39_b : _GEN_1328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1330 = 9'h28 == r_count_4_io_out ? io_r_40_b : _GEN_1329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1331 = 9'h29 == r_count_4_io_out ? io_r_41_b : _GEN_1330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1332 = 9'h2a == r_count_4_io_out ? io_r_42_b : _GEN_1331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1333 = 9'h2b == r_count_4_io_out ? io_r_43_b : _GEN_1332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1334 = 9'h2c == r_count_4_io_out ? io_r_44_b : _GEN_1333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1335 = 9'h2d == r_count_4_io_out ? io_r_45_b : _GEN_1334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1336 = 9'h2e == r_count_4_io_out ? io_r_46_b : _GEN_1335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1337 = 9'h2f == r_count_4_io_out ? io_r_47_b : _GEN_1336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1338 = 9'h30 == r_count_4_io_out ? io_r_48_b : _GEN_1337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1339 = 9'h31 == r_count_4_io_out ? io_r_49_b : _GEN_1338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1340 = 9'h32 == r_count_4_io_out ? io_r_50_b : _GEN_1339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1341 = 9'h33 == r_count_4_io_out ? io_r_51_b : _GEN_1340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1342 = 9'h34 == r_count_4_io_out ? io_r_52_b : _GEN_1341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1343 = 9'h35 == r_count_4_io_out ? io_r_53_b : _GEN_1342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1344 = 9'h36 == r_count_4_io_out ? io_r_54_b : _GEN_1343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1345 = 9'h37 == r_count_4_io_out ? io_r_55_b : _GEN_1344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1346 = 9'h38 == r_count_4_io_out ? io_r_56_b : _GEN_1345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1347 = 9'h39 == r_count_4_io_out ? io_r_57_b : _GEN_1346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1348 = 9'h3a == r_count_4_io_out ? io_r_58_b : _GEN_1347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1349 = 9'h3b == r_count_4_io_out ? io_r_59_b : _GEN_1348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1350 = 9'h3c == r_count_4_io_out ? io_r_60_b : _GEN_1349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1351 = 9'h3d == r_count_4_io_out ? io_r_61_b : _GEN_1350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1352 = 9'h3e == r_count_4_io_out ? io_r_62_b : _GEN_1351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1353 = 9'h3f == r_count_4_io_out ? io_r_63_b : _GEN_1352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1354 = 9'h40 == r_count_4_io_out ? io_r_64_b : _GEN_1353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1355 = 9'h41 == r_count_4_io_out ? io_r_65_b : _GEN_1354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1356 = 9'h42 == r_count_4_io_out ? io_r_66_b : _GEN_1355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1357 = 9'h43 == r_count_4_io_out ? io_r_67_b : _GEN_1356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1358 = 9'h44 == r_count_4_io_out ? io_r_68_b : _GEN_1357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1359 = 9'h45 == r_count_4_io_out ? io_r_69_b : _GEN_1358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1360 = 9'h46 == r_count_4_io_out ? io_r_70_b : _GEN_1359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1361 = 9'h47 == r_count_4_io_out ? io_r_71_b : _GEN_1360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1362 = 9'h48 == r_count_4_io_out ? io_r_72_b : _GEN_1361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1363 = 9'h49 == r_count_4_io_out ? io_r_73_b : _GEN_1362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1364 = 9'h4a == r_count_4_io_out ? io_r_74_b : _GEN_1363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1365 = 9'h4b == r_count_4_io_out ? io_r_75_b : _GEN_1364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1366 = 9'h4c == r_count_4_io_out ? io_r_76_b : _GEN_1365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1367 = 9'h4d == r_count_4_io_out ? io_r_77_b : _GEN_1366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1368 = 9'h4e == r_count_4_io_out ? io_r_78_b : _GEN_1367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1369 = 9'h4f == r_count_4_io_out ? io_r_79_b : _GEN_1368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1370 = 9'h50 == r_count_4_io_out ? io_r_80_b : _GEN_1369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1371 = 9'h51 == r_count_4_io_out ? io_r_81_b : _GEN_1370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1372 = 9'h52 == r_count_4_io_out ? io_r_82_b : _GEN_1371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1373 = 9'h53 == r_count_4_io_out ? io_r_83_b : _GEN_1372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1374 = 9'h54 == r_count_4_io_out ? io_r_84_b : _GEN_1373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1375 = 9'h55 == r_count_4_io_out ? io_r_85_b : _GEN_1374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1376 = 9'h56 == r_count_4_io_out ? io_r_86_b : _GEN_1375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1377 = 9'h57 == r_count_4_io_out ? io_r_87_b : _GEN_1376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1378 = 9'h58 == r_count_4_io_out ? io_r_88_b : _GEN_1377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1379 = 9'h59 == r_count_4_io_out ? io_r_89_b : _GEN_1378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1380 = 9'h5a == r_count_4_io_out ? io_r_90_b : _GEN_1379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1381 = 9'h5b == r_count_4_io_out ? io_r_91_b : _GEN_1380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1382 = 9'h5c == r_count_4_io_out ? io_r_92_b : _GEN_1381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1383 = 9'h5d == r_count_4_io_out ? io_r_93_b : _GEN_1382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1384 = 9'h5e == r_count_4_io_out ? io_r_94_b : _GEN_1383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1385 = 9'h5f == r_count_4_io_out ? io_r_95_b : _GEN_1384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1386 = 9'h60 == r_count_4_io_out ? io_r_96_b : _GEN_1385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1387 = 9'h61 == r_count_4_io_out ? io_r_97_b : _GEN_1386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1388 = 9'h62 == r_count_4_io_out ? io_r_98_b : _GEN_1387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1389 = 9'h63 == r_count_4_io_out ? io_r_99_b : _GEN_1388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1390 = 9'h64 == r_count_4_io_out ? io_r_100_b : _GEN_1389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1391 = 9'h65 == r_count_4_io_out ? io_r_101_b : _GEN_1390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1392 = 9'h66 == r_count_4_io_out ? io_r_102_b : _GEN_1391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1393 = 9'h67 == r_count_4_io_out ? io_r_103_b : _GEN_1392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1394 = 9'h68 == r_count_4_io_out ? io_r_104_b : _GEN_1393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1395 = 9'h69 == r_count_4_io_out ? io_r_105_b : _GEN_1394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1396 = 9'h6a == r_count_4_io_out ? io_r_106_b : _GEN_1395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1397 = 9'h6b == r_count_4_io_out ? io_r_107_b : _GEN_1396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1398 = 9'h6c == r_count_4_io_out ? io_r_108_b : _GEN_1397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1399 = 9'h6d == r_count_4_io_out ? io_r_109_b : _GEN_1398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1400 = 9'h6e == r_count_4_io_out ? io_r_110_b : _GEN_1399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1401 = 9'h6f == r_count_4_io_out ? io_r_111_b : _GEN_1400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1402 = 9'h70 == r_count_4_io_out ? io_r_112_b : _GEN_1401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1403 = 9'h71 == r_count_4_io_out ? io_r_113_b : _GEN_1402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1404 = 9'h72 == r_count_4_io_out ? io_r_114_b : _GEN_1403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1405 = 9'h73 == r_count_4_io_out ? io_r_115_b : _GEN_1404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1406 = 9'h74 == r_count_4_io_out ? io_r_116_b : _GEN_1405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1407 = 9'h75 == r_count_4_io_out ? io_r_117_b : _GEN_1406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1408 = 9'h76 == r_count_4_io_out ? io_r_118_b : _GEN_1407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1409 = 9'h77 == r_count_4_io_out ? io_r_119_b : _GEN_1408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1410 = 9'h78 == r_count_4_io_out ? io_r_120_b : _GEN_1409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1411 = 9'h79 == r_count_4_io_out ? io_r_121_b : _GEN_1410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1412 = 9'h7a == r_count_4_io_out ? io_r_122_b : _GEN_1411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1413 = 9'h7b == r_count_4_io_out ? io_r_123_b : _GEN_1412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1414 = 9'h7c == r_count_4_io_out ? io_r_124_b : _GEN_1413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1415 = 9'h7d == r_count_4_io_out ? io_r_125_b : _GEN_1414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1416 = 9'h7e == r_count_4_io_out ? io_r_126_b : _GEN_1415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1417 = 9'h7f == r_count_4_io_out ? io_r_127_b : _GEN_1416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1418 = 9'h80 == r_count_4_io_out ? io_r_128_b : _GEN_1417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1419 = 9'h81 == r_count_4_io_out ? io_r_129_b : _GEN_1418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1420 = 9'h82 == r_count_4_io_out ? io_r_130_b : _GEN_1419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1421 = 9'h83 == r_count_4_io_out ? io_r_131_b : _GEN_1420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1422 = 9'h84 == r_count_4_io_out ? io_r_132_b : _GEN_1421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1423 = 9'h85 == r_count_4_io_out ? io_r_133_b : _GEN_1422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1424 = 9'h86 == r_count_4_io_out ? io_r_134_b : _GEN_1423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1425 = 9'h87 == r_count_4_io_out ? io_r_135_b : _GEN_1424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1426 = 9'h88 == r_count_4_io_out ? io_r_136_b : _GEN_1425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1427 = 9'h89 == r_count_4_io_out ? io_r_137_b : _GEN_1426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1428 = 9'h8a == r_count_4_io_out ? io_r_138_b : _GEN_1427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1429 = 9'h8b == r_count_4_io_out ? io_r_139_b : _GEN_1428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1430 = 9'h8c == r_count_4_io_out ? io_r_140_b : _GEN_1429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1431 = 9'h8d == r_count_4_io_out ? io_r_141_b : _GEN_1430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1432 = 9'h8e == r_count_4_io_out ? io_r_142_b : _GEN_1431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1433 = 9'h8f == r_count_4_io_out ? io_r_143_b : _GEN_1432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1434 = 9'h90 == r_count_4_io_out ? io_r_144_b : _GEN_1433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1435 = 9'h91 == r_count_4_io_out ? io_r_145_b : _GEN_1434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1436 = 9'h92 == r_count_4_io_out ? io_r_146_b : _GEN_1435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1437 = 9'h93 == r_count_4_io_out ? io_r_147_b : _GEN_1436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1438 = 9'h94 == r_count_4_io_out ? io_r_148_b : _GEN_1437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1439 = 9'h95 == r_count_4_io_out ? io_r_149_b : _GEN_1438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1440 = 9'h96 == r_count_4_io_out ? io_r_150_b : _GEN_1439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1441 = 9'h97 == r_count_4_io_out ? io_r_151_b : _GEN_1440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1442 = 9'h98 == r_count_4_io_out ? io_r_152_b : _GEN_1441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1443 = 9'h99 == r_count_4_io_out ? io_r_153_b : _GEN_1442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1444 = 9'h9a == r_count_4_io_out ? io_r_154_b : _GEN_1443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1445 = 9'h9b == r_count_4_io_out ? io_r_155_b : _GEN_1444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1446 = 9'h9c == r_count_4_io_out ? io_r_156_b : _GEN_1445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1447 = 9'h9d == r_count_4_io_out ? io_r_157_b : _GEN_1446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1448 = 9'h9e == r_count_4_io_out ? io_r_158_b : _GEN_1447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1449 = 9'h9f == r_count_4_io_out ? io_r_159_b : _GEN_1448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1450 = 9'ha0 == r_count_4_io_out ? io_r_160_b : _GEN_1449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1451 = 9'ha1 == r_count_4_io_out ? io_r_161_b : _GEN_1450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1452 = 9'ha2 == r_count_4_io_out ? io_r_162_b : _GEN_1451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1453 = 9'ha3 == r_count_4_io_out ? io_r_163_b : _GEN_1452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1454 = 9'ha4 == r_count_4_io_out ? io_r_164_b : _GEN_1453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1455 = 9'ha5 == r_count_4_io_out ? io_r_165_b : _GEN_1454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1456 = 9'ha6 == r_count_4_io_out ? io_r_166_b : _GEN_1455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1457 = 9'ha7 == r_count_4_io_out ? io_r_167_b : _GEN_1456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1458 = 9'ha8 == r_count_4_io_out ? io_r_168_b : _GEN_1457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1459 = 9'ha9 == r_count_4_io_out ? io_r_169_b : _GEN_1458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1460 = 9'haa == r_count_4_io_out ? io_r_170_b : _GEN_1459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1461 = 9'hab == r_count_4_io_out ? io_r_171_b : _GEN_1460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1462 = 9'hac == r_count_4_io_out ? io_r_172_b : _GEN_1461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1463 = 9'had == r_count_4_io_out ? io_r_173_b : _GEN_1462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1464 = 9'hae == r_count_4_io_out ? io_r_174_b : _GEN_1463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1465 = 9'haf == r_count_4_io_out ? io_r_175_b : _GEN_1464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1466 = 9'hb0 == r_count_4_io_out ? io_r_176_b : _GEN_1465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1467 = 9'hb1 == r_count_4_io_out ? io_r_177_b : _GEN_1466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1468 = 9'hb2 == r_count_4_io_out ? io_r_178_b : _GEN_1467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1469 = 9'hb3 == r_count_4_io_out ? io_r_179_b : _GEN_1468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1470 = 9'hb4 == r_count_4_io_out ? io_r_180_b : _GEN_1469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1471 = 9'hb5 == r_count_4_io_out ? io_r_181_b : _GEN_1470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1472 = 9'hb6 == r_count_4_io_out ? io_r_182_b : _GEN_1471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1473 = 9'hb7 == r_count_4_io_out ? io_r_183_b : _GEN_1472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1474 = 9'hb8 == r_count_4_io_out ? io_r_184_b : _GEN_1473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1475 = 9'hb9 == r_count_4_io_out ? io_r_185_b : _GEN_1474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1476 = 9'hba == r_count_4_io_out ? io_r_186_b : _GEN_1475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1477 = 9'hbb == r_count_4_io_out ? io_r_187_b : _GEN_1476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1478 = 9'hbc == r_count_4_io_out ? io_r_188_b : _GEN_1477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1479 = 9'hbd == r_count_4_io_out ? io_r_189_b : _GEN_1478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1480 = 9'hbe == r_count_4_io_out ? io_r_190_b : _GEN_1479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1481 = 9'hbf == r_count_4_io_out ? io_r_191_b : _GEN_1480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1482 = 9'hc0 == r_count_4_io_out ? io_r_192_b : _GEN_1481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1483 = 9'hc1 == r_count_4_io_out ? io_r_193_b : _GEN_1482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1484 = 9'hc2 == r_count_4_io_out ? io_r_194_b : _GEN_1483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1485 = 9'hc3 == r_count_4_io_out ? io_r_195_b : _GEN_1484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1486 = 9'hc4 == r_count_4_io_out ? io_r_196_b : _GEN_1485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1487 = 9'hc5 == r_count_4_io_out ? io_r_197_b : _GEN_1486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1488 = 9'hc6 == r_count_4_io_out ? io_r_198_b : _GEN_1487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1489 = 9'hc7 == r_count_4_io_out ? io_r_199_b : _GEN_1488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1490 = 9'hc8 == r_count_4_io_out ? io_r_200_b : _GEN_1489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1491 = 9'hc9 == r_count_4_io_out ? io_r_201_b : _GEN_1490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1492 = 9'hca == r_count_4_io_out ? io_r_202_b : _GEN_1491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1493 = 9'hcb == r_count_4_io_out ? io_r_203_b : _GEN_1492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1494 = 9'hcc == r_count_4_io_out ? io_r_204_b : _GEN_1493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1495 = 9'hcd == r_count_4_io_out ? io_r_205_b : _GEN_1494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1496 = 9'hce == r_count_4_io_out ? io_r_206_b : _GEN_1495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1497 = 9'hcf == r_count_4_io_out ? io_r_207_b : _GEN_1496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1498 = 9'hd0 == r_count_4_io_out ? io_r_208_b : _GEN_1497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1499 = 9'hd1 == r_count_4_io_out ? io_r_209_b : _GEN_1498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1500 = 9'hd2 == r_count_4_io_out ? io_r_210_b : _GEN_1499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1501 = 9'hd3 == r_count_4_io_out ? io_r_211_b : _GEN_1500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1502 = 9'hd4 == r_count_4_io_out ? io_r_212_b : _GEN_1501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1503 = 9'hd5 == r_count_4_io_out ? io_r_213_b : _GEN_1502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1504 = 9'hd6 == r_count_4_io_out ? io_r_214_b : _GEN_1503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1505 = 9'hd7 == r_count_4_io_out ? io_r_215_b : _GEN_1504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1506 = 9'hd8 == r_count_4_io_out ? io_r_216_b : _GEN_1505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1507 = 9'hd9 == r_count_4_io_out ? io_r_217_b : _GEN_1506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1508 = 9'hda == r_count_4_io_out ? io_r_218_b : _GEN_1507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1509 = 9'hdb == r_count_4_io_out ? io_r_219_b : _GEN_1508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1510 = 9'hdc == r_count_4_io_out ? io_r_220_b : _GEN_1509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1511 = 9'hdd == r_count_4_io_out ? io_r_221_b : _GEN_1510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1512 = 9'hde == r_count_4_io_out ? io_r_222_b : _GEN_1511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1513 = 9'hdf == r_count_4_io_out ? io_r_223_b : _GEN_1512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1514 = 9'he0 == r_count_4_io_out ? io_r_224_b : _GEN_1513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1515 = 9'he1 == r_count_4_io_out ? io_r_225_b : _GEN_1514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1516 = 9'he2 == r_count_4_io_out ? io_r_226_b : _GEN_1515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1517 = 9'he3 == r_count_4_io_out ? io_r_227_b : _GEN_1516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1518 = 9'he4 == r_count_4_io_out ? io_r_228_b : _GEN_1517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1519 = 9'he5 == r_count_4_io_out ? io_r_229_b : _GEN_1518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1520 = 9'he6 == r_count_4_io_out ? io_r_230_b : _GEN_1519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1521 = 9'he7 == r_count_4_io_out ? io_r_231_b : _GEN_1520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1522 = 9'he8 == r_count_4_io_out ? io_r_232_b : _GEN_1521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1523 = 9'he9 == r_count_4_io_out ? io_r_233_b : _GEN_1522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1524 = 9'hea == r_count_4_io_out ? io_r_234_b : _GEN_1523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1525 = 9'heb == r_count_4_io_out ? io_r_235_b : _GEN_1524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1526 = 9'hec == r_count_4_io_out ? io_r_236_b : _GEN_1525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1527 = 9'hed == r_count_4_io_out ? io_r_237_b : _GEN_1526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1528 = 9'hee == r_count_4_io_out ? io_r_238_b : _GEN_1527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1529 = 9'hef == r_count_4_io_out ? io_r_239_b : _GEN_1528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1530 = 9'hf0 == r_count_4_io_out ? io_r_240_b : _GEN_1529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1531 = 9'hf1 == r_count_4_io_out ? io_r_241_b : _GEN_1530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1532 = 9'hf2 == r_count_4_io_out ? io_r_242_b : _GEN_1531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1533 = 9'hf3 == r_count_4_io_out ? io_r_243_b : _GEN_1532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1534 = 9'hf4 == r_count_4_io_out ? io_r_244_b : _GEN_1533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1535 = 9'hf5 == r_count_4_io_out ? io_r_245_b : _GEN_1534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1536 = 9'hf6 == r_count_4_io_out ? io_r_246_b : _GEN_1535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1537 = 9'hf7 == r_count_4_io_out ? io_r_247_b : _GEN_1536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1538 = 9'hf8 == r_count_4_io_out ? io_r_248_b : _GEN_1537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1539 = 9'hf9 == r_count_4_io_out ? io_r_249_b : _GEN_1538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1540 = 9'hfa == r_count_4_io_out ? io_r_250_b : _GEN_1539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1541 = 9'hfb == r_count_4_io_out ? io_r_251_b : _GEN_1540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1542 = 9'hfc == r_count_4_io_out ? io_r_252_b : _GEN_1541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1543 = 9'hfd == r_count_4_io_out ? io_r_253_b : _GEN_1542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1544 = 9'hfe == r_count_4_io_out ? io_r_254_b : _GEN_1543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1545 = 9'hff == r_count_4_io_out ? io_r_255_b : _GEN_1544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1546 = 9'h100 == r_count_4_io_out ? io_r_256_b : _GEN_1545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1547 = 9'h101 == r_count_4_io_out ? io_r_257_b : _GEN_1546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1548 = 9'h102 == r_count_4_io_out ? io_r_258_b : _GEN_1547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1549 = 9'h103 == r_count_4_io_out ? io_r_259_b : _GEN_1548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1550 = 9'h104 == r_count_4_io_out ? io_r_260_b : _GEN_1549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1551 = 9'h105 == r_count_4_io_out ? io_r_261_b : _GEN_1550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1552 = 9'h106 == r_count_4_io_out ? io_r_262_b : _GEN_1551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1553 = 9'h107 == r_count_4_io_out ? io_r_263_b : _GEN_1552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1554 = 9'h108 == r_count_4_io_out ? io_r_264_b : _GEN_1553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1555 = 9'h109 == r_count_4_io_out ? io_r_265_b : _GEN_1554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1556 = 9'h10a == r_count_4_io_out ? io_r_266_b : _GEN_1555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1557 = 9'h10b == r_count_4_io_out ? io_r_267_b : _GEN_1556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1558 = 9'h10c == r_count_4_io_out ? io_r_268_b : _GEN_1557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1559 = 9'h10d == r_count_4_io_out ? io_r_269_b : _GEN_1558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1560 = 9'h10e == r_count_4_io_out ? io_r_270_b : _GEN_1559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1561 = 9'h10f == r_count_4_io_out ? io_r_271_b : _GEN_1560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1562 = 9'h110 == r_count_4_io_out ? io_r_272_b : _GEN_1561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1563 = 9'h111 == r_count_4_io_out ? io_r_273_b : _GEN_1562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1564 = 9'h112 == r_count_4_io_out ? io_r_274_b : _GEN_1563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1565 = 9'h113 == r_count_4_io_out ? io_r_275_b : _GEN_1564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1566 = 9'h114 == r_count_4_io_out ? io_r_276_b : _GEN_1565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1567 = 9'h115 == r_count_4_io_out ? io_r_277_b : _GEN_1566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1568 = 9'h116 == r_count_4_io_out ? io_r_278_b : _GEN_1567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1569 = 9'h117 == r_count_4_io_out ? io_r_279_b : _GEN_1568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1570 = 9'h118 == r_count_4_io_out ? io_r_280_b : _GEN_1569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1571 = 9'h119 == r_count_4_io_out ? io_r_281_b : _GEN_1570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1572 = 9'h11a == r_count_4_io_out ? io_r_282_b : _GEN_1571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1573 = 9'h11b == r_count_4_io_out ? io_r_283_b : _GEN_1572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1574 = 9'h11c == r_count_4_io_out ? io_r_284_b : _GEN_1573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1575 = 9'h11d == r_count_4_io_out ? io_r_285_b : _GEN_1574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1576 = 9'h11e == r_count_4_io_out ? io_r_286_b : _GEN_1575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1577 = 9'h11f == r_count_4_io_out ? io_r_287_b : _GEN_1576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1578 = 9'h120 == r_count_4_io_out ? io_r_288_b : _GEN_1577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1579 = 9'h121 == r_count_4_io_out ? io_r_289_b : _GEN_1578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1580 = 9'h122 == r_count_4_io_out ? io_r_290_b : _GEN_1579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1581 = 9'h123 == r_count_4_io_out ? io_r_291_b : _GEN_1580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1582 = 9'h124 == r_count_4_io_out ? io_r_292_b : _GEN_1581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1583 = 9'h125 == r_count_4_io_out ? io_r_293_b : _GEN_1582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1584 = 9'h126 == r_count_4_io_out ? io_r_294_b : _GEN_1583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1585 = 9'h127 == r_count_4_io_out ? io_r_295_b : _GEN_1584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1586 = 9'h128 == r_count_4_io_out ? io_r_296_b : _GEN_1585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1587 = 9'h129 == r_count_4_io_out ? io_r_297_b : _GEN_1586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1588 = 9'h12a == r_count_4_io_out ? io_r_298_b : _GEN_1587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1591 = 9'h1 == r_count_5_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1592 = 9'h2 == r_count_5_io_out ? io_r_2_b : _GEN_1591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1593 = 9'h3 == r_count_5_io_out ? io_r_3_b : _GEN_1592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1594 = 9'h4 == r_count_5_io_out ? io_r_4_b : _GEN_1593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1595 = 9'h5 == r_count_5_io_out ? io_r_5_b : _GEN_1594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1596 = 9'h6 == r_count_5_io_out ? io_r_6_b : _GEN_1595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1597 = 9'h7 == r_count_5_io_out ? io_r_7_b : _GEN_1596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1598 = 9'h8 == r_count_5_io_out ? io_r_8_b : _GEN_1597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1599 = 9'h9 == r_count_5_io_out ? io_r_9_b : _GEN_1598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1600 = 9'ha == r_count_5_io_out ? io_r_10_b : _GEN_1599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1601 = 9'hb == r_count_5_io_out ? io_r_11_b : _GEN_1600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1602 = 9'hc == r_count_5_io_out ? io_r_12_b : _GEN_1601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1603 = 9'hd == r_count_5_io_out ? io_r_13_b : _GEN_1602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1604 = 9'he == r_count_5_io_out ? io_r_14_b : _GEN_1603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1605 = 9'hf == r_count_5_io_out ? io_r_15_b : _GEN_1604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1606 = 9'h10 == r_count_5_io_out ? io_r_16_b : _GEN_1605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1607 = 9'h11 == r_count_5_io_out ? io_r_17_b : _GEN_1606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1608 = 9'h12 == r_count_5_io_out ? io_r_18_b : _GEN_1607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1609 = 9'h13 == r_count_5_io_out ? io_r_19_b : _GEN_1608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1610 = 9'h14 == r_count_5_io_out ? io_r_20_b : _GEN_1609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1611 = 9'h15 == r_count_5_io_out ? io_r_21_b : _GEN_1610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1612 = 9'h16 == r_count_5_io_out ? io_r_22_b : _GEN_1611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1613 = 9'h17 == r_count_5_io_out ? io_r_23_b : _GEN_1612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1614 = 9'h18 == r_count_5_io_out ? io_r_24_b : _GEN_1613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1615 = 9'h19 == r_count_5_io_out ? io_r_25_b : _GEN_1614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1616 = 9'h1a == r_count_5_io_out ? io_r_26_b : _GEN_1615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1617 = 9'h1b == r_count_5_io_out ? io_r_27_b : _GEN_1616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1618 = 9'h1c == r_count_5_io_out ? io_r_28_b : _GEN_1617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1619 = 9'h1d == r_count_5_io_out ? io_r_29_b : _GEN_1618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1620 = 9'h1e == r_count_5_io_out ? io_r_30_b : _GEN_1619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1621 = 9'h1f == r_count_5_io_out ? io_r_31_b : _GEN_1620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1622 = 9'h20 == r_count_5_io_out ? io_r_32_b : _GEN_1621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1623 = 9'h21 == r_count_5_io_out ? io_r_33_b : _GEN_1622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1624 = 9'h22 == r_count_5_io_out ? io_r_34_b : _GEN_1623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1625 = 9'h23 == r_count_5_io_out ? io_r_35_b : _GEN_1624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1626 = 9'h24 == r_count_5_io_out ? io_r_36_b : _GEN_1625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1627 = 9'h25 == r_count_5_io_out ? io_r_37_b : _GEN_1626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1628 = 9'h26 == r_count_5_io_out ? io_r_38_b : _GEN_1627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1629 = 9'h27 == r_count_5_io_out ? io_r_39_b : _GEN_1628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1630 = 9'h28 == r_count_5_io_out ? io_r_40_b : _GEN_1629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1631 = 9'h29 == r_count_5_io_out ? io_r_41_b : _GEN_1630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1632 = 9'h2a == r_count_5_io_out ? io_r_42_b : _GEN_1631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1633 = 9'h2b == r_count_5_io_out ? io_r_43_b : _GEN_1632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1634 = 9'h2c == r_count_5_io_out ? io_r_44_b : _GEN_1633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1635 = 9'h2d == r_count_5_io_out ? io_r_45_b : _GEN_1634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1636 = 9'h2e == r_count_5_io_out ? io_r_46_b : _GEN_1635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1637 = 9'h2f == r_count_5_io_out ? io_r_47_b : _GEN_1636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1638 = 9'h30 == r_count_5_io_out ? io_r_48_b : _GEN_1637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1639 = 9'h31 == r_count_5_io_out ? io_r_49_b : _GEN_1638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1640 = 9'h32 == r_count_5_io_out ? io_r_50_b : _GEN_1639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1641 = 9'h33 == r_count_5_io_out ? io_r_51_b : _GEN_1640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1642 = 9'h34 == r_count_5_io_out ? io_r_52_b : _GEN_1641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1643 = 9'h35 == r_count_5_io_out ? io_r_53_b : _GEN_1642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1644 = 9'h36 == r_count_5_io_out ? io_r_54_b : _GEN_1643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1645 = 9'h37 == r_count_5_io_out ? io_r_55_b : _GEN_1644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1646 = 9'h38 == r_count_5_io_out ? io_r_56_b : _GEN_1645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1647 = 9'h39 == r_count_5_io_out ? io_r_57_b : _GEN_1646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1648 = 9'h3a == r_count_5_io_out ? io_r_58_b : _GEN_1647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1649 = 9'h3b == r_count_5_io_out ? io_r_59_b : _GEN_1648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1650 = 9'h3c == r_count_5_io_out ? io_r_60_b : _GEN_1649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1651 = 9'h3d == r_count_5_io_out ? io_r_61_b : _GEN_1650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1652 = 9'h3e == r_count_5_io_out ? io_r_62_b : _GEN_1651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1653 = 9'h3f == r_count_5_io_out ? io_r_63_b : _GEN_1652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1654 = 9'h40 == r_count_5_io_out ? io_r_64_b : _GEN_1653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1655 = 9'h41 == r_count_5_io_out ? io_r_65_b : _GEN_1654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1656 = 9'h42 == r_count_5_io_out ? io_r_66_b : _GEN_1655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1657 = 9'h43 == r_count_5_io_out ? io_r_67_b : _GEN_1656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1658 = 9'h44 == r_count_5_io_out ? io_r_68_b : _GEN_1657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1659 = 9'h45 == r_count_5_io_out ? io_r_69_b : _GEN_1658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1660 = 9'h46 == r_count_5_io_out ? io_r_70_b : _GEN_1659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1661 = 9'h47 == r_count_5_io_out ? io_r_71_b : _GEN_1660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1662 = 9'h48 == r_count_5_io_out ? io_r_72_b : _GEN_1661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1663 = 9'h49 == r_count_5_io_out ? io_r_73_b : _GEN_1662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1664 = 9'h4a == r_count_5_io_out ? io_r_74_b : _GEN_1663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1665 = 9'h4b == r_count_5_io_out ? io_r_75_b : _GEN_1664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1666 = 9'h4c == r_count_5_io_out ? io_r_76_b : _GEN_1665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1667 = 9'h4d == r_count_5_io_out ? io_r_77_b : _GEN_1666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1668 = 9'h4e == r_count_5_io_out ? io_r_78_b : _GEN_1667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1669 = 9'h4f == r_count_5_io_out ? io_r_79_b : _GEN_1668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1670 = 9'h50 == r_count_5_io_out ? io_r_80_b : _GEN_1669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1671 = 9'h51 == r_count_5_io_out ? io_r_81_b : _GEN_1670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1672 = 9'h52 == r_count_5_io_out ? io_r_82_b : _GEN_1671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1673 = 9'h53 == r_count_5_io_out ? io_r_83_b : _GEN_1672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1674 = 9'h54 == r_count_5_io_out ? io_r_84_b : _GEN_1673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1675 = 9'h55 == r_count_5_io_out ? io_r_85_b : _GEN_1674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1676 = 9'h56 == r_count_5_io_out ? io_r_86_b : _GEN_1675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1677 = 9'h57 == r_count_5_io_out ? io_r_87_b : _GEN_1676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1678 = 9'h58 == r_count_5_io_out ? io_r_88_b : _GEN_1677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1679 = 9'h59 == r_count_5_io_out ? io_r_89_b : _GEN_1678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1680 = 9'h5a == r_count_5_io_out ? io_r_90_b : _GEN_1679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1681 = 9'h5b == r_count_5_io_out ? io_r_91_b : _GEN_1680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1682 = 9'h5c == r_count_5_io_out ? io_r_92_b : _GEN_1681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1683 = 9'h5d == r_count_5_io_out ? io_r_93_b : _GEN_1682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1684 = 9'h5e == r_count_5_io_out ? io_r_94_b : _GEN_1683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1685 = 9'h5f == r_count_5_io_out ? io_r_95_b : _GEN_1684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1686 = 9'h60 == r_count_5_io_out ? io_r_96_b : _GEN_1685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1687 = 9'h61 == r_count_5_io_out ? io_r_97_b : _GEN_1686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1688 = 9'h62 == r_count_5_io_out ? io_r_98_b : _GEN_1687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1689 = 9'h63 == r_count_5_io_out ? io_r_99_b : _GEN_1688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1690 = 9'h64 == r_count_5_io_out ? io_r_100_b : _GEN_1689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1691 = 9'h65 == r_count_5_io_out ? io_r_101_b : _GEN_1690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1692 = 9'h66 == r_count_5_io_out ? io_r_102_b : _GEN_1691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1693 = 9'h67 == r_count_5_io_out ? io_r_103_b : _GEN_1692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1694 = 9'h68 == r_count_5_io_out ? io_r_104_b : _GEN_1693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1695 = 9'h69 == r_count_5_io_out ? io_r_105_b : _GEN_1694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1696 = 9'h6a == r_count_5_io_out ? io_r_106_b : _GEN_1695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1697 = 9'h6b == r_count_5_io_out ? io_r_107_b : _GEN_1696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1698 = 9'h6c == r_count_5_io_out ? io_r_108_b : _GEN_1697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1699 = 9'h6d == r_count_5_io_out ? io_r_109_b : _GEN_1698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1700 = 9'h6e == r_count_5_io_out ? io_r_110_b : _GEN_1699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1701 = 9'h6f == r_count_5_io_out ? io_r_111_b : _GEN_1700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1702 = 9'h70 == r_count_5_io_out ? io_r_112_b : _GEN_1701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1703 = 9'h71 == r_count_5_io_out ? io_r_113_b : _GEN_1702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1704 = 9'h72 == r_count_5_io_out ? io_r_114_b : _GEN_1703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1705 = 9'h73 == r_count_5_io_out ? io_r_115_b : _GEN_1704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1706 = 9'h74 == r_count_5_io_out ? io_r_116_b : _GEN_1705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1707 = 9'h75 == r_count_5_io_out ? io_r_117_b : _GEN_1706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1708 = 9'h76 == r_count_5_io_out ? io_r_118_b : _GEN_1707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1709 = 9'h77 == r_count_5_io_out ? io_r_119_b : _GEN_1708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1710 = 9'h78 == r_count_5_io_out ? io_r_120_b : _GEN_1709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1711 = 9'h79 == r_count_5_io_out ? io_r_121_b : _GEN_1710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1712 = 9'h7a == r_count_5_io_out ? io_r_122_b : _GEN_1711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1713 = 9'h7b == r_count_5_io_out ? io_r_123_b : _GEN_1712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1714 = 9'h7c == r_count_5_io_out ? io_r_124_b : _GEN_1713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1715 = 9'h7d == r_count_5_io_out ? io_r_125_b : _GEN_1714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1716 = 9'h7e == r_count_5_io_out ? io_r_126_b : _GEN_1715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1717 = 9'h7f == r_count_5_io_out ? io_r_127_b : _GEN_1716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1718 = 9'h80 == r_count_5_io_out ? io_r_128_b : _GEN_1717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1719 = 9'h81 == r_count_5_io_out ? io_r_129_b : _GEN_1718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1720 = 9'h82 == r_count_5_io_out ? io_r_130_b : _GEN_1719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1721 = 9'h83 == r_count_5_io_out ? io_r_131_b : _GEN_1720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1722 = 9'h84 == r_count_5_io_out ? io_r_132_b : _GEN_1721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1723 = 9'h85 == r_count_5_io_out ? io_r_133_b : _GEN_1722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1724 = 9'h86 == r_count_5_io_out ? io_r_134_b : _GEN_1723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1725 = 9'h87 == r_count_5_io_out ? io_r_135_b : _GEN_1724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1726 = 9'h88 == r_count_5_io_out ? io_r_136_b : _GEN_1725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1727 = 9'h89 == r_count_5_io_out ? io_r_137_b : _GEN_1726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1728 = 9'h8a == r_count_5_io_out ? io_r_138_b : _GEN_1727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1729 = 9'h8b == r_count_5_io_out ? io_r_139_b : _GEN_1728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1730 = 9'h8c == r_count_5_io_out ? io_r_140_b : _GEN_1729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1731 = 9'h8d == r_count_5_io_out ? io_r_141_b : _GEN_1730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1732 = 9'h8e == r_count_5_io_out ? io_r_142_b : _GEN_1731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1733 = 9'h8f == r_count_5_io_out ? io_r_143_b : _GEN_1732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1734 = 9'h90 == r_count_5_io_out ? io_r_144_b : _GEN_1733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1735 = 9'h91 == r_count_5_io_out ? io_r_145_b : _GEN_1734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1736 = 9'h92 == r_count_5_io_out ? io_r_146_b : _GEN_1735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1737 = 9'h93 == r_count_5_io_out ? io_r_147_b : _GEN_1736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1738 = 9'h94 == r_count_5_io_out ? io_r_148_b : _GEN_1737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1739 = 9'h95 == r_count_5_io_out ? io_r_149_b : _GEN_1738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1740 = 9'h96 == r_count_5_io_out ? io_r_150_b : _GEN_1739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1741 = 9'h97 == r_count_5_io_out ? io_r_151_b : _GEN_1740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1742 = 9'h98 == r_count_5_io_out ? io_r_152_b : _GEN_1741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1743 = 9'h99 == r_count_5_io_out ? io_r_153_b : _GEN_1742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1744 = 9'h9a == r_count_5_io_out ? io_r_154_b : _GEN_1743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1745 = 9'h9b == r_count_5_io_out ? io_r_155_b : _GEN_1744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1746 = 9'h9c == r_count_5_io_out ? io_r_156_b : _GEN_1745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1747 = 9'h9d == r_count_5_io_out ? io_r_157_b : _GEN_1746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1748 = 9'h9e == r_count_5_io_out ? io_r_158_b : _GEN_1747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1749 = 9'h9f == r_count_5_io_out ? io_r_159_b : _GEN_1748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1750 = 9'ha0 == r_count_5_io_out ? io_r_160_b : _GEN_1749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1751 = 9'ha1 == r_count_5_io_out ? io_r_161_b : _GEN_1750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1752 = 9'ha2 == r_count_5_io_out ? io_r_162_b : _GEN_1751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1753 = 9'ha3 == r_count_5_io_out ? io_r_163_b : _GEN_1752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1754 = 9'ha4 == r_count_5_io_out ? io_r_164_b : _GEN_1753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1755 = 9'ha5 == r_count_5_io_out ? io_r_165_b : _GEN_1754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1756 = 9'ha6 == r_count_5_io_out ? io_r_166_b : _GEN_1755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1757 = 9'ha7 == r_count_5_io_out ? io_r_167_b : _GEN_1756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1758 = 9'ha8 == r_count_5_io_out ? io_r_168_b : _GEN_1757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1759 = 9'ha9 == r_count_5_io_out ? io_r_169_b : _GEN_1758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1760 = 9'haa == r_count_5_io_out ? io_r_170_b : _GEN_1759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1761 = 9'hab == r_count_5_io_out ? io_r_171_b : _GEN_1760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1762 = 9'hac == r_count_5_io_out ? io_r_172_b : _GEN_1761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1763 = 9'had == r_count_5_io_out ? io_r_173_b : _GEN_1762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1764 = 9'hae == r_count_5_io_out ? io_r_174_b : _GEN_1763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1765 = 9'haf == r_count_5_io_out ? io_r_175_b : _GEN_1764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1766 = 9'hb0 == r_count_5_io_out ? io_r_176_b : _GEN_1765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1767 = 9'hb1 == r_count_5_io_out ? io_r_177_b : _GEN_1766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1768 = 9'hb2 == r_count_5_io_out ? io_r_178_b : _GEN_1767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1769 = 9'hb3 == r_count_5_io_out ? io_r_179_b : _GEN_1768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1770 = 9'hb4 == r_count_5_io_out ? io_r_180_b : _GEN_1769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1771 = 9'hb5 == r_count_5_io_out ? io_r_181_b : _GEN_1770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1772 = 9'hb6 == r_count_5_io_out ? io_r_182_b : _GEN_1771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1773 = 9'hb7 == r_count_5_io_out ? io_r_183_b : _GEN_1772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1774 = 9'hb8 == r_count_5_io_out ? io_r_184_b : _GEN_1773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1775 = 9'hb9 == r_count_5_io_out ? io_r_185_b : _GEN_1774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1776 = 9'hba == r_count_5_io_out ? io_r_186_b : _GEN_1775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1777 = 9'hbb == r_count_5_io_out ? io_r_187_b : _GEN_1776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1778 = 9'hbc == r_count_5_io_out ? io_r_188_b : _GEN_1777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1779 = 9'hbd == r_count_5_io_out ? io_r_189_b : _GEN_1778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1780 = 9'hbe == r_count_5_io_out ? io_r_190_b : _GEN_1779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1781 = 9'hbf == r_count_5_io_out ? io_r_191_b : _GEN_1780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1782 = 9'hc0 == r_count_5_io_out ? io_r_192_b : _GEN_1781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1783 = 9'hc1 == r_count_5_io_out ? io_r_193_b : _GEN_1782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1784 = 9'hc2 == r_count_5_io_out ? io_r_194_b : _GEN_1783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1785 = 9'hc3 == r_count_5_io_out ? io_r_195_b : _GEN_1784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1786 = 9'hc4 == r_count_5_io_out ? io_r_196_b : _GEN_1785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1787 = 9'hc5 == r_count_5_io_out ? io_r_197_b : _GEN_1786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1788 = 9'hc6 == r_count_5_io_out ? io_r_198_b : _GEN_1787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1789 = 9'hc7 == r_count_5_io_out ? io_r_199_b : _GEN_1788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1790 = 9'hc8 == r_count_5_io_out ? io_r_200_b : _GEN_1789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1791 = 9'hc9 == r_count_5_io_out ? io_r_201_b : _GEN_1790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1792 = 9'hca == r_count_5_io_out ? io_r_202_b : _GEN_1791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1793 = 9'hcb == r_count_5_io_out ? io_r_203_b : _GEN_1792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1794 = 9'hcc == r_count_5_io_out ? io_r_204_b : _GEN_1793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1795 = 9'hcd == r_count_5_io_out ? io_r_205_b : _GEN_1794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1796 = 9'hce == r_count_5_io_out ? io_r_206_b : _GEN_1795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1797 = 9'hcf == r_count_5_io_out ? io_r_207_b : _GEN_1796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1798 = 9'hd0 == r_count_5_io_out ? io_r_208_b : _GEN_1797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1799 = 9'hd1 == r_count_5_io_out ? io_r_209_b : _GEN_1798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1800 = 9'hd2 == r_count_5_io_out ? io_r_210_b : _GEN_1799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1801 = 9'hd3 == r_count_5_io_out ? io_r_211_b : _GEN_1800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1802 = 9'hd4 == r_count_5_io_out ? io_r_212_b : _GEN_1801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1803 = 9'hd5 == r_count_5_io_out ? io_r_213_b : _GEN_1802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1804 = 9'hd6 == r_count_5_io_out ? io_r_214_b : _GEN_1803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1805 = 9'hd7 == r_count_5_io_out ? io_r_215_b : _GEN_1804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1806 = 9'hd8 == r_count_5_io_out ? io_r_216_b : _GEN_1805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1807 = 9'hd9 == r_count_5_io_out ? io_r_217_b : _GEN_1806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1808 = 9'hda == r_count_5_io_out ? io_r_218_b : _GEN_1807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1809 = 9'hdb == r_count_5_io_out ? io_r_219_b : _GEN_1808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1810 = 9'hdc == r_count_5_io_out ? io_r_220_b : _GEN_1809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1811 = 9'hdd == r_count_5_io_out ? io_r_221_b : _GEN_1810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1812 = 9'hde == r_count_5_io_out ? io_r_222_b : _GEN_1811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1813 = 9'hdf == r_count_5_io_out ? io_r_223_b : _GEN_1812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1814 = 9'he0 == r_count_5_io_out ? io_r_224_b : _GEN_1813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1815 = 9'he1 == r_count_5_io_out ? io_r_225_b : _GEN_1814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1816 = 9'he2 == r_count_5_io_out ? io_r_226_b : _GEN_1815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1817 = 9'he3 == r_count_5_io_out ? io_r_227_b : _GEN_1816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1818 = 9'he4 == r_count_5_io_out ? io_r_228_b : _GEN_1817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1819 = 9'he5 == r_count_5_io_out ? io_r_229_b : _GEN_1818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1820 = 9'he6 == r_count_5_io_out ? io_r_230_b : _GEN_1819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1821 = 9'he7 == r_count_5_io_out ? io_r_231_b : _GEN_1820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1822 = 9'he8 == r_count_5_io_out ? io_r_232_b : _GEN_1821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1823 = 9'he9 == r_count_5_io_out ? io_r_233_b : _GEN_1822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1824 = 9'hea == r_count_5_io_out ? io_r_234_b : _GEN_1823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1825 = 9'heb == r_count_5_io_out ? io_r_235_b : _GEN_1824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1826 = 9'hec == r_count_5_io_out ? io_r_236_b : _GEN_1825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1827 = 9'hed == r_count_5_io_out ? io_r_237_b : _GEN_1826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1828 = 9'hee == r_count_5_io_out ? io_r_238_b : _GEN_1827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1829 = 9'hef == r_count_5_io_out ? io_r_239_b : _GEN_1828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1830 = 9'hf0 == r_count_5_io_out ? io_r_240_b : _GEN_1829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1831 = 9'hf1 == r_count_5_io_out ? io_r_241_b : _GEN_1830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1832 = 9'hf2 == r_count_5_io_out ? io_r_242_b : _GEN_1831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1833 = 9'hf3 == r_count_5_io_out ? io_r_243_b : _GEN_1832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1834 = 9'hf4 == r_count_5_io_out ? io_r_244_b : _GEN_1833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1835 = 9'hf5 == r_count_5_io_out ? io_r_245_b : _GEN_1834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1836 = 9'hf6 == r_count_5_io_out ? io_r_246_b : _GEN_1835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1837 = 9'hf7 == r_count_5_io_out ? io_r_247_b : _GEN_1836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1838 = 9'hf8 == r_count_5_io_out ? io_r_248_b : _GEN_1837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1839 = 9'hf9 == r_count_5_io_out ? io_r_249_b : _GEN_1838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1840 = 9'hfa == r_count_5_io_out ? io_r_250_b : _GEN_1839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1841 = 9'hfb == r_count_5_io_out ? io_r_251_b : _GEN_1840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1842 = 9'hfc == r_count_5_io_out ? io_r_252_b : _GEN_1841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1843 = 9'hfd == r_count_5_io_out ? io_r_253_b : _GEN_1842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1844 = 9'hfe == r_count_5_io_out ? io_r_254_b : _GEN_1843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1845 = 9'hff == r_count_5_io_out ? io_r_255_b : _GEN_1844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1846 = 9'h100 == r_count_5_io_out ? io_r_256_b : _GEN_1845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1847 = 9'h101 == r_count_5_io_out ? io_r_257_b : _GEN_1846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1848 = 9'h102 == r_count_5_io_out ? io_r_258_b : _GEN_1847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1849 = 9'h103 == r_count_5_io_out ? io_r_259_b : _GEN_1848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1850 = 9'h104 == r_count_5_io_out ? io_r_260_b : _GEN_1849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1851 = 9'h105 == r_count_5_io_out ? io_r_261_b : _GEN_1850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1852 = 9'h106 == r_count_5_io_out ? io_r_262_b : _GEN_1851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1853 = 9'h107 == r_count_5_io_out ? io_r_263_b : _GEN_1852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1854 = 9'h108 == r_count_5_io_out ? io_r_264_b : _GEN_1853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1855 = 9'h109 == r_count_5_io_out ? io_r_265_b : _GEN_1854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1856 = 9'h10a == r_count_5_io_out ? io_r_266_b : _GEN_1855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1857 = 9'h10b == r_count_5_io_out ? io_r_267_b : _GEN_1856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1858 = 9'h10c == r_count_5_io_out ? io_r_268_b : _GEN_1857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1859 = 9'h10d == r_count_5_io_out ? io_r_269_b : _GEN_1858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1860 = 9'h10e == r_count_5_io_out ? io_r_270_b : _GEN_1859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1861 = 9'h10f == r_count_5_io_out ? io_r_271_b : _GEN_1860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1862 = 9'h110 == r_count_5_io_out ? io_r_272_b : _GEN_1861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1863 = 9'h111 == r_count_5_io_out ? io_r_273_b : _GEN_1862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1864 = 9'h112 == r_count_5_io_out ? io_r_274_b : _GEN_1863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1865 = 9'h113 == r_count_5_io_out ? io_r_275_b : _GEN_1864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1866 = 9'h114 == r_count_5_io_out ? io_r_276_b : _GEN_1865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1867 = 9'h115 == r_count_5_io_out ? io_r_277_b : _GEN_1866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1868 = 9'h116 == r_count_5_io_out ? io_r_278_b : _GEN_1867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1869 = 9'h117 == r_count_5_io_out ? io_r_279_b : _GEN_1868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1870 = 9'h118 == r_count_5_io_out ? io_r_280_b : _GEN_1869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1871 = 9'h119 == r_count_5_io_out ? io_r_281_b : _GEN_1870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1872 = 9'h11a == r_count_5_io_out ? io_r_282_b : _GEN_1871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1873 = 9'h11b == r_count_5_io_out ? io_r_283_b : _GEN_1872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1874 = 9'h11c == r_count_5_io_out ? io_r_284_b : _GEN_1873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1875 = 9'h11d == r_count_5_io_out ? io_r_285_b : _GEN_1874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1876 = 9'h11e == r_count_5_io_out ? io_r_286_b : _GEN_1875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1877 = 9'h11f == r_count_5_io_out ? io_r_287_b : _GEN_1876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1878 = 9'h120 == r_count_5_io_out ? io_r_288_b : _GEN_1877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1879 = 9'h121 == r_count_5_io_out ? io_r_289_b : _GEN_1878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1880 = 9'h122 == r_count_5_io_out ? io_r_290_b : _GEN_1879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1881 = 9'h123 == r_count_5_io_out ? io_r_291_b : _GEN_1880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1882 = 9'h124 == r_count_5_io_out ? io_r_292_b : _GEN_1881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1883 = 9'h125 == r_count_5_io_out ? io_r_293_b : _GEN_1882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1884 = 9'h126 == r_count_5_io_out ? io_r_294_b : _GEN_1883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1885 = 9'h127 == r_count_5_io_out ? io_r_295_b : _GEN_1884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1886 = 9'h128 == r_count_5_io_out ? io_r_296_b : _GEN_1885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1887 = 9'h129 == r_count_5_io_out ? io_r_297_b : _GEN_1886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1888 = 9'h12a == r_count_5_io_out ? io_r_298_b : _GEN_1887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1891 = 9'h1 == r_count_6_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1892 = 9'h2 == r_count_6_io_out ? io_r_2_b : _GEN_1891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1893 = 9'h3 == r_count_6_io_out ? io_r_3_b : _GEN_1892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1894 = 9'h4 == r_count_6_io_out ? io_r_4_b : _GEN_1893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1895 = 9'h5 == r_count_6_io_out ? io_r_5_b : _GEN_1894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1896 = 9'h6 == r_count_6_io_out ? io_r_6_b : _GEN_1895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1897 = 9'h7 == r_count_6_io_out ? io_r_7_b : _GEN_1896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1898 = 9'h8 == r_count_6_io_out ? io_r_8_b : _GEN_1897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1899 = 9'h9 == r_count_6_io_out ? io_r_9_b : _GEN_1898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1900 = 9'ha == r_count_6_io_out ? io_r_10_b : _GEN_1899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1901 = 9'hb == r_count_6_io_out ? io_r_11_b : _GEN_1900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1902 = 9'hc == r_count_6_io_out ? io_r_12_b : _GEN_1901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1903 = 9'hd == r_count_6_io_out ? io_r_13_b : _GEN_1902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1904 = 9'he == r_count_6_io_out ? io_r_14_b : _GEN_1903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1905 = 9'hf == r_count_6_io_out ? io_r_15_b : _GEN_1904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1906 = 9'h10 == r_count_6_io_out ? io_r_16_b : _GEN_1905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1907 = 9'h11 == r_count_6_io_out ? io_r_17_b : _GEN_1906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1908 = 9'h12 == r_count_6_io_out ? io_r_18_b : _GEN_1907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1909 = 9'h13 == r_count_6_io_out ? io_r_19_b : _GEN_1908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1910 = 9'h14 == r_count_6_io_out ? io_r_20_b : _GEN_1909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1911 = 9'h15 == r_count_6_io_out ? io_r_21_b : _GEN_1910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1912 = 9'h16 == r_count_6_io_out ? io_r_22_b : _GEN_1911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1913 = 9'h17 == r_count_6_io_out ? io_r_23_b : _GEN_1912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1914 = 9'h18 == r_count_6_io_out ? io_r_24_b : _GEN_1913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1915 = 9'h19 == r_count_6_io_out ? io_r_25_b : _GEN_1914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1916 = 9'h1a == r_count_6_io_out ? io_r_26_b : _GEN_1915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1917 = 9'h1b == r_count_6_io_out ? io_r_27_b : _GEN_1916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1918 = 9'h1c == r_count_6_io_out ? io_r_28_b : _GEN_1917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1919 = 9'h1d == r_count_6_io_out ? io_r_29_b : _GEN_1918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1920 = 9'h1e == r_count_6_io_out ? io_r_30_b : _GEN_1919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1921 = 9'h1f == r_count_6_io_out ? io_r_31_b : _GEN_1920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1922 = 9'h20 == r_count_6_io_out ? io_r_32_b : _GEN_1921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1923 = 9'h21 == r_count_6_io_out ? io_r_33_b : _GEN_1922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1924 = 9'h22 == r_count_6_io_out ? io_r_34_b : _GEN_1923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1925 = 9'h23 == r_count_6_io_out ? io_r_35_b : _GEN_1924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1926 = 9'h24 == r_count_6_io_out ? io_r_36_b : _GEN_1925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1927 = 9'h25 == r_count_6_io_out ? io_r_37_b : _GEN_1926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1928 = 9'h26 == r_count_6_io_out ? io_r_38_b : _GEN_1927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1929 = 9'h27 == r_count_6_io_out ? io_r_39_b : _GEN_1928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1930 = 9'h28 == r_count_6_io_out ? io_r_40_b : _GEN_1929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1931 = 9'h29 == r_count_6_io_out ? io_r_41_b : _GEN_1930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1932 = 9'h2a == r_count_6_io_out ? io_r_42_b : _GEN_1931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1933 = 9'h2b == r_count_6_io_out ? io_r_43_b : _GEN_1932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1934 = 9'h2c == r_count_6_io_out ? io_r_44_b : _GEN_1933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1935 = 9'h2d == r_count_6_io_out ? io_r_45_b : _GEN_1934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1936 = 9'h2e == r_count_6_io_out ? io_r_46_b : _GEN_1935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1937 = 9'h2f == r_count_6_io_out ? io_r_47_b : _GEN_1936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1938 = 9'h30 == r_count_6_io_out ? io_r_48_b : _GEN_1937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1939 = 9'h31 == r_count_6_io_out ? io_r_49_b : _GEN_1938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1940 = 9'h32 == r_count_6_io_out ? io_r_50_b : _GEN_1939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1941 = 9'h33 == r_count_6_io_out ? io_r_51_b : _GEN_1940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1942 = 9'h34 == r_count_6_io_out ? io_r_52_b : _GEN_1941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1943 = 9'h35 == r_count_6_io_out ? io_r_53_b : _GEN_1942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1944 = 9'h36 == r_count_6_io_out ? io_r_54_b : _GEN_1943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1945 = 9'h37 == r_count_6_io_out ? io_r_55_b : _GEN_1944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1946 = 9'h38 == r_count_6_io_out ? io_r_56_b : _GEN_1945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1947 = 9'h39 == r_count_6_io_out ? io_r_57_b : _GEN_1946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1948 = 9'h3a == r_count_6_io_out ? io_r_58_b : _GEN_1947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1949 = 9'h3b == r_count_6_io_out ? io_r_59_b : _GEN_1948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1950 = 9'h3c == r_count_6_io_out ? io_r_60_b : _GEN_1949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1951 = 9'h3d == r_count_6_io_out ? io_r_61_b : _GEN_1950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1952 = 9'h3e == r_count_6_io_out ? io_r_62_b : _GEN_1951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1953 = 9'h3f == r_count_6_io_out ? io_r_63_b : _GEN_1952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1954 = 9'h40 == r_count_6_io_out ? io_r_64_b : _GEN_1953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1955 = 9'h41 == r_count_6_io_out ? io_r_65_b : _GEN_1954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1956 = 9'h42 == r_count_6_io_out ? io_r_66_b : _GEN_1955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1957 = 9'h43 == r_count_6_io_out ? io_r_67_b : _GEN_1956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1958 = 9'h44 == r_count_6_io_out ? io_r_68_b : _GEN_1957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1959 = 9'h45 == r_count_6_io_out ? io_r_69_b : _GEN_1958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1960 = 9'h46 == r_count_6_io_out ? io_r_70_b : _GEN_1959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1961 = 9'h47 == r_count_6_io_out ? io_r_71_b : _GEN_1960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1962 = 9'h48 == r_count_6_io_out ? io_r_72_b : _GEN_1961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1963 = 9'h49 == r_count_6_io_out ? io_r_73_b : _GEN_1962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1964 = 9'h4a == r_count_6_io_out ? io_r_74_b : _GEN_1963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1965 = 9'h4b == r_count_6_io_out ? io_r_75_b : _GEN_1964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1966 = 9'h4c == r_count_6_io_out ? io_r_76_b : _GEN_1965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1967 = 9'h4d == r_count_6_io_out ? io_r_77_b : _GEN_1966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1968 = 9'h4e == r_count_6_io_out ? io_r_78_b : _GEN_1967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1969 = 9'h4f == r_count_6_io_out ? io_r_79_b : _GEN_1968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1970 = 9'h50 == r_count_6_io_out ? io_r_80_b : _GEN_1969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1971 = 9'h51 == r_count_6_io_out ? io_r_81_b : _GEN_1970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1972 = 9'h52 == r_count_6_io_out ? io_r_82_b : _GEN_1971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1973 = 9'h53 == r_count_6_io_out ? io_r_83_b : _GEN_1972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1974 = 9'h54 == r_count_6_io_out ? io_r_84_b : _GEN_1973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1975 = 9'h55 == r_count_6_io_out ? io_r_85_b : _GEN_1974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1976 = 9'h56 == r_count_6_io_out ? io_r_86_b : _GEN_1975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1977 = 9'h57 == r_count_6_io_out ? io_r_87_b : _GEN_1976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1978 = 9'h58 == r_count_6_io_out ? io_r_88_b : _GEN_1977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1979 = 9'h59 == r_count_6_io_out ? io_r_89_b : _GEN_1978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1980 = 9'h5a == r_count_6_io_out ? io_r_90_b : _GEN_1979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1981 = 9'h5b == r_count_6_io_out ? io_r_91_b : _GEN_1980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1982 = 9'h5c == r_count_6_io_out ? io_r_92_b : _GEN_1981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1983 = 9'h5d == r_count_6_io_out ? io_r_93_b : _GEN_1982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1984 = 9'h5e == r_count_6_io_out ? io_r_94_b : _GEN_1983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1985 = 9'h5f == r_count_6_io_out ? io_r_95_b : _GEN_1984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1986 = 9'h60 == r_count_6_io_out ? io_r_96_b : _GEN_1985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1987 = 9'h61 == r_count_6_io_out ? io_r_97_b : _GEN_1986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1988 = 9'h62 == r_count_6_io_out ? io_r_98_b : _GEN_1987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1989 = 9'h63 == r_count_6_io_out ? io_r_99_b : _GEN_1988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1990 = 9'h64 == r_count_6_io_out ? io_r_100_b : _GEN_1989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1991 = 9'h65 == r_count_6_io_out ? io_r_101_b : _GEN_1990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1992 = 9'h66 == r_count_6_io_out ? io_r_102_b : _GEN_1991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1993 = 9'h67 == r_count_6_io_out ? io_r_103_b : _GEN_1992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1994 = 9'h68 == r_count_6_io_out ? io_r_104_b : _GEN_1993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1995 = 9'h69 == r_count_6_io_out ? io_r_105_b : _GEN_1994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1996 = 9'h6a == r_count_6_io_out ? io_r_106_b : _GEN_1995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1997 = 9'h6b == r_count_6_io_out ? io_r_107_b : _GEN_1996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1998 = 9'h6c == r_count_6_io_out ? io_r_108_b : _GEN_1997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1999 = 9'h6d == r_count_6_io_out ? io_r_109_b : _GEN_1998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2000 = 9'h6e == r_count_6_io_out ? io_r_110_b : _GEN_1999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2001 = 9'h6f == r_count_6_io_out ? io_r_111_b : _GEN_2000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2002 = 9'h70 == r_count_6_io_out ? io_r_112_b : _GEN_2001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2003 = 9'h71 == r_count_6_io_out ? io_r_113_b : _GEN_2002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2004 = 9'h72 == r_count_6_io_out ? io_r_114_b : _GEN_2003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2005 = 9'h73 == r_count_6_io_out ? io_r_115_b : _GEN_2004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2006 = 9'h74 == r_count_6_io_out ? io_r_116_b : _GEN_2005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2007 = 9'h75 == r_count_6_io_out ? io_r_117_b : _GEN_2006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2008 = 9'h76 == r_count_6_io_out ? io_r_118_b : _GEN_2007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2009 = 9'h77 == r_count_6_io_out ? io_r_119_b : _GEN_2008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2010 = 9'h78 == r_count_6_io_out ? io_r_120_b : _GEN_2009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2011 = 9'h79 == r_count_6_io_out ? io_r_121_b : _GEN_2010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2012 = 9'h7a == r_count_6_io_out ? io_r_122_b : _GEN_2011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2013 = 9'h7b == r_count_6_io_out ? io_r_123_b : _GEN_2012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2014 = 9'h7c == r_count_6_io_out ? io_r_124_b : _GEN_2013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2015 = 9'h7d == r_count_6_io_out ? io_r_125_b : _GEN_2014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2016 = 9'h7e == r_count_6_io_out ? io_r_126_b : _GEN_2015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2017 = 9'h7f == r_count_6_io_out ? io_r_127_b : _GEN_2016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2018 = 9'h80 == r_count_6_io_out ? io_r_128_b : _GEN_2017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2019 = 9'h81 == r_count_6_io_out ? io_r_129_b : _GEN_2018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2020 = 9'h82 == r_count_6_io_out ? io_r_130_b : _GEN_2019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2021 = 9'h83 == r_count_6_io_out ? io_r_131_b : _GEN_2020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2022 = 9'h84 == r_count_6_io_out ? io_r_132_b : _GEN_2021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2023 = 9'h85 == r_count_6_io_out ? io_r_133_b : _GEN_2022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2024 = 9'h86 == r_count_6_io_out ? io_r_134_b : _GEN_2023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2025 = 9'h87 == r_count_6_io_out ? io_r_135_b : _GEN_2024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2026 = 9'h88 == r_count_6_io_out ? io_r_136_b : _GEN_2025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2027 = 9'h89 == r_count_6_io_out ? io_r_137_b : _GEN_2026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2028 = 9'h8a == r_count_6_io_out ? io_r_138_b : _GEN_2027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2029 = 9'h8b == r_count_6_io_out ? io_r_139_b : _GEN_2028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2030 = 9'h8c == r_count_6_io_out ? io_r_140_b : _GEN_2029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2031 = 9'h8d == r_count_6_io_out ? io_r_141_b : _GEN_2030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2032 = 9'h8e == r_count_6_io_out ? io_r_142_b : _GEN_2031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2033 = 9'h8f == r_count_6_io_out ? io_r_143_b : _GEN_2032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2034 = 9'h90 == r_count_6_io_out ? io_r_144_b : _GEN_2033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2035 = 9'h91 == r_count_6_io_out ? io_r_145_b : _GEN_2034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2036 = 9'h92 == r_count_6_io_out ? io_r_146_b : _GEN_2035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2037 = 9'h93 == r_count_6_io_out ? io_r_147_b : _GEN_2036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2038 = 9'h94 == r_count_6_io_out ? io_r_148_b : _GEN_2037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2039 = 9'h95 == r_count_6_io_out ? io_r_149_b : _GEN_2038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2040 = 9'h96 == r_count_6_io_out ? io_r_150_b : _GEN_2039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2041 = 9'h97 == r_count_6_io_out ? io_r_151_b : _GEN_2040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2042 = 9'h98 == r_count_6_io_out ? io_r_152_b : _GEN_2041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2043 = 9'h99 == r_count_6_io_out ? io_r_153_b : _GEN_2042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2044 = 9'h9a == r_count_6_io_out ? io_r_154_b : _GEN_2043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2045 = 9'h9b == r_count_6_io_out ? io_r_155_b : _GEN_2044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2046 = 9'h9c == r_count_6_io_out ? io_r_156_b : _GEN_2045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2047 = 9'h9d == r_count_6_io_out ? io_r_157_b : _GEN_2046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2048 = 9'h9e == r_count_6_io_out ? io_r_158_b : _GEN_2047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2049 = 9'h9f == r_count_6_io_out ? io_r_159_b : _GEN_2048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2050 = 9'ha0 == r_count_6_io_out ? io_r_160_b : _GEN_2049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2051 = 9'ha1 == r_count_6_io_out ? io_r_161_b : _GEN_2050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2052 = 9'ha2 == r_count_6_io_out ? io_r_162_b : _GEN_2051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2053 = 9'ha3 == r_count_6_io_out ? io_r_163_b : _GEN_2052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2054 = 9'ha4 == r_count_6_io_out ? io_r_164_b : _GEN_2053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2055 = 9'ha5 == r_count_6_io_out ? io_r_165_b : _GEN_2054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2056 = 9'ha6 == r_count_6_io_out ? io_r_166_b : _GEN_2055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2057 = 9'ha7 == r_count_6_io_out ? io_r_167_b : _GEN_2056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2058 = 9'ha8 == r_count_6_io_out ? io_r_168_b : _GEN_2057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2059 = 9'ha9 == r_count_6_io_out ? io_r_169_b : _GEN_2058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2060 = 9'haa == r_count_6_io_out ? io_r_170_b : _GEN_2059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2061 = 9'hab == r_count_6_io_out ? io_r_171_b : _GEN_2060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2062 = 9'hac == r_count_6_io_out ? io_r_172_b : _GEN_2061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2063 = 9'had == r_count_6_io_out ? io_r_173_b : _GEN_2062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2064 = 9'hae == r_count_6_io_out ? io_r_174_b : _GEN_2063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2065 = 9'haf == r_count_6_io_out ? io_r_175_b : _GEN_2064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2066 = 9'hb0 == r_count_6_io_out ? io_r_176_b : _GEN_2065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2067 = 9'hb1 == r_count_6_io_out ? io_r_177_b : _GEN_2066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2068 = 9'hb2 == r_count_6_io_out ? io_r_178_b : _GEN_2067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2069 = 9'hb3 == r_count_6_io_out ? io_r_179_b : _GEN_2068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2070 = 9'hb4 == r_count_6_io_out ? io_r_180_b : _GEN_2069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2071 = 9'hb5 == r_count_6_io_out ? io_r_181_b : _GEN_2070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2072 = 9'hb6 == r_count_6_io_out ? io_r_182_b : _GEN_2071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2073 = 9'hb7 == r_count_6_io_out ? io_r_183_b : _GEN_2072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2074 = 9'hb8 == r_count_6_io_out ? io_r_184_b : _GEN_2073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2075 = 9'hb9 == r_count_6_io_out ? io_r_185_b : _GEN_2074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2076 = 9'hba == r_count_6_io_out ? io_r_186_b : _GEN_2075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2077 = 9'hbb == r_count_6_io_out ? io_r_187_b : _GEN_2076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2078 = 9'hbc == r_count_6_io_out ? io_r_188_b : _GEN_2077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2079 = 9'hbd == r_count_6_io_out ? io_r_189_b : _GEN_2078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2080 = 9'hbe == r_count_6_io_out ? io_r_190_b : _GEN_2079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2081 = 9'hbf == r_count_6_io_out ? io_r_191_b : _GEN_2080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2082 = 9'hc0 == r_count_6_io_out ? io_r_192_b : _GEN_2081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2083 = 9'hc1 == r_count_6_io_out ? io_r_193_b : _GEN_2082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2084 = 9'hc2 == r_count_6_io_out ? io_r_194_b : _GEN_2083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2085 = 9'hc3 == r_count_6_io_out ? io_r_195_b : _GEN_2084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2086 = 9'hc4 == r_count_6_io_out ? io_r_196_b : _GEN_2085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2087 = 9'hc5 == r_count_6_io_out ? io_r_197_b : _GEN_2086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2088 = 9'hc6 == r_count_6_io_out ? io_r_198_b : _GEN_2087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2089 = 9'hc7 == r_count_6_io_out ? io_r_199_b : _GEN_2088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2090 = 9'hc8 == r_count_6_io_out ? io_r_200_b : _GEN_2089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2091 = 9'hc9 == r_count_6_io_out ? io_r_201_b : _GEN_2090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2092 = 9'hca == r_count_6_io_out ? io_r_202_b : _GEN_2091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2093 = 9'hcb == r_count_6_io_out ? io_r_203_b : _GEN_2092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2094 = 9'hcc == r_count_6_io_out ? io_r_204_b : _GEN_2093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2095 = 9'hcd == r_count_6_io_out ? io_r_205_b : _GEN_2094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2096 = 9'hce == r_count_6_io_out ? io_r_206_b : _GEN_2095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2097 = 9'hcf == r_count_6_io_out ? io_r_207_b : _GEN_2096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2098 = 9'hd0 == r_count_6_io_out ? io_r_208_b : _GEN_2097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2099 = 9'hd1 == r_count_6_io_out ? io_r_209_b : _GEN_2098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2100 = 9'hd2 == r_count_6_io_out ? io_r_210_b : _GEN_2099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2101 = 9'hd3 == r_count_6_io_out ? io_r_211_b : _GEN_2100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2102 = 9'hd4 == r_count_6_io_out ? io_r_212_b : _GEN_2101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2103 = 9'hd5 == r_count_6_io_out ? io_r_213_b : _GEN_2102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2104 = 9'hd6 == r_count_6_io_out ? io_r_214_b : _GEN_2103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2105 = 9'hd7 == r_count_6_io_out ? io_r_215_b : _GEN_2104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2106 = 9'hd8 == r_count_6_io_out ? io_r_216_b : _GEN_2105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2107 = 9'hd9 == r_count_6_io_out ? io_r_217_b : _GEN_2106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2108 = 9'hda == r_count_6_io_out ? io_r_218_b : _GEN_2107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2109 = 9'hdb == r_count_6_io_out ? io_r_219_b : _GEN_2108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2110 = 9'hdc == r_count_6_io_out ? io_r_220_b : _GEN_2109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2111 = 9'hdd == r_count_6_io_out ? io_r_221_b : _GEN_2110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2112 = 9'hde == r_count_6_io_out ? io_r_222_b : _GEN_2111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2113 = 9'hdf == r_count_6_io_out ? io_r_223_b : _GEN_2112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2114 = 9'he0 == r_count_6_io_out ? io_r_224_b : _GEN_2113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2115 = 9'he1 == r_count_6_io_out ? io_r_225_b : _GEN_2114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2116 = 9'he2 == r_count_6_io_out ? io_r_226_b : _GEN_2115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2117 = 9'he3 == r_count_6_io_out ? io_r_227_b : _GEN_2116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2118 = 9'he4 == r_count_6_io_out ? io_r_228_b : _GEN_2117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2119 = 9'he5 == r_count_6_io_out ? io_r_229_b : _GEN_2118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2120 = 9'he6 == r_count_6_io_out ? io_r_230_b : _GEN_2119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2121 = 9'he7 == r_count_6_io_out ? io_r_231_b : _GEN_2120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2122 = 9'he8 == r_count_6_io_out ? io_r_232_b : _GEN_2121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2123 = 9'he9 == r_count_6_io_out ? io_r_233_b : _GEN_2122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2124 = 9'hea == r_count_6_io_out ? io_r_234_b : _GEN_2123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2125 = 9'heb == r_count_6_io_out ? io_r_235_b : _GEN_2124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2126 = 9'hec == r_count_6_io_out ? io_r_236_b : _GEN_2125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2127 = 9'hed == r_count_6_io_out ? io_r_237_b : _GEN_2126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2128 = 9'hee == r_count_6_io_out ? io_r_238_b : _GEN_2127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2129 = 9'hef == r_count_6_io_out ? io_r_239_b : _GEN_2128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2130 = 9'hf0 == r_count_6_io_out ? io_r_240_b : _GEN_2129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2131 = 9'hf1 == r_count_6_io_out ? io_r_241_b : _GEN_2130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2132 = 9'hf2 == r_count_6_io_out ? io_r_242_b : _GEN_2131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2133 = 9'hf3 == r_count_6_io_out ? io_r_243_b : _GEN_2132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2134 = 9'hf4 == r_count_6_io_out ? io_r_244_b : _GEN_2133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2135 = 9'hf5 == r_count_6_io_out ? io_r_245_b : _GEN_2134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2136 = 9'hf6 == r_count_6_io_out ? io_r_246_b : _GEN_2135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2137 = 9'hf7 == r_count_6_io_out ? io_r_247_b : _GEN_2136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2138 = 9'hf8 == r_count_6_io_out ? io_r_248_b : _GEN_2137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2139 = 9'hf9 == r_count_6_io_out ? io_r_249_b : _GEN_2138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2140 = 9'hfa == r_count_6_io_out ? io_r_250_b : _GEN_2139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2141 = 9'hfb == r_count_6_io_out ? io_r_251_b : _GEN_2140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2142 = 9'hfc == r_count_6_io_out ? io_r_252_b : _GEN_2141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2143 = 9'hfd == r_count_6_io_out ? io_r_253_b : _GEN_2142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2144 = 9'hfe == r_count_6_io_out ? io_r_254_b : _GEN_2143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2145 = 9'hff == r_count_6_io_out ? io_r_255_b : _GEN_2144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2146 = 9'h100 == r_count_6_io_out ? io_r_256_b : _GEN_2145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2147 = 9'h101 == r_count_6_io_out ? io_r_257_b : _GEN_2146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2148 = 9'h102 == r_count_6_io_out ? io_r_258_b : _GEN_2147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2149 = 9'h103 == r_count_6_io_out ? io_r_259_b : _GEN_2148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2150 = 9'h104 == r_count_6_io_out ? io_r_260_b : _GEN_2149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2151 = 9'h105 == r_count_6_io_out ? io_r_261_b : _GEN_2150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2152 = 9'h106 == r_count_6_io_out ? io_r_262_b : _GEN_2151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2153 = 9'h107 == r_count_6_io_out ? io_r_263_b : _GEN_2152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2154 = 9'h108 == r_count_6_io_out ? io_r_264_b : _GEN_2153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2155 = 9'h109 == r_count_6_io_out ? io_r_265_b : _GEN_2154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2156 = 9'h10a == r_count_6_io_out ? io_r_266_b : _GEN_2155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2157 = 9'h10b == r_count_6_io_out ? io_r_267_b : _GEN_2156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2158 = 9'h10c == r_count_6_io_out ? io_r_268_b : _GEN_2157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2159 = 9'h10d == r_count_6_io_out ? io_r_269_b : _GEN_2158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2160 = 9'h10e == r_count_6_io_out ? io_r_270_b : _GEN_2159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2161 = 9'h10f == r_count_6_io_out ? io_r_271_b : _GEN_2160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2162 = 9'h110 == r_count_6_io_out ? io_r_272_b : _GEN_2161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2163 = 9'h111 == r_count_6_io_out ? io_r_273_b : _GEN_2162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2164 = 9'h112 == r_count_6_io_out ? io_r_274_b : _GEN_2163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2165 = 9'h113 == r_count_6_io_out ? io_r_275_b : _GEN_2164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2166 = 9'h114 == r_count_6_io_out ? io_r_276_b : _GEN_2165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2167 = 9'h115 == r_count_6_io_out ? io_r_277_b : _GEN_2166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2168 = 9'h116 == r_count_6_io_out ? io_r_278_b : _GEN_2167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2169 = 9'h117 == r_count_6_io_out ? io_r_279_b : _GEN_2168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2170 = 9'h118 == r_count_6_io_out ? io_r_280_b : _GEN_2169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2171 = 9'h119 == r_count_6_io_out ? io_r_281_b : _GEN_2170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2172 = 9'h11a == r_count_6_io_out ? io_r_282_b : _GEN_2171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2173 = 9'h11b == r_count_6_io_out ? io_r_283_b : _GEN_2172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2174 = 9'h11c == r_count_6_io_out ? io_r_284_b : _GEN_2173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2175 = 9'h11d == r_count_6_io_out ? io_r_285_b : _GEN_2174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2176 = 9'h11e == r_count_6_io_out ? io_r_286_b : _GEN_2175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2177 = 9'h11f == r_count_6_io_out ? io_r_287_b : _GEN_2176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2178 = 9'h120 == r_count_6_io_out ? io_r_288_b : _GEN_2177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2179 = 9'h121 == r_count_6_io_out ? io_r_289_b : _GEN_2178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2180 = 9'h122 == r_count_6_io_out ? io_r_290_b : _GEN_2179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2181 = 9'h123 == r_count_6_io_out ? io_r_291_b : _GEN_2180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2182 = 9'h124 == r_count_6_io_out ? io_r_292_b : _GEN_2181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2183 = 9'h125 == r_count_6_io_out ? io_r_293_b : _GEN_2182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2184 = 9'h126 == r_count_6_io_out ? io_r_294_b : _GEN_2183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2185 = 9'h127 == r_count_6_io_out ? io_r_295_b : _GEN_2184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2186 = 9'h128 == r_count_6_io_out ? io_r_296_b : _GEN_2185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2187 = 9'h129 == r_count_6_io_out ? io_r_297_b : _GEN_2186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2188 = 9'h12a == r_count_6_io_out ? io_r_298_b : _GEN_2187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2191 = 9'h1 == r_count_7_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2192 = 9'h2 == r_count_7_io_out ? io_r_2_b : _GEN_2191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2193 = 9'h3 == r_count_7_io_out ? io_r_3_b : _GEN_2192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2194 = 9'h4 == r_count_7_io_out ? io_r_4_b : _GEN_2193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2195 = 9'h5 == r_count_7_io_out ? io_r_5_b : _GEN_2194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2196 = 9'h6 == r_count_7_io_out ? io_r_6_b : _GEN_2195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2197 = 9'h7 == r_count_7_io_out ? io_r_7_b : _GEN_2196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2198 = 9'h8 == r_count_7_io_out ? io_r_8_b : _GEN_2197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2199 = 9'h9 == r_count_7_io_out ? io_r_9_b : _GEN_2198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2200 = 9'ha == r_count_7_io_out ? io_r_10_b : _GEN_2199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2201 = 9'hb == r_count_7_io_out ? io_r_11_b : _GEN_2200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2202 = 9'hc == r_count_7_io_out ? io_r_12_b : _GEN_2201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2203 = 9'hd == r_count_7_io_out ? io_r_13_b : _GEN_2202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2204 = 9'he == r_count_7_io_out ? io_r_14_b : _GEN_2203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2205 = 9'hf == r_count_7_io_out ? io_r_15_b : _GEN_2204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2206 = 9'h10 == r_count_7_io_out ? io_r_16_b : _GEN_2205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2207 = 9'h11 == r_count_7_io_out ? io_r_17_b : _GEN_2206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2208 = 9'h12 == r_count_7_io_out ? io_r_18_b : _GEN_2207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2209 = 9'h13 == r_count_7_io_out ? io_r_19_b : _GEN_2208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2210 = 9'h14 == r_count_7_io_out ? io_r_20_b : _GEN_2209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2211 = 9'h15 == r_count_7_io_out ? io_r_21_b : _GEN_2210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2212 = 9'h16 == r_count_7_io_out ? io_r_22_b : _GEN_2211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2213 = 9'h17 == r_count_7_io_out ? io_r_23_b : _GEN_2212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2214 = 9'h18 == r_count_7_io_out ? io_r_24_b : _GEN_2213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2215 = 9'h19 == r_count_7_io_out ? io_r_25_b : _GEN_2214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2216 = 9'h1a == r_count_7_io_out ? io_r_26_b : _GEN_2215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2217 = 9'h1b == r_count_7_io_out ? io_r_27_b : _GEN_2216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2218 = 9'h1c == r_count_7_io_out ? io_r_28_b : _GEN_2217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2219 = 9'h1d == r_count_7_io_out ? io_r_29_b : _GEN_2218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2220 = 9'h1e == r_count_7_io_out ? io_r_30_b : _GEN_2219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2221 = 9'h1f == r_count_7_io_out ? io_r_31_b : _GEN_2220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2222 = 9'h20 == r_count_7_io_out ? io_r_32_b : _GEN_2221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2223 = 9'h21 == r_count_7_io_out ? io_r_33_b : _GEN_2222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2224 = 9'h22 == r_count_7_io_out ? io_r_34_b : _GEN_2223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2225 = 9'h23 == r_count_7_io_out ? io_r_35_b : _GEN_2224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2226 = 9'h24 == r_count_7_io_out ? io_r_36_b : _GEN_2225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2227 = 9'h25 == r_count_7_io_out ? io_r_37_b : _GEN_2226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2228 = 9'h26 == r_count_7_io_out ? io_r_38_b : _GEN_2227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2229 = 9'h27 == r_count_7_io_out ? io_r_39_b : _GEN_2228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2230 = 9'h28 == r_count_7_io_out ? io_r_40_b : _GEN_2229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2231 = 9'h29 == r_count_7_io_out ? io_r_41_b : _GEN_2230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2232 = 9'h2a == r_count_7_io_out ? io_r_42_b : _GEN_2231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2233 = 9'h2b == r_count_7_io_out ? io_r_43_b : _GEN_2232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2234 = 9'h2c == r_count_7_io_out ? io_r_44_b : _GEN_2233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2235 = 9'h2d == r_count_7_io_out ? io_r_45_b : _GEN_2234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2236 = 9'h2e == r_count_7_io_out ? io_r_46_b : _GEN_2235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2237 = 9'h2f == r_count_7_io_out ? io_r_47_b : _GEN_2236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2238 = 9'h30 == r_count_7_io_out ? io_r_48_b : _GEN_2237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2239 = 9'h31 == r_count_7_io_out ? io_r_49_b : _GEN_2238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2240 = 9'h32 == r_count_7_io_out ? io_r_50_b : _GEN_2239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2241 = 9'h33 == r_count_7_io_out ? io_r_51_b : _GEN_2240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2242 = 9'h34 == r_count_7_io_out ? io_r_52_b : _GEN_2241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2243 = 9'h35 == r_count_7_io_out ? io_r_53_b : _GEN_2242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2244 = 9'h36 == r_count_7_io_out ? io_r_54_b : _GEN_2243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2245 = 9'h37 == r_count_7_io_out ? io_r_55_b : _GEN_2244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2246 = 9'h38 == r_count_7_io_out ? io_r_56_b : _GEN_2245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2247 = 9'h39 == r_count_7_io_out ? io_r_57_b : _GEN_2246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2248 = 9'h3a == r_count_7_io_out ? io_r_58_b : _GEN_2247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2249 = 9'h3b == r_count_7_io_out ? io_r_59_b : _GEN_2248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2250 = 9'h3c == r_count_7_io_out ? io_r_60_b : _GEN_2249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2251 = 9'h3d == r_count_7_io_out ? io_r_61_b : _GEN_2250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2252 = 9'h3e == r_count_7_io_out ? io_r_62_b : _GEN_2251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2253 = 9'h3f == r_count_7_io_out ? io_r_63_b : _GEN_2252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2254 = 9'h40 == r_count_7_io_out ? io_r_64_b : _GEN_2253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2255 = 9'h41 == r_count_7_io_out ? io_r_65_b : _GEN_2254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2256 = 9'h42 == r_count_7_io_out ? io_r_66_b : _GEN_2255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2257 = 9'h43 == r_count_7_io_out ? io_r_67_b : _GEN_2256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2258 = 9'h44 == r_count_7_io_out ? io_r_68_b : _GEN_2257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2259 = 9'h45 == r_count_7_io_out ? io_r_69_b : _GEN_2258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2260 = 9'h46 == r_count_7_io_out ? io_r_70_b : _GEN_2259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2261 = 9'h47 == r_count_7_io_out ? io_r_71_b : _GEN_2260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2262 = 9'h48 == r_count_7_io_out ? io_r_72_b : _GEN_2261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2263 = 9'h49 == r_count_7_io_out ? io_r_73_b : _GEN_2262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2264 = 9'h4a == r_count_7_io_out ? io_r_74_b : _GEN_2263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2265 = 9'h4b == r_count_7_io_out ? io_r_75_b : _GEN_2264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2266 = 9'h4c == r_count_7_io_out ? io_r_76_b : _GEN_2265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2267 = 9'h4d == r_count_7_io_out ? io_r_77_b : _GEN_2266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2268 = 9'h4e == r_count_7_io_out ? io_r_78_b : _GEN_2267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2269 = 9'h4f == r_count_7_io_out ? io_r_79_b : _GEN_2268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2270 = 9'h50 == r_count_7_io_out ? io_r_80_b : _GEN_2269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2271 = 9'h51 == r_count_7_io_out ? io_r_81_b : _GEN_2270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2272 = 9'h52 == r_count_7_io_out ? io_r_82_b : _GEN_2271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2273 = 9'h53 == r_count_7_io_out ? io_r_83_b : _GEN_2272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2274 = 9'h54 == r_count_7_io_out ? io_r_84_b : _GEN_2273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2275 = 9'h55 == r_count_7_io_out ? io_r_85_b : _GEN_2274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2276 = 9'h56 == r_count_7_io_out ? io_r_86_b : _GEN_2275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2277 = 9'h57 == r_count_7_io_out ? io_r_87_b : _GEN_2276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2278 = 9'h58 == r_count_7_io_out ? io_r_88_b : _GEN_2277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2279 = 9'h59 == r_count_7_io_out ? io_r_89_b : _GEN_2278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2280 = 9'h5a == r_count_7_io_out ? io_r_90_b : _GEN_2279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2281 = 9'h5b == r_count_7_io_out ? io_r_91_b : _GEN_2280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2282 = 9'h5c == r_count_7_io_out ? io_r_92_b : _GEN_2281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2283 = 9'h5d == r_count_7_io_out ? io_r_93_b : _GEN_2282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2284 = 9'h5e == r_count_7_io_out ? io_r_94_b : _GEN_2283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2285 = 9'h5f == r_count_7_io_out ? io_r_95_b : _GEN_2284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2286 = 9'h60 == r_count_7_io_out ? io_r_96_b : _GEN_2285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2287 = 9'h61 == r_count_7_io_out ? io_r_97_b : _GEN_2286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2288 = 9'h62 == r_count_7_io_out ? io_r_98_b : _GEN_2287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2289 = 9'h63 == r_count_7_io_out ? io_r_99_b : _GEN_2288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2290 = 9'h64 == r_count_7_io_out ? io_r_100_b : _GEN_2289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2291 = 9'h65 == r_count_7_io_out ? io_r_101_b : _GEN_2290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2292 = 9'h66 == r_count_7_io_out ? io_r_102_b : _GEN_2291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2293 = 9'h67 == r_count_7_io_out ? io_r_103_b : _GEN_2292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2294 = 9'h68 == r_count_7_io_out ? io_r_104_b : _GEN_2293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2295 = 9'h69 == r_count_7_io_out ? io_r_105_b : _GEN_2294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2296 = 9'h6a == r_count_7_io_out ? io_r_106_b : _GEN_2295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2297 = 9'h6b == r_count_7_io_out ? io_r_107_b : _GEN_2296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2298 = 9'h6c == r_count_7_io_out ? io_r_108_b : _GEN_2297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2299 = 9'h6d == r_count_7_io_out ? io_r_109_b : _GEN_2298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2300 = 9'h6e == r_count_7_io_out ? io_r_110_b : _GEN_2299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2301 = 9'h6f == r_count_7_io_out ? io_r_111_b : _GEN_2300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2302 = 9'h70 == r_count_7_io_out ? io_r_112_b : _GEN_2301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2303 = 9'h71 == r_count_7_io_out ? io_r_113_b : _GEN_2302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2304 = 9'h72 == r_count_7_io_out ? io_r_114_b : _GEN_2303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2305 = 9'h73 == r_count_7_io_out ? io_r_115_b : _GEN_2304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2306 = 9'h74 == r_count_7_io_out ? io_r_116_b : _GEN_2305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2307 = 9'h75 == r_count_7_io_out ? io_r_117_b : _GEN_2306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2308 = 9'h76 == r_count_7_io_out ? io_r_118_b : _GEN_2307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2309 = 9'h77 == r_count_7_io_out ? io_r_119_b : _GEN_2308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2310 = 9'h78 == r_count_7_io_out ? io_r_120_b : _GEN_2309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2311 = 9'h79 == r_count_7_io_out ? io_r_121_b : _GEN_2310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2312 = 9'h7a == r_count_7_io_out ? io_r_122_b : _GEN_2311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2313 = 9'h7b == r_count_7_io_out ? io_r_123_b : _GEN_2312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2314 = 9'h7c == r_count_7_io_out ? io_r_124_b : _GEN_2313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2315 = 9'h7d == r_count_7_io_out ? io_r_125_b : _GEN_2314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2316 = 9'h7e == r_count_7_io_out ? io_r_126_b : _GEN_2315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2317 = 9'h7f == r_count_7_io_out ? io_r_127_b : _GEN_2316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2318 = 9'h80 == r_count_7_io_out ? io_r_128_b : _GEN_2317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2319 = 9'h81 == r_count_7_io_out ? io_r_129_b : _GEN_2318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2320 = 9'h82 == r_count_7_io_out ? io_r_130_b : _GEN_2319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2321 = 9'h83 == r_count_7_io_out ? io_r_131_b : _GEN_2320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2322 = 9'h84 == r_count_7_io_out ? io_r_132_b : _GEN_2321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2323 = 9'h85 == r_count_7_io_out ? io_r_133_b : _GEN_2322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2324 = 9'h86 == r_count_7_io_out ? io_r_134_b : _GEN_2323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2325 = 9'h87 == r_count_7_io_out ? io_r_135_b : _GEN_2324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2326 = 9'h88 == r_count_7_io_out ? io_r_136_b : _GEN_2325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2327 = 9'h89 == r_count_7_io_out ? io_r_137_b : _GEN_2326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2328 = 9'h8a == r_count_7_io_out ? io_r_138_b : _GEN_2327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2329 = 9'h8b == r_count_7_io_out ? io_r_139_b : _GEN_2328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2330 = 9'h8c == r_count_7_io_out ? io_r_140_b : _GEN_2329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2331 = 9'h8d == r_count_7_io_out ? io_r_141_b : _GEN_2330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2332 = 9'h8e == r_count_7_io_out ? io_r_142_b : _GEN_2331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2333 = 9'h8f == r_count_7_io_out ? io_r_143_b : _GEN_2332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2334 = 9'h90 == r_count_7_io_out ? io_r_144_b : _GEN_2333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2335 = 9'h91 == r_count_7_io_out ? io_r_145_b : _GEN_2334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2336 = 9'h92 == r_count_7_io_out ? io_r_146_b : _GEN_2335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2337 = 9'h93 == r_count_7_io_out ? io_r_147_b : _GEN_2336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2338 = 9'h94 == r_count_7_io_out ? io_r_148_b : _GEN_2337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2339 = 9'h95 == r_count_7_io_out ? io_r_149_b : _GEN_2338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2340 = 9'h96 == r_count_7_io_out ? io_r_150_b : _GEN_2339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2341 = 9'h97 == r_count_7_io_out ? io_r_151_b : _GEN_2340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2342 = 9'h98 == r_count_7_io_out ? io_r_152_b : _GEN_2341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2343 = 9'h99 == r_count_7_io_out ? io_r_153_b : _GEN_2342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2344 = 9'h9a == r_count_7_io_out ? io_r_154_b : _GEN_2343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2345 = 9'h9b == r_count_7_io_out ? io_r_155_b : _GEN_2344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2346 = 9'h9c == r_count_7_io_out ? io_r_156_b : _GEN_2345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2347 = 9'h9d == r_count_7_io_out ? io_r_157_b : _GEN_2346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2348 = 9'h9e == r_count_7_io_out ? io_r_158_b : _GEN_2347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2349 = 9'h9f == r_count_7_io_out ? io_r_159_b : _GEN_2348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2350 = 9'ha0 == r_count_7_io_out ? io_r_160_b : _GEN_2349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2351 = 9'ha1 == r_count_7_io_out ? io_r_161_b : _GEN_2350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2352 = 9'ha2 == r_count_7_io_out ? io_r_162_b : _GEN_2351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2353 = 9'ha3 == r_count_7_io_out ? io_r_163_b : _GEN_2352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2354 = 9'ha4 == r_count_7_io_out ? io_r_164_b : _GEN_2353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2355 = 9'ha5 == r_count_7_io_out ? io_r_165_b : _GEN_2354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2356 = 9'ha6 == r_count_7_io_out ? io_r_166_b : _GEN_2355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2357 = 9'ha7 == r_count_7_io_out ? io_r_167_b : _GEN_2356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2358 = 9'ha8 == r_count_7_io_out ? io_r_168_b : _GEN_2357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2359 = 9'ha9 == r_count_7_io_out ? io_r_169_b : _GEN_2358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2360 = 9'haa == r_count_7_io_out ? io_r_170_b : _GEN_2359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2361 = 9'hab == r_count_7_io_out ? io_r_171_b : _GEN_2360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2362 = 9'hac == r_count_7_io_out ? io_r_172_b : _GEN_2361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2363 = 9'had == r_count_7_io_out ? io_r_173_b : _GEN_2362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2364 = 9'hae == r_count_7_io_out ? io_r_174_b : _GEN_2363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2365 = 9'haf == r_count_7_io_out ? io_r_175_b : _GEN_2364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2366 = 9'hb0 == r_count_7_io_out ? io_r_176_b : _GEN_2365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2367 = 9'hb1 == r_count_7_io_out ? io_r_177_b : _GEN_2366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2368 = 9'hb2 == r_count_7_io_out ? io_r_178_b : _GEN_2367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2369 = 9'hb3 == r_count_7_io_out ? io_r_179_b : _GEN_2368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2370 = 9'hb4 == r_count_7_io_out ? io_r_180_b : _GEN_2369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2371 = 9'hb5 == r_count_7_io_out ? io_r_181_b : _GEN_2370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2372 = 9'hb6 == r_count_7_io_out ? io_r_182_b : _GEN_2371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2373 = 9'hb7 == r_count_7_io_out ? io_r_183_b : _GEN_2372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2374 = 9'hb8 == r_count_7_io_out ? io_r_184_b : _GEN_2373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2375 = 9'hb9 == r_count_7_io_out ? io_r_185_b : _GEN_2374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2376 = 9'hba == r_count_7_io_out ? io_r_186_b : _GEN_2375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2377 = 9'hbb == r_count_7_io_out ? io_r_187_b : _GEN_2376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2378 = 9'hbc == r_count_7_io_out ? io_r_188_b : _GEN_2377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2379 = 9'hbd == r_count_7_io_out ? io_r_189_b : _GEN_2378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2380 = 9'hbe == r_count_7_io_out ? io_r_190_b : _GEN_2379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2381 = 9'hbf == r_count_7_io_out ? io_r_191_b : _GEN_2380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2382 = 9'hc0 == r_count_7_io_out ? io_r_192_b : _GEN_2381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2383 = 9'hc1 == r_count_7_io_out ? io_r_193_b : _GEN_2382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2384 = 9'hc2 == r_count_7_io_out ? io_r_194_b : _GEN_2383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2385 = 9'hc3 == r_count_7_io_out ? io_r_195_b : _GEN_2384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2386 = 9'hc4 == r_count_7_io_out ? io_r_196_b : _GEN_2385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2387 = 9'hc5 == r_count_7_io_out ? io_r_197_b : _GEN_2386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2388 = 9'hc6 == r_count_7_io_out ? io_r_198_b : _GEN_2387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2389 = 9'hc7 == r_count_7_io_out ? io_r_199_b : _GEN_2388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2390 = 9'hc8 == r_count_7_io_out ? io_r_200_b : _GEN_2389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2391 = 9'hc9 == r_count_7_io_out ? io_r_201_b : _GEN_2390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2392 = 9'hca == r_count_7_io_out ? io_r_202_b : _GEN_2391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2393 = 9'hcb == r_count_7_io_out ? io_r_203_b : _GEN_2392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2394 = 9'hcc == r_count_7_io_out ? io_r_204_b : _GEN_2393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2395 = 9'hcd == r_count_7_io_out ? io_r_205_b : _GEN_2394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2396 = 9'hce == r_count_7_io_out ? io_r_206_b : _GEN_2395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2397 = 9'hcf == r_count_7_io_out ? io_r_207_b : _GEN_2396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2398 = 9'hd0 == r_count_7_io_out ? io_r_208_b : _GEN_2397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2399 = 9'hd1 == r_count_7_io_out ? io_r_209_b : _GEN_2398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2400 = 9'hd2 == r_count_7_io_out ? io_r_210_b : _GEN_2399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2401 = 9'hd3 == r_count_7_io_out ? io_r_211_b : _GEN_2400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2402 = 9'hd4 == r_count_7_io_out ? io_r_212_b : _GEN_2401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2403 = 9'hd5 == r_count_7_io_out ? io_r_213_b : _GEN_2402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2404 = 9'hd6 == r_count_7_io_out ? io_r_214_b : _GEN_2403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2405 = 9'hd7 == r_count_7_io_out ? io_r_215_b : _GEN_2404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2406 = 9'hd8 == r_count_7_io_out ? io_r_216_b : _GEN_2405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2407 = 9'hd9 == r_count_7_io_out ? io_r_217_b : _GEN_2406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2408 = 9'hda == r_count_7_io_out ? io_r_218_b : _GEN_2407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2409 = 9'hdb == r_count_7_io_out ? io_r_219_b : _GEN_2408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2410 = 9'hdc == r_count_7_io_out ? io_r_220_b : _GEN_2409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2411 = 9'hdd == r_count_7_io_out ? io_r_221_b : _GEN_2410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2412 = 9'hde == r_count_7_io_out ? io_r_222_b : _GEN_2411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2413 = 9'hdf == r_count_7_io_out ? io_r_223_b : _GEN_2412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2414 = 9'he0 == r_count_7_io_out ? io_r_224_b : _GEN_2413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2415 = 9'he1 == r_count_7_io_out ? io_r_225_b : _GEN_2414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2416 = 9'he2 == r_count_7_io_out ? io_r_226_b : _GEN_2415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2417 = 9'he3 == r_count_7_io_out ? io_r_227_b : _GEN_2416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2418 = 9'he4 == r_count_7_io_out ? io_r_228_b : _GEN_2417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2419 = 9'he5 == r_count_7_io_out ? io_r_229_b : _GEN_2418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2420 = 9'he6 == r_count_7_io_out ? io_r_230_b : _GEN_2419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2421 = 9'he7 == r_count_7_io_out ? io_r_231_b : _GEN_2420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2422 = 9'he8 == r_count_7_io_out ? io_r_232_b : _GEN_2421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2423 = 9'he9 == r_count_7_io_out ? io_r_233_b : _GEN_2422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2424 = 9'hea == r_count_7_io_out ? io_r_234_b : _GEN_2423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2425 = 9'heb == r_count_7_io_out ? io_r_235_b : _GEN_2424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2426 = 9'hec == r_count_7_io_out ? io_r_236_b : _GEN_2425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2427 = 9'hed == r_count_7_io_out ? io_r_237_b : _GEN_2426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2428 = 9'hee == r_count_7_io_out ? io_r_238_b : _GEN_2427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2429 = 9'hef == r_count_7_io_out ? io_r_239_b : _GEN_2428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2430 = 9'hf0 == r_count_7_io_out ? io_r_240_b : _GEN_2429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2431 = 9'hf1 == r_count_7_io_out ? io_r_241_b : _GEN_2430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2432 = 9'hf2 == r_count_7_io_out ? io_r_242_b : _GEN_2431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2433 = 9'hf3 == r_count_7_io_out ? io_r_243_b : _GEN_2432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2434 = 9'hf4 == r_count_7_io_out ? io_r_244_b : _GEN_2433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2435 = 9'hf5 == r_count_7_io_out ? io_r_245_b : _GEN_2434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2436 = 9'hf6 == r_count_7_io_out ? io_r_246_b : _GEN_2435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2437 = 9'hf7 == r_count_7_io_out ? io_r_247_b : _GEN_2436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2438 = 9'hf8 == r_count_7_io_out ? io_r_248_b : _GEN_2437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2439 = 9'hf9 == r_count_7_io_out ? io_r_249_b : _GEN_2438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2440 = 9'hfa == r_count_7_io_out ? io_r_250_b : _GEN_2439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2441 = 9'hfb == r_count_7_io_out ? io_r_251_b : _GEN_2440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2442 = 9'hfc == r_count_7_io_out ? io_r_252_b : _GEN_2441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2443 = 9'hfd == r_count_7_io_out ? io_r_253_b : _GEN_2442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2444 = 9'hfe == r_count_7_io_out ? io_r_254_b : _GEN_2443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2445 = 9'hff == r_count_7_io_out ? io_r_255_b : _GEN_2444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2446 = 9'h100 == r_count_7_io_out ? io_r_256_b : _GEN_2445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2447 = 9'h101 == r_count_7_io_out ? io_r_257_b : _GEN_2446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2448 = 9'h102 == r_count_7_io_out ? io_r_258_b : _GEN_2447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2449 = 9'h103 == r_count_7_io_out ? io_r_259_b : _GEN_2448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2450 = 9'h104 == r_count_7_io_out ? io_r_260_b : _GEN_2449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2451 = 9'h105 == r_count_7_io_out ? io_r_261_b : _GEN_2450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2452 = 9'h106 == r_count_7_io_out ? io_r_262_b : _GEN_2451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2453 = 9'h107 == r_count_7_io_out ? io_r_263_b : _GEN_2452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2454 = 9'h108 == r_count_7_io_out ? io_r_264_b : _GEN_2453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2455 = 9'h109 == r_count_7_io_out ? io_r_265_b : _GEN_2454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2456 = 9'h10a == r_count_7_io_out ? io_r_266_b : _GEN_2455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2457 = 9'h10b == r_count_7_io_out ? io_r_267_b : _GEN_2456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2458 = 9'h10c == r_count_7_io_out ? io_r_268_b : _GEN_2457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2459 = 9'h10d == r_count_7_io_out ? io_r_269_b : _GEN_2458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2460 = 9'h10e == r_count_7_io_out ? io_r_270_b : _GEN_2459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2461 = 9'h10f == r_count_7_io_out ? io_r_271_b : _GEN_2460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2462 = 9'h110 == r_count_7_io_out ? io_r_272_b : _GEN_2461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2463 = 9'h111 == r_count_7_io_out ? io_r_273_b : _GEN_2462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2464 = 9'h112 == r_count_7_io_out ? io_r_274_b : _GEN_2463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2465 = 9'h113 == r_count_7_io_out ? io_r_275_b : _GEN_2464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2466 = 9'h114 == r_count_7_io_out ? io_r_276_b : _GEN_2465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2467 = 9'h115 == r_count_7_io_out ? io_r_277_b : _GEN_2466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2468 = 9'h116 == r_count_7_io_out ? io_r_278_b : _GEN_2467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2469 = 9'h117 == r_count_7_io_out ? io_r_279_b : _GEN_2468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2470 = 9'h118 == r_count_7_io_out ? io_r_280_b : _GEN_2469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2471 = 9'h119 == r_count_7_io_out ? io_r_281_b : _GEN_2470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2472 = 9'h11a == r_count_7_io_out ? io_r_282_b : _GEN_2471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2473 = 9'h11b == r_count_7_io_out ? io_r_283_b : _GEN_2472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2474 = 9'h11c == r_count_7_io_out ? io_r_284_b : _GEN_2473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2475 = 9'h11d == r_count_7_io_out ? io_r_285_b : _GEN_2474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2476 = 9'h11e == r_count_7_io_out ? io_r_286_b : _GEN_2475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2477 = 9'h11f == r_count_7_io_out ? io_r_287_b : _GEN_2476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2478 = 9'h120 == r_count_7_io_out ? io_r_288_b : _GEN_2477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2479 = 9'h121 == r_count_7_io_out ? io_r_289_b : _GEN_2478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2480 = 9'h122 == r_count_7_io_out ? io_r_290_b : _GEN_2479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2481 = 9'h123 == r_count_7_io_out ? io_r_291_b : _GEN_2480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2482 = 9'h124 == r_count_7_io_out ? io_r_292_b : _GEN_2481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2483 = 9'h125 == r_count_7_io_out ? io_r_293_b : _GEN_2482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2484 = 9'h126 == r_count_7_io_out ? io_r_294_b : _GEN_2483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2485 = 9'h127 == r_count_7_io_out ? io_r_295_b : _GEN_2484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2486 = 9'h128 == r_count_7_io_out ? io_r_296_b : _GEN_2485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2487 = 9'h129 == r_count_7_io_out ? io_r_297_b : _GEN_2486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2488 = 9'h12a == r_count_7_io_out ? io_r_298_b : _GEN_2487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2491 = 9'h1 == r_count_8_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2492 = 9'h2 == r_count_8_io_out ? io_r_2_b : _GEN_2491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2493 = 9'h3 == r_count_8_io_out ? io_r_3_b : _GEN_2492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2494 = 9'h4 == r_count_8_io_out ? io_r_4_b : _GEN_2493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2495 = 9'h5 == r_count_8_io_out ? io_r_5_b : _GEN_2494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2496 = 9'h6 == r_count_8_io_out ? io_r_6_b : _GEN_2495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2497 = 9'h7 == r_count_8_io_out ? io_r_7_b : _GEN_2496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2498 = 9'h8 == r_count_8_io_out ? io_r_8_b : _GEN_2497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2499 = 9'h9 == r_count_8_io_out ? io_r_9_b : _GEN_2498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2500 = 9'ha == r_count_8_io_out ? io_r_10_b : _GEN_2499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2501 = 9'hb == r_count_8_io_out ? io_r_11_b : _GEN_2500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2502 = 9'hc == r_count_8_io_out ? io_r_12_b : _GEN_2501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2503 = 9'hd == r_count_8_io_out ? io_r_13_b : _GEN_2502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2504 = 9'he == r_count_8_io_out ? io_r_14_b : _GEN_2503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2505 = 9'hf == r_count_8_io_out ? io_r_15_b : _GEN_2504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2506 = 9'h10 == r_count_8_io_out ? io_r_16_b : _GEN_2505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2507 = 9'h11 == r_count_8_io_out ? io_r_17_b : _GEN_2506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2508 = 9'h12 == r_count_8_io_out ? io_r_18_b : _GEN_2507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2509 = 9'h13 == r_count_8_io_out ? io_r_19_b : _GEN_2508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2510 = 9'h14 == r_count_8_io_out ? io_r_20_b : _GEN_2509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2511 = 9'h15 == r_count_8_io_out ? io_r_21_b : _GEN_2510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2512 = 9'h16 == r_count_8_io_out ? io_r_22_b : _GEN_2511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2513 = 9'h17 == r_count_8_io_out ? io_r_23_b : _GEN_2512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2514 = 9'h18 == r_count_8_io_out ? io_r_24_b : _GEN_2513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2515 = 9'h19 == r_count_8_io_out ? io_r_25_b : _GEN_2514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2516 = 9'h1a == r_count_8_io_out ? io_r_26_b : _GEN_2515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2517 = 9'h1b == r_count_8_io_out ? io_r_27_b : _GEN_2516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2518 = 9'h1c == r_count_8_io_out ? io_r_28_b : _GEN_2517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2519 = 9'h1d == r_count_8_io_out ? io_r_29_b : _GEN_2518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2520 = 9'h1e == r_count_8_io_out ? io_r_30_b : _GEN_2519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2521 = 9'h1f == r_count_8_io_out ? io_r_31_b : _GEN_2520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2522 = 9'h20 == r_count_8_io_out ? io_r_32_b : _GEN_2521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2523 = 9'h21 == r_count_8_io_out ? io_r_33_b : _GEN_2522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2524 = 9'h22 == r_count_8_io_out ? io_r_34_b : _GEN_2523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2525 = 9'h23 == r_count_8_io_out ? io_r_35_b : _GEN_2524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2526 = 9'h24 == r_count_8_io_out ? io_r_36_b : _GEN_2525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2527 = 9'h25 == r_count_8_io_out ? io_r_37_b : _GEN_2526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2528 = 9'h26 == r_count_8_io_out ? io_r_38_b : _GEN_2527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2529 = 9'h27 == r_count_8_io_out ? io_r_39_b : _GEN_2528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2530 = 9'h28 == r_count_8_io_out ? io_r_40_b : _GEN_2529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2531 = 9'h29 == r_count_8_io_out ? io_r_41_b : _GEN_2530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2532 = 9'h2a == r_count_8_io_out ? io_r_42_b : _GEN_2531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2533 = 9'h2b == r_count_8_io_out ? io_r_43_b : _GEN_2532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2534 = 9'h2c == r_count_8_io_out ? io_r_44_b : _GEN_2533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2535 = 9'h2d == r_count_8_io_out ? io_r_45_b : _GEN_2534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2536 = 9'h2e == r_count_8_io_out ? io_r_46_b : _GEN_2535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2537 = 9'h2f == r_count_8_io_out ? io_r_47_b : _GEN_2536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2538 = 9'h30 == r_count_8_io_out ? io_r_48_b : _GEN_2537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2539 = 9'h31 == r_count_8_io_out ? io_r_49_b : _GEN_2538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2540 = 9'h32 == r_count_8_io_out ? io_r_50_b : _GEN_2539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2541 = 9'h33 == r_count_8_io_out ? io_r_51_b : _GEN_2540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2542 = 9'h34 == r_count_8_io_out ? io_r_52_b : _GEN_2541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2543 = 9'h35 == r_count_8_io_out ? io_r_53_b : _GEN_2542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2544 = 9'h36 == r_count_8_io_out ? io_r_54_b : _GEN_2543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2545 = 9'h37 == r_count_8_io_out ? io_r_55_b : _GEN_2544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2546 = 9'h38 == r_count_8_io_out ? io_r_56_b : _GEN_2545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2547 = 9'h39 == r_count_8_io_out ? io_r_57_b : _GEN_2546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2548 = 9'h3a == r_count_8_io_out ? io_r_58_b : _GEN_2547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2549 = 9'h3b == r_count_8_io_out ? io_r_59_b : _GEN_2548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2550 = 9'h3c == r_count_8_io_out ? io_r_60_b : _GEN_2549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2551 = 9'h3d == r_count_8_io_out ? io_r_61_b : _GEN_2550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2552 = 9'h3e == r_count_8_io_out ? io_r_62_b : _GEN_2551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2553 = 9'h3f == r_count_8_io_out ? io_r_63_b : _GEN_2552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2554 = 9'h40 == r_count_8_io_out ? io_r_64_b : _GEN_2553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2555 = 9'h41 == r_count_8_io_out ? io_r_65_b : _GEN_2554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2556 = 9'h42 == r_count_8_io_out ? io_r_66_b : _GEN_2555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2557 = 9'h43 == r_count_8_io_out ? io_r_67_b : _GEN_2556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2558 = 9'h44 == r_count_8_io_out ? io_r_68_b : _GEN_2557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2559 = 9'h45 == r_count_8_io_out ? io_r_69_b : _GEN_2558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2560 = 9'h46 == r_count_8_io_out ? io_r_70_b : _GEN_2559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2561 = 9'h47 == r_count_8_io_out ? io_r_71_b : _GEN_2560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2562 = 9'h48 == r_count_8_io_out ? io_r_72_b : _GEN_2561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2563 = 9'h49 == r_count_8_io_out ? io_r_73_b : _GEN_2562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2564 = 9'h4a == r_count_8_io_out ? io_r_74_b : _GEN_2563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2565 = 9'h4b == r_count_8_io_out ? io_r_75_b : _GEN_2564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2566 = 9'h4c == r_count_8_io_out ? io_r_76_b : _GEN_2565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2567 = 9'h4d == r_count_8_io_out ? io_r_77_b : _GEN_2566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2568 = 9'h4e == r_count_8_io_out ? io_r_78_b : _GEN_2567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2569 = 9'h4f == r_count_8_io_out ? io_r_79_b : _GEN_2568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2570 = 9'h50 == r_count_8_io_out ? io_r_80_b : _GEN_2569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2571 = 9'h51 == r_count_8_io_out ? io_r_81_b : _GEN_2570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2572 = 9'h52 == r_count_8_io_out ? io_r_82_b : _GEN_2571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2573 = 9'h53 == r_count_8_io_out ? io_r_83_b : _GEN_2572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2574 = 9'h54 == r_count_8_io_out ? io_r_84_b : _GEN_2573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2575 = 9'h55 == r_count_8_io_out ? io_r_85_b : _GEN_2574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2576 = 9'h56 == r_count_8_io_out ? io_r_86_b : _GEN_2575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2577 = 9'h57 == r_count_8_io_out ? io_r_87_b : _GEN_2576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2578 = 9'h58 == r_count_8_io_out ? io_r_88_b : _GEN_2577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2579 = 9'h59 == r_count_8_io_out ? io_r_89_b : _GEN_2578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2580 = 9'h5a == r_count_8_io_out ? io_r_90_b : _GEN_2579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2581 = 9'h5b == r_count_8_io_out ? io_r_91_b : _GEN_2580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2582 = 9'h5c == r_count_8_io_out ? io_r_92_b : _GEN_2581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2583 = 9'h5d == r_count_8_io_out ? io_r_93_b : _GEN_2582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2584 = 9'h5e == r_count_8_io_out ? io_r_94_b : _GEN_2583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2585 = 9'h5f == r_count_8_io_out ? io_r_95_b : _GEN_2584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2586 = 9'h60 == r_count_8_io_out ? io_r_96_b : _GEN_2585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2587 = 9'h61 == r_count_8_io_out ? io_r_97_b : _GEN_2586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2588 = 9'h62 == r_count_8_io_out ? io_r_98_b : _GEN_2587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2589 = 9'h63 == r_count_8_io_out ? io_r_99_b : _GEN_2588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2590 = 9'h64 == r_count_8_io_out ? io_r_100_b : _GEN_2589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2591 = 9'h65 == r_count_8_io_out ? io_r_101_b : _GEN_2590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2592 = 9'h66 == r_count_8_io_out ? io_r_102_b : _GEN_2591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2593 = 9'h67 == r_count_8_io_out ? io_r_103_b : _GEN_2592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2594 = 9'h68 == r_count_8_io_out ? io_r_104_b : _GEN_2593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2595 = 9'h69 == r_count_8_io_out ? io_r_105_b : _GEN_2594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2596 = 9'h6a == r_count_8_io_out ? io_r_106_b : _GEN_2595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2597 = 9'h6b == r_count_8_io_out ? io_r_107_b : _GEN_2596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2598 = 9'h6c == r_count_8_io_out ? io_r_108_b : _GEN_2597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2599 = 9'h6d == r_count_8_io_out ? io_r_109_b : _GEN_2598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2600 = 9'h6e == r_count_8_io_out ? io_r_110_b : _GEN_2599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2601 = 9'h6f == r_count_8_io_out ? io_r_111_b : _GEN_2600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2602 = 9'h70 == r_count_8_io_out ? io_r_112_b : _GEN_2601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2603 = 9'h71 == r_count_8_io_out ? io_r_113_b : _GEN_2602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2604 = 9'h72 == r_count_8_io_out ? io_r_114_b : _GEN_2603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2605 = 9'h73 == r_count_8_io_out ? io_r_115_b : _GEN_2604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2606 = 9'h74 == r_count_8_io_out ? io_r_116_b : _GEN_2605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2607 = 9'h75 == r_count_8_io_out ? io_r_117_b : _GEN_2606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2608 = 9'h76 == r_count_8_io_out ? io_r_118_b : _GEN_2607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2609 = 9'h77 == r_count_8_io_out ? io_r_119_b : _GEN_2608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2610 = 9'h78 == r_count_8_io_out ? io_r_120_b : _GEN_2609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2611 = 9'h79 == r_count_8_io_out ? io_r_121_b : _GEN_2610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2612 = 9'h7a == r_count_8_io_out ? io_r_122_b : _GEN_2611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2613 = 9'h7b == r_count_8_io_out ? io_r_123_b : _GEN_2612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2614 = 9'h7c == r_count_8_io_out ? io_r_124_b : _GEN_2613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2615 = 9'h7d == r_count_8_io_out ? io_r_125_b : _GEN_2614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2616 = 9'h7e == r_count_8_io_out ? io_r_126_b : _GEN_2615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2617 = 9'h7f == r_count_8_io_out ? io_r_127_b : _GEN_2616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2618 = 9'h80 == r_count_8_io_out ? io_r_128_b : _GEN_2617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2619 = 9'h81 == r_count_8_io_out ? io_r_129_b : _GEN_2618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2620 = 9'h82 == r_count_8_io_out ? io_r_130_b : _GEN_2619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2621 = 9'h83 == r_count_8_io_out ? io_r_131_b : _GEN_2620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2622 = 9'h84 == r_count_8_io_out ? io_r_132_b : _GEN_2621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2623 = 9'h85 == r_count_8_io_out ? io_r_133_b : _GEN_2622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2624 = 9'h86 == r_count_8_io_out ? io_r_134_b : _GEN_2623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2625 = 9'h87 == r_count_8_io_out ? io_r_135_b : _GEN_2624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2626 = 9'h88 == r_count_8_io_out ? io_r_136_b : _GEN_2625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2627 = 9'h89 == r_count_8_io_out ? io_r_137_b : _GEN_2626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2628 = 9'h8a == r_count_8_io_out ? io_r_138_b : _GEN_2627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2629 = 9'h8b == r_count_8_io_out ? io_r_139_b : _GEN_2628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2630 = 9'h8c == r_count_8_io_out ? io_r_140_b : _GEN_2629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2631 = 9'h8d == r_count_8_io_out ? io_r_141_b : _GEN_2630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2632 = 9'h8e == r_count_8_io_out ? io_r_142_b : _GEN_2631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2633 = 9'h8f == r_count_8_io_out ? io_r_143_b : _GEN_2632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2634 = 9'h90 == r_count_8_io_out ? io_r_144_b : _GEN_2633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2635 = 9'h91 == r_count_8_io_out ? io_r_145_b : _GEN_2634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2636 = 9'h92 == r_count_8_io_out ? io_r_146_b : _GEN_2635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2637 = 9'h93 == r_count_8_io_out ? io_r_147_b : _GEN_2636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2638 = 9'h94 == r_count_8_io_out ? io_r_148_b : _GEN_2637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2639 = 9'h95 == r_count_8_io_out ? io_r_149_b : _GEN_2638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2640 = 9'h96 == r_count_8_io_out ? io_r_150_b : _GEN_2639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2641 = 9'h97 == r_count_8_io_out ? io_r_151_b : _GEN_2640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2642 = 9'h98 == r_count_8_io_out ? io_r_152_b : _GEN_2641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2643 = 9'h99 == r_count_8_io_out ? io_r_153_b : _GEN_2642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2644 = 9'h9a == r_count_8_io_out ? io_r_154_b : _GEN_2643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2645 = 9'h9b == r_count_8_io_out ? io_r_155_b : _GEN_2644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2646 = 9'h9c == r_count_8_io_out ? io_r_156_b : _GEN_2645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2647 = 9'h9d == r_count_8_io_out ? io_r_157_b : _GEN_2646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2648 = 9'h9e == r_count_8_io_out ? io_r_158_b : _GEN_2647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2649 = 9'h9f == r_count_8_io_out ? io_r_159_b : _GEN_2648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2650 = 9'ha0 == r_count_8_io_out ? io_r_160_b : _GEN_2649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2651 = 9'ha1 == r_count_8_io_out ? io_r_161_b : _GEN_2650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2652 = 9'ha2 == r_count_8_io_out ? io_r_162_b : _GEN_2651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2653 = 9'ha3 == r_count_8_io_out ? io_r_163_b : _GEN_2652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2654 = 9'ha4 == r_count_8_io_out ? io_r_164_b : _GEN_2653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2655 = 9'ha5 == r_count_8_io_out ? io_r_165_b : _GEN_2654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2656 = 9'ha6 == r_count_8_io_out ? io_r_166_b : _GEN_2655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2657 = 9'ha7 == r_count_8_io_out ? io_r_167_b : _GEN_2656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2658 = 9'ha8 == r_count_8_io_out ? io_r_168_b : _GEN_2657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2659 = 9'ha9 == r_count_8_io_out ? io_r_169_b : _GEN_2658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2660 = 9'haa == r_count_8_io_out ? io_r_170_b : _GEN_2659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2661 = 9'hab == r_count_8_io_out ? io_r_171_b : _GEN_2660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2662 = 9'hac == r_count_8_io_out ? io_r_172_b : _GEN_2661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2663 = 9'had == r_count_8_io_out ? io_r_173_b : _GEN_2662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2664 = 9'hae == r_count_8_io_out ? io_r_174_b : _GEN_2663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2665 = 9'haf == r_count_8_io_out ? io_r_175_b : _GEN_2664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2666 = 9'hb0 == r_count_8_io_out ? io_r_176_b : _GEN_2665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2667 = 9'hb1 == r_count_8_io_out ? io_r_177_b : _GEN_2666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2668 = 9'hb2 == r_count_8_io_out ? io_r_178_b : _GEN_2667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2669 = 9'hb3 == r_count_8_io_out ? io_r_179_b : _GEN_2668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2670 = 9'hb4 == r_count_8_io_out ? io_r_180_b : _GEN_2669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2671 = 9'hb5 == r_count_8_io_out ? io_r_181_b : _GEN_2670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2672 = 9'hb6 == r_count_8_io_out ? io_r_182_b : _GEN_2671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2673 = 9'hb7 == r_count_8_io_out ? io_r_183_b : _GEN_2672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2674 = 9'hb8 == r_count_8_io_out ? io_r_184_b : _GEN_2673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2675 = 9'hb9 == r_count_8_io_out ? io_r_185_b : _GEN_2674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2676 = 9'hba == r_count_8_io_out ? io_r_186_b : _GEN_2675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2677 = 9'hbb == r_count_8_io_out ? io_r_187_b : _GEN_2676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2678 = 9'hbc == r_count_8_io_out ? io_r_188_b : _GEN_2677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2679 = 9'hbd == r_count_8_io_out ? io_r_189_b : _GEN_2678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2680 = 9'hbe == r_count_8_io_out ? io_r_190_b : _GEN_2679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2681 = 9'hbf == r_count_8_io_out ? io_r_191_b : _GEN_2680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2682 = 9'hc0 == r_count_8_io_out ? io_r_192_b : _GEN_2681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2683 = 9'hc1 == r_count_8_io_out ? io_r_193_b : _GEN_2682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2684 = 9'hc2 == r_count_8_io_out ? io_r_194_b : _GEN_2683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2685 = 9'hc3 == r_count_8_io_out ? io_r_195_b : _GEN_2684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2686 = 9'hc4 == r_count_8_io_out ? io_r_196_b : _GEN_2685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2687 = 9'hc5 == r_count_8_io_out ? io_r_197_b : _GEN_2686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2688 = 9'hc6 == r_count_8_io_out ? io_r_198_b : _GEN_2687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2689 = 9'hc7 == r_count_8_io_out ? io_r_199_b : _GEN_2688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2690 = 9'hc8 == r_count_8_io_out ? io_r_200_b : _GEN_2689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2691 = 9'hc9 == r_count_8_io_out ? io_r_201_b : _GEN_2690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2692 = 9'hca == r_count_8_io_out ? io_r_202_b : _GEN_2691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2693 = 9'hcb == r_count_8_io_out ? io_r_203_b : _GEN_2692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2694 = 9'hcc == r_count_8_io_out ? io_r_204_b : _GEN_2693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2695 = 9'hcd == r_count_8_io_out ? io_r_205_b : _GEN_2694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2696 = 9'hce == r_count_8_io_out ? io_r_206_b : _GEN_2695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2697 = 9'hcf == r_count_8_io_out ? io_r_207_b : _GEN_2696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2698 = 9'hd0 == r_count_8_io_out ? io_r_208_b : _GEN_2697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2699 = 9'hd1 == r_count_8_io_out ? io_r_209_b : _GEN_2698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2700 = 9'hd2 == r_count_8_io_out ? io_r_210_b : _GEN_2699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2701 = 9'hd3 == r_count_8_io_out ? io_r_211_b : _GEN_2700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2702 = 9'hd4 == r_count_8_io_out ? io_r_212_b : _GEN_2701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2703 = 9'hd5 == r_count_8_io_out ? io_r_213_b : _GEN_2702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2704 = 9'hd6 == r_count_8_io_out ? io_r_214_b : _GEN_2703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2705 = 9'hd7 == r_count_8_io_out ? io_r_215_b : _GEN_2704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2706 = 9'hd8 == r_count_8_io_out ? io_r_216_b : _GEN_2705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2707 = 9'hd9 == r_count_8_io_out ? io_r_217_b : _GEN_2706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2708 = 9'hda == r_count_8_io_out ? io_r_218_b : _GEN_2707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2709 = 9'hdb == r_count_8_io_out ? io_r_219_b : _GEN_2708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2710 = 9'hdc == r_count_8_io_out ? io_r_220_b : _GEN_2709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2711 = 9'hdd == r_count_8_io_out ? io_r_221_b : _GEN_2710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2712 = 9'hde == r_count_8_io_out ? io_r_222_b : _GEN_2711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2713 = 9'hdf == r_count_8_io_out ? io_r_223_b : _GEN_2712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2714 = 9'he0 == r_count_8_io_out ? io_r_224_b : _GEN_2713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2715 = 9'he1 == r_count_8_io_out ? io_r_225_b : _GEN_2714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2716 = 9'he2 == r_count_8_io_out ? io_r_226_b : _GEN_2715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2717 = 9'he3 == r_count_8_io_out ? io_r_227_b : _GEN_2716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2718 = 9'he4 == r_count_8_io_out ? io_r_228_b : _GEN_2717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2719 = 9'he5 == r_count_8_io_out ? io_r_229_b : _GEN_2718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2720 = 9'he6 == r_count_8_io_out ? io_r_230_b : _GEN_2719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2721 = 9'he7 == r_count_8_io_out ? io_r_231_b : _GEN_2720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2722 = 9'he8 == r_count_8_io_out ? io_r_232_b : _GEN_2721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2723 = 9'he9 == r_count_8_io_out ? io_r_233_b : _GEN_2722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2724 = 9'hea == r_count_8_io_out ? io_r_234_b : _GEN_2723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2725 = 9'heb == r_count_8_io_out ? io_r_235_b : _GEN_2724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2726 = 9'hec == r_count_8_io_out ? io_r_236_b : _GEN_2725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2727 = 9'hed == r_count_8_io_out ? io_r_237_b : _GEN_2726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2728 = 9'hee == r_count_8_io_out ? io_r_238_b : _GEN_2727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2729 = 9'hef == r_count_8_io_out ? io_r_239_b : _GEN_2728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2730 = 9'hf0 == r_count_8_io_out ? io_r_240_b : _GEN_2729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2731 = 9'hf1 == r_count_8_io_out ? io_r_241_b : _GEN_2730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2732 = 9'hf2 == r_count_8_io_out ? io_r_242_b : _GEN_2731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2733 = 9'hf3 == r_count_8_io_out ? io_r_243_b : _GEN_2732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2734 = 9'hf4 == r_count_8_io_out ? io_r_244_b : _GEN_2733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2735 = 9'hf5 == r_count_8_io_out ? io_r_245_b : _GEN_2734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2736 = 9'hf6 == r_count_8_io_out ? io_r_246_b : _GEN_2735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2737 = 9'hf7 == r_count_8_io_out ? io_r_247_b : _GEN_2736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2738 = 9'hf8 == r_count_8_io_out ? io_r_248_b : _GEN_2737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2739 = 9'hf9 == r_count_8_io_out ? io_r_249_b : _GEN_2738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2740 = 9'hfa == r_count_8_io_out ? io_r_250_b : _GEN_2739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2741 = 9'hfb == r_count_8_io_out ? io_r_251_b : _GEN_2740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2742 = 9'hfc == r_count_8_io_out ? io_r_252_b : _GEN_2741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2743 = 9'hfd == r_count_8_io_out ? io_r_253_b : _GEN_2742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2744 = 9'hfe == r_count_8_io_out ? io_r_254_b : _GEN_2743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2745 = 9'hff == r_count_8_io_out ? io_r_255_b : _GEN_2744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2746 = 9'h100 == r_count_8_io_out ? io_r_256_b : _GEN_2745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2747 = 9'h101 == r_count_8_io_out ? io_r_257_b : _GEN_2746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2748 = 9'h102 == r_count_8_io_out ? io_r_258_b : _GEN_2747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2749 = 9'h103 == r_count_8_io_out ? io_r_259_b : _GEN_2748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2750 = 9'h104 == r_count_8_io_out ? io_r_260_b : _GEN_2749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2751 = 9'h105 == r_count_8_io_out ? io_r_261_b : _GEN_2750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2752 = 9'h106 == r_count_8_io_out ? io_r_262_b : _GEN_2751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2753 = 9'h107 == r_count_8_io_out ? io_r_263_b : _GEN_2752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2754 = 9'h108 == r_count_8_io_out ? io_r_264_b : _GEN_2753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2755 = 9'h109 == r_count_8_io_out ? io_r_265_b : _GEN_2754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2756 = 9'h10a == r_count_8_io_out ? io_r_266_b : _GEN_2755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2757 = 9'h10b == r_count_8_io_out ? io_r_267_b : _GEN_2756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2758 = 9'h10c == r_count_8_io_out ? io_r_268_b : _GEN_2757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2759 = 9'h10d == r_count_8_io_out ? io_r_269_b : _GEN_2758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2760 = 9'h10e == r_count_8_io_out ? io_r_270_b : _GEN_2759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2761 = 9'h10f == r_count_8_io_out ? io_r_271_b : _GEN_2760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2762 = 9'h110 == r_count_8_io_out ? io_r_272_b : _GEN_2761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2763 = 9'h111 == r_count_8_io_out ? io_r_273_b : _GEN_2762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2764 = 9'h112 == r_count_8_io_out ? io_r_274_b : _GEN_2763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2765 = 9'h113 == r_count_8_io_out ? io_r_275_b : _GEN_2764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2766 = 9'h114 == r_count_8_io_out ? io_r_276_b : _GEN_2765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2767 = 9'h115 == r_count_8_io_out ? io_r_277_b : _GEN_2766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2768 = 9'h116 == r_count_8_io_out ? io_r_278_b : _GEN_2767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2769 = 9'h117 == r_count_8_io_out ? io_r_279_b : _GEN_2768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2770 = 9'h118 == r_count_8_io_out ? io_r_280_b : _GEN_2769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2771 = 9'h119 == r_count_8_io_out ? io_r_281_b : _GEN_2770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2772 = 9'h11a == r_count_8_io_out ? io_r_282_b : _GEN_2771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2773 = 9'h11b == r_count_8_io_out ? io_r_283_b : _GEN_2772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2774 = 9'h11c == r_count_8_io_out ? io_r_284_b : _GEN_2773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2775 = 9'h11d == r_count_8_io_out ? io_r_285_b : _GEN_2774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2776 = 9'h11e == r_count_8_io_out ? io_r_286_b : _GEN_2775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2777 = 9'h11f == r_count_8_io_out ? io_r_287_b : _GEN_2776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2778 = 9'h120 == r_count_8_io_out ? io_r_288_b : _GEN_2777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2779 = 9'h121 == r_count_8_io_out ? io_r_289_b : _GEN_2778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2780 = 9'h122 == r_count_8_io_out ? io_r_290_b : _GEN_2779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2781 = 9'h123 == r_count_8_io_out ? io_r_291_b : _GEN_2780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2782 = 9'h124 == r_count_8_io_out ? io_r_292_b : _GEN_2781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2783 = 9'h125 == r_count_8_io_out ? io_r_293_b : _GEN_2782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2784 = 9'h126 == r_count_8_io_out ? io_r_294_b : _GEN_2783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2785 = 9'h127 == r_count_8_io_out ? io_r_295_b : _GEN_2784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2786 = 9'h128 == r_count_8_io_out ? io_r_296_b : _GEN_2785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2787 = 9'h129 == r_count_8_io_out ? io_r_297_b : _GEN_2786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2788 = 9'h12a == r_count_8_io_out ? io_r_298_b : _GEN_2787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2791 = 9'h1 == r_count_9_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2792 = 9'h2 == r_count_9_io_out ? io_r_2_b : _GEN_2791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2793 = 9'h3 == r_count_9_io_out ? io_r_3_b : _GEN_2792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2794 = 9'h4 == r_count_9_io_out ? io_r_4_b : _GEN_2793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2795 = 9'h5 == r_count_9_io_out ? io_r_5_b : _GEN_2794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2796 = 9'h6 == r_count_9_io_out ? io_r_6_b : _GEN_2795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2797 = 9'h7 == r_count_9_io_out ? io_r_7_b : _GEN_2796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2798 = 9'h8 == r_count_9_io_out ? io_r_8_b : _GEN_2797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2799 = 9'h9 == r_count_9_io_out ? io_r_9_b : _GEN_2798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2800 = 9'ha == r_count_9_io_out ? io_r_10_b : _GEN_2799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2801 = 9'hb == r_count_9_io_out ? io_r_11_b : _GEN_2800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2802 = 9'hc == r_count_9_io_out ? io_r_12_b : _GEN_2801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2803 = 9'hd == r_count_9_io_out ? io_r_13_b : _GEN_2802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2804 = 9'he == r_count_9_io_out ? io_r_14_b : _GEN_2803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2805 = 9'hf == r_count_9_io_out ? io_r_15_b : _GEN_2804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2806 = 9'h10 == r_count_9_io_out ? io_r_16_b : _GEN_2805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2807 = 9'h11 == r_count_9_io_out ? io_r_17_b : _GEN_2806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2808 = 9'h12 == r_count_9_io_out ? io_r_18_b : _GEN_2807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2809 = 9'h13 == r_count_9_io_out ? io_r_19_b : _GEN_2808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2810 = 9'h14 == r_count_9_io_out ? io_r_20_b : _GEN_2809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2811 = 9'h15 == r_count_9_io_out ? io_r_21_b : _GEN_2810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2812 = 9'h16 == r_count_9_io_out ? io_r_22_b : _GEN_2811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2813 = 9'h17 == r_count_9_io_out ? io_r_23_b : _GEN_2812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2814 = 9'h18 == r_count_9_io_out ? io_r_24_b : _GEN_2813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2815 = 9'h19 == r_count_9_io_out ? io_r_25_b : _GEN_2814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2816 = 9'h1a == r_count_9_io_out ? io_r_26_b : _GEN_2815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2817 = 9'h1b == r_count_9_io_out ? io_r_27_b : _GEN_2816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2818 = 9'h1c == r_count_9_io_out ? io_r_28_b : _GEN_2817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2819 = 9'h1d == r_count_9_io_out ? io_r_29_b : _GEN_2818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2820 = 9'h1e == r_count_9_io_out ? io_r_30_b : _GEN_2819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2821 = 9'h1f == r_count_9_io_out ? io_r_31_b : _GEN_2820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2822 = 9'h20 == r_count_9_io_out ? io_r_32_b : _GEN_2821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2823 = 9'h21 == r_count_9_io_out ? io_r_33_b : _GEN_2822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2824 = 9'h22 == r_count_9_io_out ? io_r_34_b : _GEN_2823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2825 = 9'h23 == r_count_9_io_out ? io_r_35_b : _GEN_2824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2826 = 9'h24 == r_count_9_io_out ? io_r_36_b : _GEN_2825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2827 = 9'h25 == r_count_9_io_out ? io_r_37_b : _GEN_2826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2828 = 9'h26 == r_count_9_io_out ? io_r_38_b : _GEN_2827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2829 = 9'h27 == r_count_9_io_out ? io_r_39_b : _GEN_2828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2830 = 9'h28 == r_count_9_io_out ? io_r_40_b : _GEN_2829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2831 = 9'h29 == r_count_9_io_out ? io_r_41_b : _GEN_2830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2832 = 9'h2a == r_count_9_io_out ? io_r_42_b : _GEN_2831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2833 = 9'h2b == r_count_9_io_out ? io_r_43_b : _GEN_2832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2834 = 9'h2c == r_count_9_io_out ? io_r_44_b : _GEN_2833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2835 = 9'h2d == r_count_9_io_out ? io_r_45_b : _GEN_2834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2836 = 9'h2e == r_count_9_io_out ? io_r_46_b : _GEN_2835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2837 = 9'h2f == r_count_9_io_out ? io_r_47_b : _GEN_2836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2838 = 9'h30 == r_count_9_io_out ? io_r_48_b : _GEN_2837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2839 = 9'h31 == r_count_9_io_out ? io_r_49_b : _GEN_2838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2840 = 9'h32 == r_count_9_io_out ? io_r_50_b : _GEN_2839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2841 = 9'h33 == r_count_9_io_out ? io_r_51_b : _GEN_2840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2842 = 9'h34 == r_count_9_io_out ? io_r_52_b : _GEN_2841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2843 = 9'h35 == r_count_9_io_out ? io_r_53_b : _GEN_2842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2844 = 9'h36 == r_count_9_io_out ? io_r_54_b : _GEN_2843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2845 = 9'h37 == r_count_9_io_out ? io_r_55_b : _GEN_2844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2846 = 9'h38 == r_count_9_io_out ? io_r_56_b : _GEN_2845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2847 = 9'h39 == r_count_9_io_out ? io_r_57_b : _GEN_2846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2848 = 9'h3a == r_count_9_io_out ? io_r_58_b : _GEN_2847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2849 = 9'h3b == r_count_9_io_out ? io_r_59_b : _GEN_2848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2850 = 9'h3c == r_count_9_io_out ? io_r_60_b : _GEN_2849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2851 = 9'h3d == r_count_9_io_out ? io_r_61_b : _GEN_2850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2852 = 9'h3e == r_count_9_io_out ? io_r_62_b : _GEN_2851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2853 = 9'h3f == r_count_9_io_out ? io_r_63_b : _GEN_2852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2854 = 9'h40 == r_count_9_io_out ? io_r_64_b : _GEN_2853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2855 = 9'h41 == r_count_9_io_out ? io_r_65_b : _GEN_2854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2856 = 9'h42 == r_count_9_io_out ? io_r_66_b : _GEN_2855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2857 = 9'h43 == r_count_9_io_out ? io_r_67_b : _GEN_2856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2858 = 9'h44 == r_count_9_io_out ? io_r_68_b : _GEN_2857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2859 = 9'h45 == r_count_9_io_out ? io_r_69_b : _GEN_2858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2860 = 9'h46 == r_count_9_io_out ? io_r_70_b : _GEN_2859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2861 = 9'h47 == r_count_9_io_out ? io_r_71_b : _GEN_2860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2862 = 9'h48 == r_count_9_io_out ? io_r_72_b : _GEN_2861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2863 = 9'h49 == r_count_9_io_out ? io_r_73_b : _GEN_2862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2864 = 9'h4a == r_count_9_io_out ? io_r_74_b : _GEN_2863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2865 = 9'h4b == r_count_9_io_out ? io_r_75_b : _GEN_2864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2866 = 9'h4c == r_count_9_io_out ? io_r_76_b : _GEN_2865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2867 = 9'h4d == r_count_9_io_out ? io_r_77_b : _GEN_2866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2868 = 9'h4e == r_count_9_io_out ? io_r_78_b : _GEN_2867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2869 = 9'h4f == r_count_9_io_out ? io_r_79_b : _GEN_2868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2870 = 9'h50 == r_count_9_io_out ? io_r_80_b : _GEN_2869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2871 = 9'h51 == r_count_9_io_out ? io_r_81_b : _GEN_2870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2872 = 9'h52 == r_count_9_io_out ? io_r_82_b : _GEN_2871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2873 = 9'h53 == r_count_9_io_out ? io_r_83_b : _GEN_2872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2874 = 9'h54 == r_count_9_io_out ? io_r_84_b : _GEN_2873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2875 = 9'h55 == r_count_9_io_out ? io_r_85_b : _GEN_2874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2876 = 9'h56 == r_count_9_io_out ? io_r_86_b : _GEN_2875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2877 = 9'h57 == r_count_9_io_out ? io_r_87_b : _GEN_2876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2878 = 9'h58 == r_count_9_io_out ? io_r_88_b : _GEN_2877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2879 = 9'h59 == r_count_9_io_out ? io_r_89_b : _GEN_2878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2880 = 9'h5a == r_count_9_io_out ? io_r_90_b : _GEN_2879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2881 = 9'h5b == r_count_9_io_out ? io_r_91_b : _GEN_2880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2882 = 9'h5c == r_count_9_io_out ? io_r_92_b : _GEN_2881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2883 = 9'h5d == r_count_9_io_out ? io_r_93_b : _GEN_2882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2884 = 9'h5e == r_count_9_io_out ? io_r_94_b : _GEN_2883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2885 = 9'h5f == r_count_9_io_out ? io_r_95_b : _GEN_2884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2886 = 9'h60 == r_count_9_io_out ? io_r_96_b : _GEN_2885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2887 = 9'h61 == r_count_9_io_out ? io_r_97_b : _GEN_2886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2888 = 9'h62 == r_count_9_io_out ? io_r_98_b : _GEN_2887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2889 = 9'h63 == r_count_9_io_out ? io_r_99_b : _GEN_2888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2890 = 9'h64 == r_count_9_io_out ? io_r_100_b : _GEN_2889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2891 = 9'h65 == r_count_9_io_out ? io_r_101_b : _GEN_2890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2892 = 9'h66 == r_count_9_io_out ? io_r_102_b : _GEN_2891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2893 = 9'h67 == r_count_9_io_out ? io_r_103_b : _GEN_2892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2894 = 9'h68 == r_count_9_io_out ? io_r_104_b : _GEN_2893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2895 = 9'h69 == r_count_9_io_out ? io_r_105_b : _GEN_2894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2896 = 9'h6a == r_count_9_io_out ? io_r_106_b : _GEN_2895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2897 = 9'h6b == r_count_9_io_out ? io_r_107_b : _GEN_2896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2898 = 9'h6c == r_count_9_io_out ? io_r_108_b : _GEN_2897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2899 = 9'h6d == r_count_9_io_out ? io_r_109_b : _GEN_2898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2900 = 9'h6e == r_count_9_io_out ? io_r_110_b : _GEN_2899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2901 = 9'h6f == r_count_9_io_out ? io_r_111_b : _GEN_2900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2902 = 9'h70 == r_count_9_io_out ? io_r_112_b : _GEN_2901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2903 = 9'h71 == r_count_9_io_out ? io_r_113_b : _GEN_2902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2904 = 9'h72 == r_count_9_io_out ? io_r_114_b : _GEN_2903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2905 = 9'h73 == r_count_9_io_out ? io_r_115_b : _GEN_2904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2906 = 9'h74 == r_count_9_io_out ? io_r_116_b : _GEN_2905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2907 = 9'h75 == r_count_9_io_out ? io_r_117_b : _GEN_2906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2908 = 9'h76 == r_count_9_io_out ? io_r_118_b : _GEN_2907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2909 = 9'h77 == r_count_9_io_out ? io_r_119_b : _GEN_2908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2910 = 9'h78 == r_count_9_io_out ? io_r_120_b : _GEN_2909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2911 = 9'h79 == r_count_9_io_out ? io_r_121_b : _GEN_2910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2912 = 9'h7a == r_count_9_io_out ? io_r_122_b : _GEN_2911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2913 = 9'h7b == r_count_9_io_out ? io_r_123_b : _GEN_2912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2914 = 9'h7c == r_count_9_io_out ? io_r_124_b : _GEN_2913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2915 = 9'h7d == r_count_9_io_out ? io_r_125_b : _GEN_2914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2916 = 9'h7e == r_count_9_io_out ? io_r_126_b : _GEN_2915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2917 = 9'h7f == r_count_9_io_out ? io_r_127_b : _GEN_2916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2918 = 9'h80 == r_count_9_io_out ? io_r_128_b : _GEN_2917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2919 = 9'h81 == r_count_9_io_out ? io_r_129_b : _GEN_2918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2920 = 9'h82 == r_count_9_io_out ? io_r_130_b : _GEN_2919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2921 = 9'h83 == r_count_9_io_out ? io_r_131_b : _GEN_2920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2922 = 9'h84 == r_count_9_io_out ? io_r_132_b : _GEN_2921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2923 = 9'h85 == r_count_9_io_out ? io_r_133_b : _GEN_2922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2924 = 9'h86 == r_count_9_io_out ? io_r_134_b : _GEN_2923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2925 = 9'h87 == r_count_9_io_out ? io_r_135_b : _GEN_2924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2926 = 9'h88 == r_count_9_io_out ? io_r_136_b : _GEN_2925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2927 = 9'h89 == r_count_9_io_out ? io_r_137_b : _GEN_2926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2928 = 9'h8a == r_count_9_io_out ? io_r_138_b : _GEN_2927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2929 = 9'h8b == r_count_9_io_out ? io_r_139_b : _GEN_2928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2930 = 9'h8c == r_count_9_io_out ? io_r_140_b : _GEN_2929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2931 = 9'h8d == r_count_9_io_out ? io_r_141_b : _GEN_2930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2932 = 9'h8e == r_count_9_io_out ? io_r_142_b : _GEN_2931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2933 = 9'h8f == r_count_9_io_out ? io_r_143_b : _GEN_2932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2934 = 9'h90 == r_count_9_io_out ? io_r_144_b : _GEN_2933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2935 = 9'h91 == r_count_9_io_out ? io_r_145_b : _GEN_2934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2936 = 9'h92 == r_count_9_io_out ? io_r_146_b : _GEN_2935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2937 = 9'h93 == r_count_9_io_out ? io_r_147_b : _GEN_2936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2938 = 9'h94 == r_count_9_io_out ? io_r_148_b : _GEN_2937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2939 = 9'h95 == r_count_9_io_out ? io_r_149_b : _GEN_2938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2940 = 9'h96 == r_count_9_io_out ? io_r_150_b : _GEN_2939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2941 = 9'h97 == r_count_9_io_out ? io_r_151_b : _GEN_2940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2942 = 9'h98 == r_count_9_io_out ? io_r_152_b : _GEN_2941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2943 = 9'h99 == r_count_9_io_out ? io_r_153_b : _GEN_2942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2944 = 9'h9a == r_count_9_io_out ? io_r_154_b : _GEN_2943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2945 = 9'h9b == r_count_9_io_out ? io_r_155_b : _GEN_2944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2946 = 9'h9c == r_count_9_io_out ? io_r_156_b : _GEN_2945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2947 = 9'h9d == r_count_9_io_out ? io_r_157_b : _GEN_2946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2948 = 9'h9e == r_count_9_io_out ? io_r_158_b : _GEN_2947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2949 = 9'h9f == r_count_9_io_out ? io_r_159_b : _GEN_2948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2950 = 9'ha0 == r_count_9_io_out ? io_r_160_b : _GEN_2949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2951 = 9'ha1 == r_count_9_io_out ? io_r_161_b : _GEN_2950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2952 = 9'ha2 == r_count_9_io_out ? io_r_162_b : _GEN_2951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2953 = 9'ha3 == r_count_9_io_out ? io_r_163_b : _GEN_2952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2954 = 9'ha4 == r_count_9_io_out ? io_r_164_b : _GEN_2953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2955 = 9'ha5 == r_count_9_io_out ? io_r_165_b : _GEN_2954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2956 = 9'ha6 == r_count_9_io_out ? io_r_166_b : _GEN_2955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2957 = 9'ha7 == r_count_9_io_out ? io_r_167_b : _GEN_2956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2958 = 9'ha8 == r_count_9_io_out ? io_r_168_b : _GEN_2957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2959 = 9'ha9 == r_count_9_io_out ? io_r_169_b : _GEN_2958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2960 = 9'haa == r_count_9_io_out ? io_r_170_b : _GEN_2959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2961 = 9'hab == r_count_9_io_out ? io_r_171_b : _GEN_2960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2962 = 9'hac == r_count_9_io_out ? io_r_172_b : _GEN_2961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2963 = 9'had == r_count_9_io_out ? io_r_173_b : _GEN_2962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2964 = 9'hae == r_count_9_io_out ? io_r_174_b : _GEN_2963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2965 = 9'haf == r_count_9_io_out ? io_r_175_b : _GEN_2964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2966 = 9'hb0 == r_count_9_io_out ? io_r_176_b : _GEN_2965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2967 = 9'hb1 == r_count_9_io_out ? io_r_177_b : _GEN_2966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2968 = 9'hb2 == r_count_9_io_out ? io_r_178_b : _GEN_2967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2969 = 9'hb3 == r_count_9_io_out ? io_r_179_b : _GEN_2968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2970 = 9'hb4 == r_count_9_io_out ? io_r_180_b : _GEN_2969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2971 = 9'hb5 == r_count_9_io_out ? io_r_181_b : _GEN_2970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2972 = 9'hb6 == r_count_9_io_out ? io_r_182_b : _GEN_2971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2973 = 9'hb7 == r_count_9_io_out ? io_r_183_b : _GEN_2972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2974 = 9'hb8 == r_count_9_io_out ? io_r_184_b : _GEN_2973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2975 = 9'hb9 == r_count_9_io_out ? io_r_185_b : _GEN_2974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2976 = 9'hba == r_count_9_io_out ? io_r_186_b : _GEN_2975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2977 = 9'hbb == r_count_9_io_out ? io_r_187_b : _GEN_2976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2978 = 9'hbc == r_count_9_io_out ? io_r_188_b : _GEN_2977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2979 = 9'hbd == r_count_9_io_out ? io_r_189_b : _GEN_2978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2980 = 9'hbe == r_count_9_io_out ? io_r_190_b : _GEN_2979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2981 = 9'hbf == r_count_9_io_out ? io_r_191_b : _GEN_2980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2982 = 9'hc0 == r_count_9_io_out ? io_r_192_b : _GEN_2981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2983 = 9'hc1 == r_count_9_io_out ? io_r_193_b : _GEN_2982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2984 = 9'hc2 == r_count_9_io_out ? io_r_194_b : _GEN_2983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2985 = 9'hc3 == r_count_9_io_out ? io_r_195_b : _GEN_2984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2986 = 9'hc4 == r_count_9_io_out ? io_r_196_b : _GEN_2985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2987 = 9'hc5 == r_count_9_io_out ? io_r_197_b : _GEN_2986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2988 = 9'hc6 == r_count_9_io_out ? io_r_198_b : _GEN_2987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2989 = 9'hc7 == r_count_9_io_out ? io_r_199_b : _GEN_2988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2990 = 9'hc8 == r_count_9_io_out ? io_r_200_b : _GEN_2989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2991 = 9'hc9 == r_count_9_io_out ? io_r_201_b : _GEN_2990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2992 = 9'hca == r_count_9_io_out ? io_r_202_b : _GEN_2991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2993 = 9'hcb == r_count_9_io_out ? io_r_203_b : _GEN_2992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2994 = 9'hcc == r_count_9_io_out ? io_r_204_b : _GEN_2993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2995 = 9'hcd == r_count_9_io_out ? io_r_205_b : _GEN_2994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2996 = 9'hce == r_count_9_io_out ? io_r_206_b : _GEN_2995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2997 = 9'hcf == r_count_9_io_out ? io_r_207_b : _GEN_2996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2998 = 9'hd0 == r_count_9_io_out ? io_r_208_b : _GEN_2997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2999 = 9'hd1 == r_count_9_io_out ? io_r_209_b : _GEN_2998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3000 = 9'hd2 == r_count_9_io_out ? io_r_210_b : _GEN_2999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3001 = 9'hd3 == r_count_9_io_out ? io_r_211_b : _GEN_3000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3002 = 9'hd4 == r_count_9_io_out ? io_r_212_b : _GEN_3001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3003 = 9'hd5 == r_count_9_io_out ? io_r_213_b : _GEN_3002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3004 = 9'hd6 == r_count_9_io_out ? io_r_214_b : _GEN_3003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3005 = 9'hd7 == r_count_9_io_out ? io_r_215_b : _GEN_3004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3006 = 9'hd8 == r_count_9_io_out ? io_r_216_b : _GEN_3005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3007 = 9'hd9 == r_count_9_io_out ? io_r_217_b : _GEN_3006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3008 = 9'hda == r_count_9_io_out ? io_r_218_b : _GEN_3007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3009 = 9'hdb == r_count_9_io_out ? io_r_219_b : _GEN_3008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3010 = 9'hdc == r_count_9_io_out ? io_r_220_b : _GEN_3009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3011 = 9'hdd == r_count_9_io_out ? io_r_221_b : _GEN_3010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3012 = 9'hde == r_count_9_io_out ? io_r_222_b : _GEN_3011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3013 = 9'hdf == r_count_9_io_out ? io_r_223_b : _GEN_3012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3014 = 9'he0 == r_count_9_io_out ? io_r_224_b : _GEN_3013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3015 = 9'he1 == r_count_9_io_out ? io_r_225_b : _GEN_3014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3016 = 9'he2 == r_count_9_io_out ? io_r_226_b : _GEN_3015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3017 = 9'he3 == r_count_9_io_out ? io_r_227_b : _GEN_3016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3018 = 9'he4 == r_count_9_io_out ? io_r_228_b : _GEN_3017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3019 = 9'he5 == r_count_9_io_out ? io_r_229_b : _GEN_3018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3020 = 9'he6 == r_count_9_io_out ? io_r_230_b : _GEN_3019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3021 = 9'he7 == r_count_9_io_out ? io_r_231_b : _GEN_3020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3022 = 9'he8 == r_count_9_io_out ? io_r_232_b : _GEN_3021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3023 = 9'he9 == r_count_9_io_out ? io_r_233_b : _GEN_3022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3024 = 9'hea == r_count_9_io_out ? io_r_234_b : _GEN_3023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3025 = 9'heb == r_count_9_io_out ? io_r_235_b : _GEN_3024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3026 = 9'hec == r_count_9_io_out ? io_r_236_b : _GEN_3025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3027 = 9'hed == r_count_9_io_out ? io_r_237_b : _GEN_3026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3028 = 9'hee == r_count_9_io_out ? io_r_238_b : _GEN_3027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3029 = 9'hef == r_count_9_io_out ? io_r_239_b : _GEN_3028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3030 = 9'hf0 == r_count_9_io_out ? io_r_240_b : _GEN_3029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3031 = 9'hf1 == r_count_9_io_out ? io_r_241_b : _GEN_3030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3032 = 9'hf2 == r_count_9_io_out ? io_r_242_b : _GEN_3031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3033 = 9'hf3 == r_count_9_io_out ? io_r_243_b : _GEN_3032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3034 = 9'hf4 == r_count_9_io_out ? io_r_244_b : _GEN_3033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3035 = 9'hf5 == r_count_9_io_out ? io_r_245_b : _GEN_3034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3036 = 9'hf6 == r_count_9_io_out ? io_r_246_b : _GEN_3035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3037 = 9'hf7 == r_count_9_io_out ? io_r_247_b : _GEN_3036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3038 = 9'hf8 == r_count_9_io_out ? io_r_248_b : _GEN_3037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3039 = 9'hf9 == r_count_9_io_out ? io_r_249_b : _GEN_3038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3040 = 9'hfa == r_count_9_io_out ? io_r_250_b : _GEN_3039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3041 = 9'hfb == r_count_9_io_out ? io_r_251_b : _GEN_3040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3042 = 9'hfc == r_count_9_io_out ? io_r_252_b : _GEN_3041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3043 = 9'hfd == r_count_9_io_out ? io_r_253_b : _GEN_3042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3044 = 9'hfe == r_count_9_io_out ? io_r_254_b : _GEN_3043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3045 = 9'hff == r_count_9_io_out ? io_r_255_b : _GEN_3044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3046 = 9'h100 == r_count_9_io_out ? io_r_256_b : _GEN_3045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3047 = 9'h101 == r_count_9_io_out ? io_r_257_b : _GEN_3046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3048 = 9'h102 == r_count_9_io_out ? io_r_258_b : _GEN_3047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3049 = 9'h103 == r_count_9_io_out ? io_r_259_b : _GEN_3048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3050 = 9'h104 == r_count_9_io_out ? io_r_260_b : _GEN_3049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3051 = 9'h105 == r_count_9_io_out ? io_r_261_b : _GEN_3050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3052 = 9'h106 == r_count_9_io_out ? io_r_262_b : _GEN_3051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3053 = 9'h107 == r_count_9_io_out ? io_r_263_b : _GEN_3052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3054 = 9'h108 == r_count_9_io_out ? io_r_264_b : _GEN_3053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3055 = 9'h109 == r_count_9_io_out ? io_r_265_b : _GEN_3054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3056 = 9'h10a == r_count_9_io_out ? io_r_266_b : _GEN_3055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3057 = 9'h10b == r_count_9_io_out ? io_r_267_b : _GEN_3056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3058 = 9'h10c == r_count_9_io_out ? io_r_268_b : _GEN_3057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3059 = 9'h10d == r_count_9_io_out ? io_r_269_b : _GEN_3058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3060 = 9'h10e == r_count_9_io_out ? io_r_270_b : _GEN_3059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3061 = 9'h10f == r_count_9_io_out ? io_r_271_b : _GEN_3060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3062 = 9'h110 == r_count_9_io_out ? io_r_272_b : _GEN_3061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3063 = 9'h111 == r_count_9_io_out ? io_r_273_b : _GEN_3062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3064 = 9'h112 == r_count_9_io_out ? io_r_274_b : _GEN_3063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3065 = 9'h113 == r_count_9_io_out ? io_r_275_b : _GEN_3064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3066 = 9'h114 == r_count_9_io_out ? io_r_276_b : _GEN_3065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3067 = 9'h115 == r_count_9_io_out ? io_r_277_b : _GEN_3066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3068 = 9'h116 == r_count_9_io_out ? io_r_278_b : _GEN_3067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3069 = 9'h117 == r_count_9_io_out ? io_r_279_b : _GEN_3068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3070 = 9'h118 == r_count_9_io_out ? io_r_280_b : _GEN_3069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3071 = 9'h119 == r_count_9_io_out ? io_r_281_b : _GEN_3070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3072 = 9'h11a == r_count_9_io_out ? io_r_282_b : _GEN_3071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3073 = 9'h11b == r_count_9_io_out ? io_r_283_b : _GEN_3072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3074 = 9'h11c == r_count_9_io_out ? io_r_284_b : _GEN_3073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3075 = 9'h11d == r_count_9_io_out ? io_r_285_b : _GEN_3074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3076 = 9'h11e == r_count_9_io_out ? io_r_286_b : _GEN_3075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3077 = 9'h11f == r_count_9_io_out ? io_r_287_b : _GEN_3076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3078 = 9'h120 == r_count_9_io_out ? io_r_288_b : _GEN_3077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3079 = 9'h121 == r_count_9_io_out ? io_r_289_b : _GEN_3078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3080 = 9'h122 == r_count_9_io_out ? io_r_290_b : _GEN_3079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3081 = 9'h123 == r_count_9_io_out ? io_r_291_b : _GEN_3080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3082 = 9'h124 == r_count_9_io_out ? io_r_292_b : _GEN_3081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3083 = 9'h125 == r_count_9_io_out ? io_r_293_b : _GEN_3082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3084 = 9'h126 == r_count_9_io_out ? io_r_294_b : _GEN_3083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3085 = 9'h127 == r_count_9_io_out ? io_r_295_b : _GEN_3084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3086 = 9'h128 == r_count_9_io_out ? io_r_296_b : _GEN_3085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3087 = 9'h129 == r_count_9_io_out ? io_r_297_b : _GEN_3086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3088 = 9'h12a == r_count_9_io_out ? io_r_298_b : _GEN_3087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3091 = 9'h1 == r_count_10_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3092 = 9'h2 == r_count_10_io_out ? io_r_2_b : _GEN_3091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3093 = 9'h3 == r_count_10_io_out ? io_r_3_b : _GEN_3092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3094 = 9'h4 == r_count_10_io_out ? io_r_4_b : _GEN_3093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3095 = 9'h5 == r_count_10_io_out ? io_r_5_b : _GEN_3094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3096 = 9'h6 == r_count_10_io_out ? io_r_6_b : _GEN_3095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3097 = 9'h7 == r_count_10_io_out ? io_r_7_b : _GEN_3096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3098 = 9'h8 == r_count_10_io_out ? io_r_8_b : _GEN_3097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3099 = 9'h9 == r_count_10_io_out ? io_r_9_b : _GEN_3098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3100 = 9'ha == r_count_10_io_out ? io_r_10_b : _GEN_3099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3101 = 9'hb == r_count_10_io_out ? io_r_11_b : _GEN_3100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3102 = 9'hc == r_count_10_io_out ? io_r_12_b : _GEN_3101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3103 = 9'hd == r_count_10_io_out ? io_r_13_b : _GEN_3102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3104 = 9'he == r_count_10_io_out ? io_r_14_b : _GEN_3103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3105 = 9'hf == r_count_10_io_out ? io_r_15_b : _GEN_3104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3106 = 9'h10 == r_count_10_io_out ? io_r_16_b : _GEN_3105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3107 = 9'h11 == r_count_10_io_out ? io_r_17_b : _GEN_3106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3108 = 9'h12 == r_count_10_io_out ? io_r_18_b : _GEN_3107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3109 = 9'h13 == r_count_10_io_out ? io_r_19_b : _GEN_3108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3110 = 9'h14 == r_count_10_io_out ? io_r_20_b : _GEN_3109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3111 = 9'h15 == r_count_10_io_out ? io_r_21_b : _GEN_3110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3112 = 9'h16 == r_count_10_io_out ? io_r_22_b : _GEN_3111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3113 = 9'h17 == r_count_10_io_out ? io_r_23_b : _GEN_3112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3114 = 9'h18 == r_count_10_io_out ? io_r_24_b : _GEN_3113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3115 = 9'h19 == r_count_10_io_out ? io_r_25_b : _GEN_3114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3116 = 9'h1a == r_count_10_io_out ? io_r_26_b : _GEN_3115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3117 = 9'h1b == r_count_10_io_out ? io_r_27_b : _GEN_3116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3118 = 9'h1c == r_count_10_io_out ? io_r_28_b : _GEN_3117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3119 = 9'h1d == r_count_10_io_out ? io_r_29_b : _GEN_3118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3120 = 9'h1e == r_count_10_io_out ? io_r_30_b : _GEN_3119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3121 = 9'h1f == r_count_10_io_out ? io_r_31_b : _GEN_3120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3122 = 9'h20 == r_count_10_io_out ? io_r_32_b : _GEN_3121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3123 = 9'h21 == r_count_10_io_out ? io_r_33_b : _GEN_3122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3124 = 9'h22 == r_count_10_io_out ? io_r_34_b : _GEN_3123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3125 = 9'h23 == r_count_10_io_out ? io_r_35_b : _GEN_3124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3126 = 9'h24 == r_count_10_io_out ? io_r_36_b : _GEN_3125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3127 = 9'h25 == r_count_10_io_out ? io_r_37_b : _GEN_3126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3128 = 9'h26 == r_count_10_io_out ? io_r_38_b : _GEN_3127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3129 = 9'h27 == r_count_10_io_out ? io_r_39_b : _GEN_3128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3130 = 9'h28 == r_count_10_io_out ? io_r_40_b : _GEN_3129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3131 = 9'h29 == r_count_10_io_out ? io_r_41_b : _GEN_3130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3132 = 9'h2a == r_count_10_io_out ? io_r_42_b : _GEN_3131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3133 = 9'h2b == r_count_10_io_out ? io_r_43_b : _GEN_3132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3134 = 9'h2c == r_count_10_io_out ? io_r_44_b : _GEN_3133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3135 = 9'h2d == r_count_10_io_out ? io_r_45_b : _GEN_3134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3136 = 9'h2e == r_count_10_io_out ? io_r_46_b : _GEN_3135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3137 = 9'h2f == r_count_10_io_out ? io_r_47_b : _GEN_3136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3138 = 9'h30 == r_count_10_io_out ? io_r_48_b : _GEN_3137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3139 = 9'h31 == r_count_10_io_out ? io_r_49_b : _GEN_3138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3140 = 9'h32 == r_count_10_io_out ? io_r_50_b : _GEN_3139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3141 = 9'h33 == r_count_10_io_out ? io_r_51_b : _GEN_3140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3142 = 9'h34 == r_count_10_io_out ? io_r_52_b : _GEN_3141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3143 = 9'h35 == r_count_10_io_out ? io_r_53_b : _GEN_3142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3144 = 9'h36 == r_count_10_io_out ? io_r_54_b : _GEN_3143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3145 = 9'h37 == r_count_10_io_out ? io_r_55_b : _GEN_3144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3146 = 9'h38 == r_count_10_io_out ? io_r_56_b : _GEN_3145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3147 = 9'h39 == r_count_10_io_out ? io_r_57_b : _GEN_3146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3148 = 9'h3a == r_count_10_io_out ? io_r_58_b : _GEN_3147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3149 = 9'h3b == r_count_10_io_out ? io_r_59_b : _GEN_3148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3150 = 9'h3c == r_count_10_io_out ? io_r_60_b : _GEN_3149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3151 = 9'h3d == r_count_10_io_out ? io_r_61_b : _GEN_3150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3152 = 9'h3e == r_count_10_io_out ? io_r_62_b : _GEN_3151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3153 = 9'h3f == r_count_10_io_out ? io_r_63_b : _GEN_3152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3154 = 9'h40 == r_count_10_io_out ? io_r_64_b : _GEN_3153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3155 = 9'h41 == r_count_10_io_out ? io_r_65_b : _GEN_3154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3156 = 9'h42 == r_count_10_io_out ? io_r_66_b : _GEN_3155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3157 = 9'h43 == r_count_10_io_out ? io_r_67_b : _GEN_3156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3158 = 9'h44 == r_count_10_io_out ? io_r_68_b : _GEN_3157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3159 = 9'h45 == r_count_10_io_out ? io_r_69_b : _GEN_3158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3160 = 9'h46 == r_count_10_io_out ? io_r_70_b : _GEN_3159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3161 = 9'h47 == r_count_10_io_out ? io_r_71_b : _GEN_3160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3162 = 9'h48 == r_count_10_io_out ? io_r_72_b : _GEN_3161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3163 = 9'h49 == r_count_10_io_out ? io_r_73_b : _GEN_3162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3164 = 9'h4a == r_count_10_io_out ? io_r_74_b : _GEN_3163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3165 = 9'h4b == r_count_10_io_out ? io_r_75_b : _GEN_3164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3166 = 9'h4c == r_count_10_io_out ? io_r_76_b : _GEN_3165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3167 = 9'h4d == r_count_10_io_out ? io_r_77_b : _GEN_3166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3168 = 9'h4e == r_count_10_io_out ? io_r_78_b : _GEN_3167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3169 = 9'h4f == r_count_10_io_out ? io_r_79_b : _GEN_3168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3170 = 9'h50 == r_count_10_io_out ? io_r_80_b : _GEN_3169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3171 = 9'h51 == r_count_10_io_out ? io_r_81_b : _GEN_3170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3172 = 9'h52 == r_count_10_io_out ? io_r_82_b : _GEN_3171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3173 = 9'h53 == r_count_10_io_out ? io_r_83_b : _GEN_3172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3174 = 9'h54 == r_count_10_io_out ? io_r_84_b : _GEN_3173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3175 = 9'h55 == r_count_10_io_out ? io_r_85_b : _GEN_3174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3176 = 9'h56 == r_count_10_io_out ? io_r_86_b : _GEN_3175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3177 = 9'h57 == r_count_10_io_out ? io_r_87_b : _GEN_3176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3178 = 9'h58 == r_count_10_io_out ? io_r_88_b : _GEN_3177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3179 = 9'h59 == r_count_10_io_out ? io_r_89_b : _GEN_3178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3180 = 9'h5a == r_count_10_io_out ? io_r_90_b : _GEN_3179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3181 = 9'h5b == r_count_10_io_out ? io_r_91_b : _GEN_3180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3182 = 9'h5c == r_count_10_io_out ? io_r_92_b : _GEN_3181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3183 = 9'h5d == r_count_10_io_out ? io_r_93_b : _GEN_3182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3184 = 9'h5e == r_count_10_io_out ? io_r_94_b : _GEN_3183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3185 = 9'h5f == r_count_10_io_out ? io_r_95_b : _GEN_3184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3186 = 9'h60 == r_count_10_io_out ? io_r_96_b : _GEN_3185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3187 = 9'h61 == r_count_10_io_out ? io_r_97_b : _GEN_3186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3188 = 9'h62 == r_count_10_io_out ? io_r_98_b : _GEN_3187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3189 = 9'h63 == r_count_10_io_out ? io_r_99_b : _GEN_3188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3190 = 9'h64 == r_count_10_io_out ? io_r_100_b : _GEN_3189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3191 = 9'h65 == r_count_10_io_out ? io_r_101_b : _GEN_3190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3192 = 9'h66 == r_count_10_io_out ? io_r_102_b : _GEN_3191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3193 = 9'h67 == r_count_10_io_out ? io_r_103_b : _GEN_3192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3194 = 9'h68 == r_count_10_io_out ? io_r_104_b : _GEN_3193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3195 = 9'h69 == r_count_10_io_out ? io_r_105_b : _GEN_3194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3196 = 9'h6a == r_count_10_io_out ? io_r_106_b : _GEN_3195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3197 = 9'h6b == r_count_10_io_out ? io_r_107_b : _GEN_3196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3198 = 9'h6c == r_count_10_io_out ? io_r_108_b : _GEN_3197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3199 = 9'h6d == r_count_10_io_out ? io_r_109_b : _GEN_3198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3200 = 9'h6e == r_count_10_io_out ? io_r_110_b : _GEN_3199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3201 = 9'h6f == r_count_10_io_out ? io_r_111_b : _GEN_3200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3202 = 9'h70 == r_count_10_io_out ? io_r_112_b : _GEN_3201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3203 = 9'h71 == r_count_10_io_out ? io_r_113_b : _GEN_3202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3204 = 9'h72 == r_count_10_io_out ? io_r_114_b : _GEN_3203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3205 = 9'h73 == r_count_10_io_out ? io_r_115_b : _GEN_3204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3206 = 9'h74 == r_count_10_io_out ? io_r_116_b : _GEN_3205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3207 = 9'h75 == r_count_10_io_out ? io_r_117_b : _GEN_3206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3208 = 9'h76 == r_count_10_io_out ? io_r_118_b : _GEN_3207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3209 = 9'h77 == r_count_10_io_out ? io_r_119_b : _GEN_3208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3210 = 9'h78 == r_count_10_io_out ? io_r_120_b : _GEN_3209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3211 = 9'h79 == r_count_10_io_out ? io_r_121_b : _GEN_3210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3212 = 9'h7a == r_count_10_io_out ? io_r_122_b : _GEN_3211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3213 = 9'h7b == r_count_10_io_out ? io_r_123_b : _GEN_3212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3214 = 9'h7c == r_count_10_io_out ? io_r_124_b : _GEN_3213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3215 = 9'h7d == r_count_10_io_out ? io_r_125_b : _GEN_3214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3216 = 9'h7e == r_count_10_io_out ? io_r_126_b : _GEN_3215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3217 = 9'h7f == r_count_10_io_out ? io_r_127_b : _GEN_3216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3218 = 9'h80 == r_count_10_io_out ? io_r_128_b : _GEN_3217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3219 = 9'h81 == r_count_10_io_out ? io_r_129_b : _GEN_3218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3220 = 9'h82 == r_count_10_io_out ? io_r_130_b : _GEN_3219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3221 = 9'h83 == r_count_10_io_out ? io_r_131_b : _GEN_3220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3222 = 9'h84 == r_count_10_io_out ? io_r_132_b : _GEN_3221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3223 = 9'h85 == r_count_10_io_out ? io_r_133_b : _GEN_3222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3224 = 9'h86 == r_count_10_io_out ? io_r_134_b : _GEN_3223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3225 = 9'h87 == r_count_10_io_out ? io_r_135_b : _GEN_3224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3226 = 9'h88 == r_count_10_io_out ? io_r_136_b : _GEN_3225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3227 = 9'h89 == r_count_10_io_out ? io_r_137_b : _GEN_3226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3228 = 9'h8a == r_count_10_io_out ? io_r_138_b : _GEN_3227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3229 = 9'h8b == r_count_10_io_out ? io_r_139_b : _GEN_3228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3230 = 9'h8c == r_count_10_io_out ? io_r_140_b : _GEN_3229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3231 = 9'h8d == r_count_10_io_out ? io_r_141_b : _GEN_3230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3232 = 9'h8e == r_count_10_io_out ? io_r_142_b : _GEN_3231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3233 = 9'h8f == r_count_10_io_out ? io_r_143_b : _GEN_3232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3234 = 9'h90 == r_count_10_io_out ? io_r_144_b : _GEN_3233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3235 = 9'h91 == r_count_10_io_out ? io_r_145_b : _GEN_3234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3236 = 9'h92 == r_count_10_io_out ? io_r_146_b : _GEN_3235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3237 = 9'h93 == r_count_10_io_out ? io_r_147_b : _GEN_3236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3238 = 9'h94 == r_count_10_io_out ? io_r_148_b : _GEN_3237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3239 = 9'h95 == r_count_10_io_out ? io_r_149_b : _GEN_3238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3240 = 9'h96 == r_count_10_io_out ? io_r_150_b : _GEN_3239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3241 = 9'h97 == r_count_10_io_out ? io_r_151_b : _GEN_3240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3242 = 9'h98 == r_count_10_io_out ? io_r_152_b : _GEN_3241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3243 = 9'h99 == r_count_10_io_out ? io_r_153_b : _GEN_3242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3244 = 9'h9a == r_count_10_io_out ? io_r_154_b : _GEN_3243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3245 = 9'h9b == r_count_10_io_out ? io_r_155_b : _GEN_3244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3246 = 9'h9c == r_count_10_io_out ? io_r_156_b : _GEN_3245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3247 = 9'h9d == r_count_10_io_out ? io_r_157_b : _GEN_3246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3248 = 9'h9e == r_count_10_io_out ? io_r_158_b : _GEN_3247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3249 = 9'h9f == r_count_10_io_out ? io_r_159_b : _GEN_3248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3250 = 9'ha0 == r_count_10_io_out ? io_r_160_b : _GEN_3249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3251 = 9'ha1 == r_count_10_io_out ? io_r_161_b : _GEN_3250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3252 = 9'ha2 == r_count_10_io_out ? io_r_162_b : _GEN_3251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3253 = 9'ha3 == r_count_10_io_out ? io_r_163_b : _GEN_3252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3254 = 9'ha4 == r_count_10_io_out ? io_r_164_b : _GEN_3253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3255 = 9'ha5 == r_count_10_io_out ? io_r_165_b : _GEN_3254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3256 = 9'ha6 == r_count_10_io_out ? io_r_166_b : _GEN_3255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3257 = 9'ha7 == r_count_10_io_out ? io_r_167_b : _GEN_3256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3258 = 9'ha8 == r_count_10_io_out ? io_r_168_b : _GEN_3257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3259 = 9'ha9 == r_count_10_io_out ? io_r_169_b : _GEN_3258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3260 = 9'haa == r_count_10_io_out ? io_r_170_b : _GEN_3259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3261 = 9'hab == r_count_10_io_out ? io_r_171_b : _GEN_3260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3262 = 9'hac == r_count_10_io_out ? io_r_172_b : _GEN_3261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3263 = 9'had == r_count_10_io_out ? io_r_173_b : _GEN_3262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3264 = 9'hae == r_count_10_io_out ? io_r_174_b : _GEN_3263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3265 = 9'haf == r_count_10_io_out ? io_r_175_b : _GEN_3264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3266 = 9'hb0 == r_count_10_io_out ? io_r_176_b : _GEN_3265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3267 = 9'hb1 == r_count_10_io_out ? io_r_177_b : _GEN_3266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3268 = 9'hb2 == r_count_10_io_out ? io_r_178_b : _GEN_3267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3269 = 9'hb3 == r_count_10_io_out ? io_r_179_b : _GEN_3268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3270 = 9'hb4 == r_count_10_io_out ? io_r_180_b : _GEN_3269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3271 = 9'hb5 == r_count_10_io_out ? io_r_181_b : _GEN_3270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3272 = 9'hb6 == r_count_10_io_out ? io_r_182_b : _GEN_3271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3273 = 9'hb7 == r_count_10_io_out ? io_r_183_b : _GEN_3272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3274 = 9'hb8 == r_count_10_io_out ? io_r_184_b : _GEN_3273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3275 = 9'hb9 == r_count_10_io_out ? io_r_185_b : _GEN_3274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3276 = 9'hba == r_count_10_io_out ? io_r_186_b : _GEN_3275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3277 = 9'hbb == r_count_10_io_out ? io_r_187_b : _GEN_3276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3278 = 9'hbc == r_count_10_io_out ? io_r_188_b : _GEN_3277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3279 = 9'hbd == r_count_10_io_out ? io_r_189_b : _GEN_3278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3280 = 9'hbe == r_count_10_io_out ? io_r_190_b : _GEN_3279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3281 = 9'hbf == r_count_10_io_out ? io_r_191_b : _GEN_3280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3282 = 9'hc0 == r_count_10_io_out ? io_r_192_b : _GEN_3281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3283 = 9'hc1 == r_count_10_io_out ? io_r_193_b : _GEN_3282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3284 = 9'hc2 == r_count_10_io_out ? io_r_194_b : _GEN_3283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3285 = 9'hc3 == r_count_10_io_out ? io_r_195_b : _GEN_3284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3286 = 9'hc4 == r_count_10_io_out ? io_r_196_b : _GEN_3285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3287 = 9'hc5 == r_count_10_io_out ? io_r_197_b : _GEN_3286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3288 = 9'hc6 == r_count_10_io_out ? io_r_198_b : _GEN_3287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3289 = 9'hc7 == r_count_10_io_out ? io_r_199_b : _GEN_3288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3290 = 9'hc8 == r_count_10_io_out ? io_r_200_b : _GEN_3289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3291 = 9'hc9 == r_count_10_io_out ? io_r_201_b : _GEN_3290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3292 = 9'hca == r_count_10_io_out ? io_r_202_b : _GEN_3291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3293 = 9'hcb == r_count_10_io_out ? io_r_203_b : _GEN_3292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3294 = 9'hcc == r_count_10_io_out ? io_r_204_b : _GEN_3293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3295 = 9'hcd == r_count_10_io_out ? io_r_205_b : _GEN_3294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3296 = 9'hce == r_count_10_io_out ? io_r_206_b : _GEN_3295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3297 = 9'hcf == r_count_10_io_out ? io_r_207_b : _GEN_3296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3298 = 9'hd0 == r_count_10_io_out ? io_r_208_b : _GEN_3297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3299 = 9'hd1 == r_count_10_io_out ? io_r_209_b : _GEN_3298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3300 = 9'hd2 == r_count_10_io_out ? io_r_210_b : _GEN_3299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3301 = 9'hd3 == r_count_10_io_out ? io_r_211_b : _GEN_3300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3302 = 9'hd4 == r_count_10_io_out ? io_r_212_b : _GEN_3301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3303 = 9'hd5 == r_count_10_io_out ? io_r_213_b : _GEN_3302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3304 = 9'hd6 == r_count_10_io_out ? io_r_214_b : _GEN_3303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3305 = 9'hd7 == r_count_10_io_out ? io_r_215_b : _GEN_3304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3306 = 9'hd8 == r_count_10_io_out ? io_r_216_b : _GEN_3305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3307 = 9'hd9 == r_count_10_io_out ? io_r_217_b : _GEN_3306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3308 = 9'hda == r_count_10_io_out ? io_r_218_b : _GEN_3307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3309 = 9'hdb == r_count_10_io_out ? io_r_219_b : _GEN_3308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3310 = 9'hdc == r_count_10_io_out ? io_r_220_b : _GEN_3309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3311 = 9'hdd == r_count_10_io_out ? io_r_221_b : _GEN_3310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3312 = 9'hde == r_count_10_io_out ? io_r_222_b : _GEN_3311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3313 = 9'hdf == r_count_10_io_out ? io_r_223_b : _GEN_3312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3314 = 9'he0 == r_count_10_io_out ? io_r_224_b : _GEN_3313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3315 = 9'he1 == r_count_10_io_out ? io_r_225_b : _GEN_3314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3316 = 9'he2 == r_count_10_io_out ? io_r_226_b : _GEN_3315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3317 = 9'he3 == r_count_10_io_out ? io_r_227_b : _GEN_3316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3318 = 9'he4 == r_count_10_io_out ? io_r_228_b : _GEN_3317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3319 = 9'he5 == r_count_10_io_out ? io_r_229_b : _GEN_3318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3320 = 9'he6 == r_count_10_io_out ? io_r_230_b : _GEN_3319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3321 = 9'he7 == r_count_10_io_out ? io_r_231_b : _GEN_3320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3322 = 9'he8 == r_count_10_io_out ? io_r_232_b : _GEN_3321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3323 = 9'he9 == r_count_10_io_out ? io_r_233_b : _GEN_3322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3324 = 9'hea == r_count_10_io_out ? io_r_234_b : _GEN_3323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3325 = 9'heb == r_count_10_io_out ? io_r_235_b : _GEN_3324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3326 = 9'hec == r_count_10_io_out ? io_r_236_b : _GEN_3325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3327 = 9'hed == r_count_10_io_out ? io_r_237_b : _GEN_3326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3328 = 9'hee == r_count_10_io_out ? io_r_238_b : _GEN_3327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3329 = 9'hef == r_count_10_io_out ? io_r_239_b : _GEN_3328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3330 = 9'hf0 == r_count_10_io_out ? io_r_240_b : _GEN_3329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3331 = 9'hf1 == r_count_10_io_out ? io_r_241_b : _GEN_3330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3332 = 9'hf2 == r_count_10_io_out ? io_r_242_b : _GEN_3331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3333 = 9'hf3 == r_count_10_io_out ? io_r_243_b : _GEN_3332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3334 = 9'hf4 == r_count_10_io_out ? io_r_244_b : _GEN_3333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3335 = 9'hf5 == r_count_10_io_out ? io_r_245_b : _GEN_3334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3336 = 9'hf6 == r_count_10_io_out ? io_r_246_b : _GEN_3335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3337 = 9'hf7 == r_count_10_io_out ? io_r_247_b : _GEN_3336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3338 = 9'hf8 == r_count_10_io_out ? io_r_248_b : _GEN_3337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3339 = 9'hf9 == r_count_10_io_out ? io_r_249_b : _GEN_3338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3340 = 9'hfa == r_count_10_io_out ? io_r_250_b : _GEN_3339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3341 = 9'hfb == r_count_10_io_out ? io_r_251_b : _GEN_3340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3342 = 9'hfc == r_count_10_io_out ? io_r_252_b : _GEN_3341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3343 = 9'hfd == r_count_10_io_out ? io_r_253_b : _GEN_3342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3344 = 9'hfe == r_count_10_io_out ? io_r_254_b : _GEN_3343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3345 = 9'hff == r_count_10_io_out ? io_r_255_b : _GEN_3344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3346 = 9'h100 == r_count_10_io_out ? io_r_256_b : _GEN_3345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3347 = 9'h101 == r_count_10_io_out ? io_r_257_b : _GEN_3346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3348 = 9'h102 == r_count_10_io_out ? io_r_258_b : _GEN_3347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3349 = 9'h103 == r_count_10_io_out ? io_r_259_b : _GEN_3348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3350 = 9'h104 == r_count_10_io_out ? io_r_260_b : _GEN_3349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3351 = 9'h105 == r_count_10_io_out ? io_r_261_b : _GEN_3350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3352 = 9'h106 == r_count_10_io_out ? io_r_262_b : _GEN_3351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3353 = 9'h107 == r_count_10_io_out ? io_r_263_b : _GEN_3352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3354 = 9'h108 == r_count_10_io_out ? io_r_264_b : _GEN_3353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3355 = 9'h109 == r_count_10_io_out ? io_r_265_b : _GEN_3354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3356 = 9'h10a == r_count_10_io_out ? io_r_266_b : _GEN_3355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3357 = 9'h10b == r_count_10_io_out ? io_r_267_b : _GEN_3356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3358 = 9'h10c == r_count_10_io_out ? io_r_268_b : _GEN_3357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3359 = 9'h10d == r_count_10_io_out ? io_r_269_b : _GEN_3358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3360 = 9'h10e == r_count_10_io_out ? io_r_270_b : _GEN_3359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3361 = 9'h10f == r_count_10_io_out ? io_r_271_b : _GEN_3360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3362 = 9'h110 == r_count_10_io_out ? io_r_272_b : _GEN_3361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3363 = 9'h111 == r_count_10_io_out ? io_r_273_b : _GEN_3362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3364 = 9'h112 == r_count_10_io_out ? io_r_274_b : _GEN_3363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3365 = 9'h113 == r_count_10_io_out ? io_r_275_b : _GEN_3364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3366 = 9'h114 == r_count_10_io_out ? io_r_276_b : _GEN_3365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3367 = 9'h115 == r_count_10_io_out ? io_r_277_b : _GEN_3366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3368 = 9'h116 == r_count_10_io_out ? io_r_278_b : _GEN_3367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3369 = 9'h117 == r_count_10_io_out ? io_r_279_b : _GEN_3368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3370 = 9'h118 == r_count_10_io_out ? io_r_280_b : _GEN_3369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3371 = 9'h119 == r_count_10_io_out ? io_r_281_b : _GEN_3370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3372 = 9'h11a == r_count_10_io_out ? io_r_282_b : _GEN_3371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3373 = 9'h11b == r_count_10_io_out ? io_r_283_b : _GEN_3372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3374 = 9'h11c == r_count_10_io_out ? io_r_284_b : _GEN_3373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3375 = 9'h11d == r_count_10_io_out ? io_r_285_b : _GEN_3374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3376 = 9'h11e == r_count_10_io_out ? io_r_286_b : _GEN_3375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3377 = 9'h11f == r_count_10_io_out ? io_r_287_b : _GEN_3376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3378 = 9'h120 == r_count_10_io_out ? io_r_288_b : _GEN_3377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3379 = 9'h121 == r_count_10_io_out ? io_r_289_b : _GEN_3378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3380 = 9'h122 == r_count_10_io_out ? io_r_290_b : _GEN_3379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3381 = 9'h123 == r_count_10_io_out ? io_r_291_b : _GEN_3380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3382 = 9'h124 == r_count_10_io_out ? io_r_292_b : _GEN_3381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3383 = 9'h125 == r_count_10_io_out ? io_r_293_b : _GEN_3382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3384 = 9'h126 == r_count_10_io_out ? io_r_294_b : _GEN_3383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3385 = 9'h127 == r_count_10_io_out ? io_r_295_b : _GEN_3384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3386 = 9'h128 == r_count_10_io_out ? io_r_296_b : _GEN_3385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3387 = 9'h129 == r_count_10_io_out ? io_r_297_b : _GEN_3386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3388 = 9'h12a == r_count_10_io_out ? io_r_298_b : _GEN_3387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3391 = 9'h1 == r_count_11_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3392 = 9'h2 == r_count_11_io_out ? io_r_2_b : _GEN_3391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3393 = 9'h3 == r_count_11_io_out ? io_r_3_b : _GEN_3392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3394 = 9'h4 == r_count_11_io_out ? io_r_4_b : _GEN_3393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3395 = 9'h5 == r_count_11_io_out ? io_r_5_b : _GEN_3394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3396 = 9'h6 == r_count_11_io_out ? io_r_6_b : _GEN_3395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3397 = 9'h7 == r_count_11_io_out ? io_r_7_b : _GEN_3396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3398 = 9'h8 == r_count_11_io_out ? io_r_8_b : _GEN_3397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3399 = 9'h9 == r_count_11_io_out ? io_r_9_b : _GEN_3398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3400 = 9'ha == r_count_11_io_out ? io_r_10_b : _GEN_3399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3401 = 9'hb == r_count_11_io_out ? io_r_11_b : _GEN_3400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3402 = 9'hc == r_count_11_io_out ? io_r_12_b : _GEN_3401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3403 = 9'hd == r_count_11_io_out ? io_r_13_b : _GEN_3402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3404 = 9'he == r_count_11_io_out ? io_r_14_b : _GEN_3403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3405 = 9'hf == r_count_11_io_out ? io_r_15_b : _GEN_3404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3406 = 9'h10 == r_count_11_io_out ? io_r_16_b : _GEN_3405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3407 = 9'h11 == r_count_11_io_out ? io_r_17_b : _GEN_3406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3408 = 9'h12 == r_count_11_io_out ? io_r_18_b : _GEN_3407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3409 = 9'h13 == r_count_11_io_out ? io_r_19_b : _GEN_3408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3410 = 9'h14 == r_count_11_io_out ? io_r_20_b : _GEN_3409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3411 = 9'h15 == r_count_11_io_out ? io_r_21_b : _GEN_3410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3412 = 9'h16 == r_count_11_io_out ? io_r_22_b : _GEN_3411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3413 = 9'h17 == r_count_11_io_out ? io_r_23_b : _GEN_3412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3414 = 9'h18 == r_count_11_io_out ? io_r_24_b : _GEN_3413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3415 = 9'h19 == r_count_11_io_out ? io_r_25_b : _GEN_3414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3416 = 9'h1a == r_count_11_io_out ? io_r_26_b : _GEN_3415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3417 = 9'h1b == r_count_11_io_out ? io_r_27_b : _GEN_3416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3418 = 9'h1c == r_count_11_io_out ? io_r_28_b : _GEN_3417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3419 = 9'h1d == r_count_11_io_out ? io_r_29_b : _GEN_3418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3420 = 9'h1e == r_count_11_io_out ? io_r_30_b : _GEN_3419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3421 = 9'h1f == r_count_11_io_out ? io_r_31_b : _GEN_3420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3422 = 9'h20 == r_count_11_io_out ? io_r_32_b : _GEN_3421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3423 = 9'h21 == r_count_11_io_out ? io_r_33_b : _GEN_3422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3424 = 9'h22 == r_count_11_io_out ? io_r_34_b : _GEN_3423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3425 = 9'h23 == r_count_11_io_out ? io_r_35_b : _GEN_3424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3426 = 9'h24 == r_count_11_io_out ? io_r_36_b : _GEN_3425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3427 = 9'h25 == r_count_11_io_out ? io_r_37_b : _GEN_3426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3428 = 9'h26 == r_count_11_io_out ? io_r_38_b : _GEN_3427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3429 = 9'h27 == r_count_11_io_out ? io_r_39_b : _GEN_3428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3430 = 9'h28 == r_count_11_io_out ? io_r_40_b : _GEN_3429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3431 = 9'h29 == r_count_11_io_out ? io_r_41_b : _GEN_3430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3432 = 9'h2a == r_count_11_io_out ? io_r_42_b : _GEN_3431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3433 = 9'h2b == r_count_11_io_out ? io_r_43_b : _GEN_3432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3434 = 9'h2c == r_count_11_io_out ? io_r_44_b : _GEN_3433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3435 = 9'h2d == r_count_11_io_out ? io_r_45_b : _GEN_3434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3436 = 9'h2e == r_count_11_io_out ? io_r_46_b : _GEN_3435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3437 = 9'h2f == r_count_11_io_out ? io_r_47_b : _GEN_3436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3438 = 9'h30 == r_count_11_io_out ? io_r_48_b : _GEN_3437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3439 = 9'h31 == r_count_11_io_out ? io_r_49_b : _GEN_3438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3440 = 9'h32 == r_count_11_io_out ? io_r_50_b : _GEN_3439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3441 = 9'h33 == r_count_11_io_out ? io_r_51_b : _GEN_3440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3442 = 9'h34 == r_count_11_io_out ? io_r_52_b : _GEN_3441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3443 = 9'h35 == r_count_11_io_out ? io_r_53_b : _GEN_3442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3444 = 9'h36 == r_count_11_io_out ? io_r_54_b : _GEN_3443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3445 = 9'h37 == r_count_11_io_out ? io_r_55_b : _GEN_3444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3446 = 9'h38 == r_count_11_io_out ? io_r_56_b : _GEN_3445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3447 = 9'h39 == r_count_11_io_out ? io_r_57_b : _GEN_3446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3448 = 9'h3a == r_count_11_io_out ? io_r_58_b : _GEN_3447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3449 = 9'h3b == r_count_11_io_out ? io_r_59_b : _GEN_3448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3450 = 9'h3c == r_count_11_io_out ? io_r_60_b : _GEN_3449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3451 = 9'h3d == r_count_11_io_out ? io_r_61_b : _GEN_3450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3452 = 9'h3e == r_count_11_io_out ? io_r_62_b : _GEN_3451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3453 = 9'h3f == r_count_11_io_out ? io_r_63_b : _GEN_3452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3454 = 9'h40 == r_count_11_io_out ? io_r_64_b : _GEN_3453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3455 = 9'h41 == r_count_11_io_out ? io_r_65_b : _GEN_3454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3456 = 9'h42 == r_count_11_io_out ? io_r_66_b : _GEN_3455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3457 = 9'h43 == r_count_11_io_out ? io_r_67_b : _GEN_3456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3458 = 9'h44 == r_count_11_io_out ? io_r_68_b : _GEN_3457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3459 = 9'h45 == r_count_11_io_out ? io_r_69_b : _GEN_3458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3460 = 9'h46 == r_count_11_io_out ? io_r_70_b : _GEN_3459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3461 = 9'h47 == r_count_11_io_out ? io_r_71_b : _GEN_3460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3462 = 9'h48 == r_count_11_io_out ? io_r_72_b : _GEN_3461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3463 = 9'h49 == r_count_11_io_out ? io_r_73_b : _GEN_3462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3464 = 9'h4a == r_count_11_io_out ? io_r_74_b : _GEN_3463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3465 = 9'h4b == r_count_11_io_out ? io_r_75_b : _GEN_3464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3466 = 9'h4c == r_count_11_io_out ? io_r_76_b : _GEN_3465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3467 = 9'h4d == r_count_11_io_out ? io_r_77_b : _GEN_3466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3468 = 9'h4e == r_count_11_io_out ? io_r_78_b : _GEN_3467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3469 = 9'h4f == r_count_11_io_out ? io_r_79_b : _GEN_3468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3470 = 9'h50 == r_count_11_io_out ? io_r_80_b : _GEN_3469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3471 = 9'h51 == r_count_11_io_out ? io_r_81_b : _GEN_3470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3472 = 9'h52 == r_count_11_io_out ? io_r_82_b : _GEN_3471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3473 = 9'h53 == r_count_11_io_out ? io_r_83_b : _GEN_3472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3474 = 9'h54 == r_count_11_io_out ? io_r_84_b : _GEN_3473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3475 = 9'h55 == r_count_11_io_out ? io_r_85_b : _GEN_3474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3476 = 9'h56 == r_count_11_io_out ? io_r_86_b : _GEN_3475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3477 = 9'h57 == r_count_11_io_out ? io_r_87_b : _GEN_3476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3478 = 9'h58 == r_count_11_io_out ? io_r_88_b : _GEN_3477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3479 = 9'h59 == r_count_11_io_out ? io_r_89_b : _GEN_3478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3480 = 9'h5a == r_count_11_io_out ? io_r_90_b : _GEN_3479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3481 = 9'h5b == r_count_11_io_out ? io_r_91_b : _GEN_3480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3482 = 9'h5c == r_count_11_io_out ? io_r_92_b : _GEN_3481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3483 = 9'h5d == r_count_11_io_out ? io_r_93_b : _GEN_3482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3484 = 9'h5e == r_count_11_io_out ? io_r_94_b : _GEN_3483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3485 = 9'h5f == r_count_11_io_out ? io_r_95_b : _GEN_3484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3486 = 9'h60 == r_count_11_io_out ? io_r_96_b : _GEN_3485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3487 = 9'h61 == r_count_11_io_out ? io_r_97_b : _GEN_3486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3488 = 9'h62 == r_count_11_io_out ? io_r_98_b : _GEN_3487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3489 = 9'h63 == r_count_11_io_out ? io_r_99_b : _GEN_3488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3490 = 9'h64 == r_count_11_io_out ? io_r_100_b : _GEN_3489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3491 = 9'h65 == r_count_11_io_out ? io_r_101_b : _GEN_3490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3492 = 9'h66 == r_count_11_io_out ? io_r_102_b : _GEN_3491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3493 = 9'h67 == r_count_11_io_out ? io_r_103_b : _GEN_3492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3494 = 9'h68 == r_count_11_io_out ? io_r_104_b : _GEN_3493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3495 = 9'h69 == r_count_11_io_out ? io_r_105_b : _GEN_3494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3496 = 9'h6a == r_count_11_io_out ? io_r_106_b : _GEN_3495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3497 = 9'h6b == r_count_11_io_out ? io_r_107_b : _GEN_3496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3498 = 9'h6c == r_count_11_io_out ? io_r_108_b : _GEN_3497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3499 = 9'h6d == r_count_11_io_out ? io_r_109_b : _GEN_3498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3500 = 9'h6e == r_count_11_io_out ? io_r_110_b : _GEN_3499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3501 = 9'h6f == r_count_11_io_out ? io_r_111_b : _GEN_3500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3502 = 9'h70 == r_count_11_io_out ? io_r_112_b : _GEN_3501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3503 = 9'h71 == r_count_11_io_out ? io_r_113_b : _GEN_3502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3504 = 9'h72 == r_count_11_io_out ? io_r_114_b : _GEN_3503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3505 = 9'h73 == r_count_11_io_out ? io_r_115_b : _GEN_3504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3506 = 9'h74 == r_count_11_io_out ? io_r_116_b : _GEN_3505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3507 = 9'h75 == r_count_11_io_out ? io_r_117_b : _GEN_3506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3508 = 9'h76 == r_count_11_io_out ? io_r_118_b : _GEN_3507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3509 = 9'h77 == r_count_11_io_out ? io_r_119_b : _GEN_3508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3510 = 9'h78 == r_count_11_io_out ? io_r_120_b : _GEN_3509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3511 = 9'h79 == r_count_11_io_out ? io_r_121_b : _GEN_3510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3512 = 9'h7a == r_count_11_io_out ? io_r_122_b : _GEN_3511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3513 = 9'h7b == r_count_11_io_out ? io_r_123_b : _GEN_3512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3514 = 9'h7c == r_count_11_io_out ? io_r_124_b : _GEN_3513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3515 = 9'h7d == r_count_11_io_out ? io_r_125_b : _GEN_3514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3516 = 9'h7e == r_count_11_io_out ? io_r_126_b : _GEN_3515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3517 = 9'h7f == r_count_11_io_out ? io_r_127_b : _GEN_3516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3518 = 9'h80 == r_count_11_io_out ? io_r_128_b : _GEN_3517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3519 = 9'h81 == r_count_11_io_out ? io_r_129_b : _GEN_3518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3520 = 9'h82 == r_count_11_io_out ? io_r_130_b : _GEN_3519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3521 = 9'h83 == r_count_11_io_out ? io_r_131_b : _GEN_3520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3522 = 9'h84 == r_count_11_io_out ? io_r_132_b : _GEN_3521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3523 = 9'h85 == r_count_11_io_out ? io_r_133_b : _GEN_3522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3524 = 9'h86 == r_count_11_io_out ? io_r_134_b : _GEN_3523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3525 = 9'h87 == r_count_11_io_out ? io_r_135_b : _GEN_3524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3526 = 9'h88 == r_count_11_io_out ? io_r_136_b : _GEN_3525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3527 = 9'h89 == r_count_11_io_out ? io_r_137_b : _GEN_3526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3528 = 9'h8a == r_count_11_io_out ? io_r_138_b : _GEN_3527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3529 = 9'h8b == r_count_11_io_out ? io_r_139_b : _GEN_3528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3530 = 9'h8c == r_count_11_io_out ? io_r_140_b : _GEN_3529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3531 = 9'h8d == r_count_11_io_out ? io_r_141_b : _GEN_3530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3532 = 9'h8e == r_count_11_io_out ? io_r_142_b : _GEN_3531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3533 = 9'h8f == r_count_11_io_out ? io_r_143_b : _GEN_3532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3534 = 9'h90 == r_count_11_io_out ? io_r_144_b : _GEN_3533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3535 = 9'h91 == r_count_11_io_out ? io_r_145_b : _GEN_3534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3536 = 9'h92 == r_count_11_io_out ? io_r_146_b : _GEN_3535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3537 = 9'h93 == r_count_11_io_out ? io_r_147_b : _GEN_3536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3538 = 9'h94 == r_count_11_io_out ? io_r_148_b : _GEN_3537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3539 = 9'h95 == r_count_11_io_out ? io_r_149_b : _GEN_3538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3540 = 9'h96 == r_count_11_io_out ? io_r_150_b : _GEN_3539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3541 = 9'h97 == r_count_11_io_out ? io_r_151_b : _GEN_3540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3542 = 9'h98 == r_count_11_io_out ? io_r_152_b : _GEN_3541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3543 = 9'h99 == r_count_11_io_out ? io_r_153_b : _GEN_3542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3544 = 9'h9a == r_count_11_io_out ? io_r_154_b : _GEN_3543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3545 = 9'h9b == r_count_11_io_out ? io_r_155_b : _GEN_3544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3546 = 9'h9c == r_count_11_io_out ? io_r_156_b : _GEN_3545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3547 = 9'h9d == r_count_11_io_out ? io_r_157_b : _GEN_3546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3548 = 9'h9e == r_count_11_io_out ? io_r_158_b : _GEN_3547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3549 = 9'h9f == r_count_11_io_out ? io_r_159_b : _GEN_3548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3550 = 9'ha0 == r_count_11_io_out ? io_r_160_b : _GEN_3549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3551 = 9'ha1 == r_count_11_io_out ? io_r_161_b : _GEN_3550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3552 = 9'ha2 == r_count_11_io_out ? io_r_162_b : _GEN_3551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3553 = 9'ha3 == r_count_11_io_out ? io_r_163_b : _GEN_3552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3554 = 9'ha4 == r_count_11_io_out ? io_r_164_b : _GEN_3553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3555 = 9'ha5 == r_count_11_io_out ? io_r_165_b : _GEN_3554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3556 = 9'ha6 == r_count_11_io_out ? io_r_166_b : _GEN_3555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3557 = 9'ha7 == r_count_11_io_out ? io_r_167_b : _GEN_3556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3558 = 9'ha8 == r_count_11_io_out ? io_r_168_b : _GEN_3557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3559 = 9'ha9 == r_count_11_io_out ? io_r_169_b : _GEN_3558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3560 = 9'haa == r_count_11_io_out ? io_r_170_b : _GEN_3559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3561 = 9'hab == r_count_11_io_out ? io_r_171_b : _GEN_3560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3562 = 9'hac == r_count_11_io_out ? io_r_172_b : _GEN_3561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3563 = 9'had == r_count_11_io_out ? io_r_173_b : _GEN_3562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3564 = 9'hae == r_count_11_io_out ? io_r_174_b : _GEN_3563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3565 = 9'haf == r_count_11_io_out ? io_r_175_b : _GEN_3564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3566 = 9'hb0 == r_count_11_io_out ? io_r_176_b : _GEN_3565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3567 = 9'hb1 == r_count_11_io_out ? io_r_177_b : _GEN_3566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3568 = 9'hb2 == r_count_11_io_out ? io_r_178_b : _GEN_3567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3569 = 9'hb3 == r_count_11_io_out ? io_r_179_b : _GEN_3568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3570 = 9'hb4 == r_count_11_io_out ? io_r_180_b : _GEN_3569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3571 = 9'hb5 == r_count_11_io_out ? io_r_181_b : _GEN_3570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3572 = 9'hb6 == r_count_11_io_out ? io_r_182_b : _GEN_3571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3573 = 9'hb7 == r_count_11_io_out ? io_r_183_b : _GEN_3572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3574 = 9'hb8 == r_count_11_io_out ? io_r_184_b : _GEN_3573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3575 = 9'hb9 == r_count_11_io_out ? io_r_185_b : _GEN_3574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3576 = 9'hba == r_count_11_io_out ? io_r_186_b : _GEN_3575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3577 = 9'hbb == r_count_11_io_out ? io_r_187_b : _GEN_3576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3578 = 9'hbc == r_count_11_io_out ? io_r_188_b : _GEN_3577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3579 = 9'hbd == r_count_11_io_out ? io_r_189_b : _GEN_3578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3580 = 9'hbe == r_count_11_io_out ? io_r_190_b : _GEN_3579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3581 = 9'hbf == r_count_11_io_out ? io_r_191_b : _GEN_3580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3582 = 9'hc0 == r_count_11_io_out ? io_r_192_b : _GEN_3581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3583 = 9'hc1 == r_count_11_io_out ? io_r_193_b : _GEN_3582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3584 = 9'hc2 == r_count_11_io_out ? io_r_194_b : _GEN_3583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3585 = 9'hc3 == r_count_11_io_out ? io_r_195_b : _GEN_3584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3586 = 9'hc4 == r_count_11_io_out ? io_r_196_b : _GEN_3585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3587 = 9'hc5 == r_count_11_io_out ? io_r_197_b : _GEN_3586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3588 = 9'hc6 == r_count_11_io_out ? io_r_198_b : _GEN_3587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3589 = 9'hc7 == r_count_11_io_out ? io_r_199_b : _GEN_3588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3590 = 9'hc8 == r_count_11_io_out ? io_r_200_b : _GEN_3589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3591 = 9'hc9 == r_count_11_io_out ? io_r_201_b : _GEN_3590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3592 = 9'hca == r_count_11_io_out ? io_r_202_b : _GEN_3591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3593 = 9'hcb == r_count_11_io_out ? io_r_203_b : _GEN_3592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3594 = 9'hcc == r_count_11_io_out ? io_r_204_b : _GEN_3593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3595 = 9'hcd == r_count_11_io_out ? io_r_205_b : _GEN_3594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3596 = 9'hce == r_count_11_io_out ? io_r_206_b : _GEN_3595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3597 = 9'hcf == r_count_11_io_out ? io_r_207_b : _GEN_3596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3598 = 9'hd0 == r_count_11_io_out ? io_r_208_b : _GEN_3597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3599 = 9'hd1 == r_count_11_io_out ? io_r_209_b : _GEN_3598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3600 = 9'hd2 == r_count_11_io_out ? io_r_210_b : _GEN_3599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3601 = 9'hd3 == r_count_11_io_out ? io_r_211_b : _GEN_3600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3602 = 9'hd4 == r_count_11_io_out ? io_r_212_b : _GEN_3601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3603 = 9'hd5 == r_count_11_io_out ? io_r_213_b : _GEN_3602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3604 = 9'hd6 == r_count_11_io_out ? io_r_214_b : _GEN_3603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3605 = 9'hd7 == r_count_11_io_out ? io_r_215_b : _GEN_3604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3606 = 9'hd8 == r_count_11_io_out ? io_r_216_b : _GEN_3605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3607 = 9'hd9 == r_count_11_io_out ? io_r_217_b : _GEN_3606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3608 = 9'hda == r_count_11_io_out ? io_r_218_b : _GEN_3607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3609 = 9'hdb == r_count_11_io_out ? io_r_219_b : _GEN_3608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3610 = 9'hdc == r_count_11_io_out ? io_r_220_b : _GEN_3609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3611 = 9'hdd == r_count_11_io_out ? io_r_221_b : _GEN_3610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3612 = 9'hde == r_count_11_io_out ? io_r_222_b : _GEN_3611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3613 = 9'hdf == r_count_11_io_out ? io_r_223_b : _GEN_3612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3614 = 9'he0 == r_count_11_io_out ? io_r_224_b : _GEN_3613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3615 = 9'he1 == r_count_11_io_out ? io_r_225_b : _GEN_3614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3616 = 9'he2 == r_count_11_io_out ? io_r_226_b : _GEN_3615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3617 = 9'he3 == r_count_11_io_out ? io_r_227_b : _GEN_3616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3618 = 9'he4 == r_count_11_io_out ? io_r_228_b : _GEN_3617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3619 = 9'he5 == r_count_11_io_out ? io_r_229_b : _GEN_3618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3620 = 9'he6 == r_count_11_io_out ? io_r_230_b : _GEN_3619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3621 = 9'he7 == r_count_11_io_out ? io_r_231_b : _GEN_3620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3622 = 9'he8 == r_count_11_io_out ? io_r_232_b : _GEN_3621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3623 = 9'he9 == r_count_11_io_out ? io_r_233_b : _GEN_3622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3624 = 9'hea == r_count_11_io_out ? io_r_234_b : _GEN_3623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3625 = 9'heb == r_count_11_io_out ? io_r_235_b : _GEN_3624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3626 = 9'hec == r_count_11_io_out ? io_r_236_b : _GEN_3625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3627 = 9'hed == r_count_11_io_out ? io_r_237_b : _GEN_3626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3628 = 9'hee == r_count_11_io_out ? io_r_238_b : _GEN_3627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3629 = 9'hef == r_count_11_io_out ? io_r_239_b : _GEN_3628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3630 = 9'hf0 == r_count_11_io_out ? io_r_240_b : _GEN_3629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3631 = 9'hf1 == r_count_11_io_out ? io_r_241_b : _GEN_3630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3632 = 9'hf2 == r_count_11_io_out ? io_r_242_b : _GEN_3631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3633 = 9'hf3 == r_count_11_io_out ? io_r_243_b : _GEN_3632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3634 = 9'hf4 == r_count_11_io_out ? io_r_244_b : _GEN_3633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3635 = 9'hf5 == r_count_11_io_out ? io_r_245_b : _GEN_3634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3636 = 9'hf6 == r_count_11_io_out ? io_r_246_b : _GEN_3635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3637 = 9'hf7 == r_count_11_io_out ? io_r_247_b : _GEN_3636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3638 = 9'hf8 == r_count_11_io_out ? io_r_248_b : _GEN_3637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3639 = 9'hf9 == r_count_11_io_out ? io_r_249_b : _GEN_3638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3640 = 9'hfa == r_count_11_io_out ? io_r_250_b : _GEN_3639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3641 = 9'hfb == r_count_11_io_out ? io_r_251_b : _GEN_3640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3642 = 9'hfc == r_count_11_io_out ? io_r_252_b : _GEN_3641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3643 = 9'hfd == r_count_11_io_out ? io_r_253_b : _GEN_3642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3644 = 9'hfe == r_count_11_io_out ? io_r_254_b : _GEN_3643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3645 = 9'hff == r_count_11_io_out ? io_r_255_b : _GEN_3644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3646 = 9'h100 == r_count_11_io_out ? io_r_256_b : _GEN_3645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3647 = 9'h101 == r_count_11_io_out ? io_r_257_b : _GEN_3646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3648 = 9'h102 == r_count_11_io_out ? io_r_258_b : _GEN_3647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3649 = 9'h103 == r_count_11_io_out ? io_r_259_b : _GEN_3648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3650 = 9'h104 == r_count_11_io_out ? io_r_260_b : _GEN_3649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3651 = 9'h105 == r_count_11_io_out ? io_r_261_b : _GEN_3650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3652 = 9'h106 == r_count_11_io_out ? io_r_262_b : _GEN_3651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3653 = 9'h107 == r_count_11_io_out ? io_r_263_b : _GEN_3652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3654 = 9'h108 == r_count_11_io_out ? io_r_264_b : _GEN_3653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3655 = 9'h109 == r_count_11_io_out ? io_r_265_b : _GEN_3654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3656 = 9'h10a == r_count_11_io_out ? io_r_266_b : _GEN_3655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3657 = 9'h10b == r_count_11_io_out ? io_r_267_b : _GEN_3656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3658 = 9'h10c == r_count_11_io_out ? io_r_268_b : _GEN_3657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3659 = 9'h10d == r_count_11_io_out ? io_r_269_b : _GEN_3658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3660 = 9'h10e == r_count_11_io_out ? io_r_270_b : _GEN_3659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3661 = 9'h10f == r_count_11_io_out ? io_r_271_b : _GEN_3660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3662 = 9'h110 == r_count_11_io_out ? io_r_272_b : _GEN_3661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3663 = 9'h111 == r_count_11_io_out ? io_r_273_b : _GEN_3662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3664 = 9'h112 == r_count_11_io_out ? io_r_274_b : _GEN_3663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3665 = 9'h113 == r_count_11_io_out ? io_r_275_b : _GEN_3664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3666 = 9'h114 == r_count_11_io_out ? io_r_276_b : _GEN_3665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3667 = 9'h115 == r_count_11_io_out ? io_r_277_b : _GEN_3666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3668 = 9'h116 == r_count_11_io_out ? io_r_278_b : _GEN_3667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3669 = 9'h117 == r_count_11_io_out ? io_r_279_b : _GEN_3668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3670 = 9'h118 == r_count_11_io_out ? io_r_280_b : _GEN_3669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3671 = 9'h119 == r_count_11_io_out ? io_r_281_b : _GEN_3670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3672 = 9'h11a == r_count_11_io_out ? io_r_282_b : _GEN_3671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3673 = 9'h11b == r_count_11_io_out ? io_r_283_b : _GEN_3672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3674 = 9'h11c == r_count_11_io_out ? io_r_284_b : _GEN_3673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3675 = 9'h11d == r_count_11_io_out ? io_r_285_b : _GEN_3674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3676 = 9'h11e == r_count_11_io_out ? io_r_286_b : _GEN_3675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3677 = 9'h11f == r_count_11_io_out ? io_r_287_b : _GEN_3676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3678 = 9'h120 == r_count_11_io_out ? io_r_288_b : _GEN_3677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3679 = 9'h121 == r_count_11_io_out ? io_r_289_b : _GEN_3678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3680 = 9'h122 == r_count_11_io_out ? io_r_290_b : _GEN_3679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3681 = 9'h123 == r_count_11_io_out ? io_r_291_b : _GEN_3680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3682 = 9'h124 == r_count_11_io_out ? io_r_292_b : _GEN_3681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3683 = 9'h125 == r_count_11_io_out ? io_r_293_b : _GEN_3682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3684 = 9'h126 == r_count_11_io_out ? io_r_294_b : _GEN_3683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3685 = 9'h127 == r_count_11_io_out ? io_r_295_b : _GEN_3684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3686 = 9'h128 == r_count_11_io_out ? io_r_296_b : _GEN_3685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3687 = 9'h129 == r_count_11_io_out ? io_r_297_b : _GEN_3686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3688 = 9'h12a == r_count_11_io_out ? io_r_298_b : _GEN_3687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3691 = 9'h1 == r_count_12_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3692 = 9'h2 == r_count_12_io_out ? io_r_2_b : _GEN_3691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3693 = 9'h3 == r_count_12_io_out ? io_r_3_b : _GEN_3692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3694 = 9'h4 == r_count_12_io_out ? io_r_4_b : _GEN_3693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3695 = 9'h5 == r_count_12_io_out ? io_r_5_b : _GEN_3694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3696 = 9'h6 == r_count_12_io_out ? io_r_6_b : _GEN_3695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3697 = 9'h7 == r_count_12_io_out ? io_r_7_b : _GEN_3696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3698 = 9'h8 == r_count_12_io_out ? io_r_8_b : _GEN_3697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3699 = 9'h9 == r_count_12_io_out ? io_r_9_b : _GEN_3698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3700 = 9'ha == r_count_12_io_out ? io_r_10_b : _GEN_3699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3701 = 9'hb == r_count_12_io_out ? io_r_11_b : _GEN_3700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3702 = 9'hc == r_count_12_io_out ? io_r_12_b : _GEN_3701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3703 = 9'hd == r_count_12_io_out ? io_r_13_b : _GEN_3702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3704 = 9'he == r_count_12_io_out ? io_r_14_b : _GEN_3703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3705 = 9'hf == r_count_12_io_out ? io_r_15_b : _GEN_3704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3706 = 9'h10 == r_count_12_io_out ? io_r_16_b : _GEN_3705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3707 = 9'h11 == r_count_12_io_out ? io_r_17_b : _GEN_3706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3708 = 9'h12 == r_count_12_io_out ? io_r_18_b : _GEN_3707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3709 = 9'h13 == r_count_12_io_out ? io_r_19_b : _GEN_3708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3710 = 9'h14 == r_count_12_io_out ? io_r_20_b : _GEN_3709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3711 = 9'h15 == r_count_12_io_out ? io_r_21_b : _GEN_3710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3712 = 9'h16 == r_count_12_io_out ? io_r_22_b : _GEN_3711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3713 = 9'h17 == r_count_12_io_out ? io_r_23_b : _GEN_3712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3714 = 9'h18 == r_count_12_io_out ? io_r_24_b : _GEN_3713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3715 = 9'h19 == r_count_12_io_out ? io_r_25_b : _GEN_3714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3716 = 9'h1a == r_count_12_io_out ? io_r_26_b : _GEN_3715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3717 = 9'h1b == r_count_12_io_out ? io_r_27_b : _GEN_3716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3718 = 9'h1c == r_count_12_io_out ? io_r_28_b : _GEN_3717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3719 = 9'h1d == r_count_12_io_out ? io_r_29_b : _GEN_3718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3720 = 9'h1e == r_count_12_io_out ? io_r_30_b : _GEN_3719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3721 = 9'h1f == r_count_12_io_out ? io_r_31_b : _GEN_3720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3722 = 9'h20 == r_count_12_io_out ? io_r_32_b : _GEN_3721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3723 = 9'h21 == r_count_12_io_out ? io_r_33_b : _GEN_3722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3724 = 9'h22 == r_count_12_io_out ? io_r_34_b : _GEN_3723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3725 = 9'h23 == r_count_12_io_out ? io_r_35_b : _GEN_3724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3726 = 9'h24 == r_count_12_io_out ? io_r_36_b : _GEN_3725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3727 = 9'h25 == r_count_12_io_out ? io_r_37_b : _GEN_3726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3728 = 9'h26 == r_count_12_io_out ? io_r_38_b : _GEN_3727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3729 = 9'h27 == r_count_12_io_out ? io_r_39_b : _GEN_3728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3730 = 9'h28 == r_count_12_io_out ? io_r_40_b : _GEN_3729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3731 = 9'h29 == r_count_12_io_out ? io_r_41_b : _GEN_3730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3732 = 9'h2a == r_count_12_io_out ? io_r_42_b : _GEN_3731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3733 = 9'h2b == r_count_12_io_out ? io_r_43_b : _GEN_3732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3734 = 9'h2c == r_count_12_io_out ? io_r_44_b : _GEN_3733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3735 = 9'h2d == r_count_12_io_out ? io_r_45_b : _GEN_3734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3736 = 9'h2e == r_count_12_io_out ? io_r_46_b : _GEN_3735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3737 = 9'h2f == r_count_12_io_out ? io_r_47_b : _GEN_3736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3738 = 9'h30 == r_count_12_io_out ? io_r_48_b : _GEN_3737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3739 = 9'h31 == r_count_12_io_out ? io_r_49_b : _GEN_3738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3740 = 9'h32 == r_count_12_io_out ? io_r_50_b : _GEN_3739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3741 = 9'h33 == r_count_12_io_out ? io_r_51_b : _GEN_3740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3742 = 9'h34 == r_count_12_io_out ? io_r_52_b : _GEN_3741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3743 = 9'h35 == r_count_12_io_out ? io_r_53_b : _GEN_3742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3744 = 9'h36 == r_count_12_io_out ? io_r_54_b : _GEN_3743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3745 = 9'h37 == r_count_12_io_out ? io_r_55_b : _GEN_3744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3746 = 9'h38 == r_count_12_io_out ? io_r_56_b : _GEN_3745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3747 = 9'h39 == r_count_12_io_out ? io_r_57_b : _GEN_3746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3748 = 9'h3a == r_count_12_io_out ? io_r_58_b : _GEN_3747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3749 = 9'h3b == r_count_12_io_out ? io_r_59_b : _GEN_3748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3750 = 9'h3c == r_count_12_io_out ? io_r_60_b : _GEN_3749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3751 = 9'h3d == r_count_12_io_out ? io_r_61_b : _GEN_3750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3752 = 9'h3e == r_count_12_io_out ? io_r_62_b : _GEN_3751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3753 = 9'h3f == r_count_12_io_out ? io_r_63_b : _GEN_3752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3754 = 9'h40 == r_count_12_io_out ? io_r_64_b : _GEN_3753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3755 = 9'h41 == r_count_12_io_out ? io_r_65_b : _GEN_3754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3756 = 9'h42 == r_count_12_io_out ? io_r_66_b : _GEN_3755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3757 = 9'h43 == r_count_12_io_out ? io_r_67_b : _GEN_3756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3758 = 9'h44 == r_count_12_io_out ? io_r_68_b : _GEN_3757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3759 = 9'h45 == r_count_12_io_out ? io_r_69_b : _GEN_3758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3760 = 9'h46 == r_count_12_io_out ? io_r_70_b : _GEN_3759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3761 = 9'h47 == r_count_12_io_out ? io_r_71_b : _GEN_3760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3762 = 9'h48 == r_count_12_io_out ? io_r_72_b : _GEN_3761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3763 = 9'h49 == r_count_12_io_out ? io_r_73_b : _GEN_3762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3764 = 9'h4a == r_count_12_io_out ? io_r_74_b : _GEN_3763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3765 = 9'h4b == r_count_12_io_out ? io_r_75_b : _GEN_3764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3766 = 9'h4c == r_count_12_io_out ? io_r_76_b : _GEN_3765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3767 = 9'h4d == r_count_12_io_out ? io_r_77_b : _GEN_3766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3768 = 9'h4e == r_count_12_io_out ? io_r_78_b : _GEN_3767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3769 = 9'h4f == r_count_12_io_out ? io_r_79_b : _GEN_3768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3770 = 9'h50 == r_count_12_io_out ? io_r_80_b : _GEN_3769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3771 = 9'h51 == r_count_12_io_out ? io_r_81_b : _GEN_3770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3772 = 9'h52 == r_count_12_io_out ? io_r_82_b : _GEN_3771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3773 = 9'h53 == r_count_12_io_out ? io_r_83_b : _GEN_3772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3774 = 9'h54 == r_count_12_io_out ? io_r_84_b : _GEN_3773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3775 = 9'h55 == r_count_12_io_out ? io_r_85_b : _GEN_3774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3776 = 9'h56 == r_count_12_io_out ? io_r_86_b : _GEN_3775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3777 = 9'h57 == r_count_12_io_out ? io_r_87_b : _GEN_3776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3778 = 9'h58 == r_count_12_io_out ? io_r_88_b : _GEN_3777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3779 = 9'h59 == r_count_12_io_out ? io_r_89_b : _GEN_3778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3780 = 9'h5a == r_count_12_io_out ? io_r_90_b : _GEN_3779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3781 = 9'h5b == r_count_12_io_out ? io_r_91_b : _GEN_3780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3782 = 9'h5c == r_count_12_io_out ? io_r_92_b : _GEN_3781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3783 = 9'h5d == r_count_12_io_out ? io_r_93_b : _GEN_3782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3784 = 9'h5e == r_count_12_io_out ? io_r_94_b : _GEN_3783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3785 = 9'h5f == r_count_12_io_out ? io_r_95_b : _GEN_3784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3786 = 9'h60 == r_count_12_io_out ? io_r_96_b : _GEN_3785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3787 = 9'h61 == r_count_12_io_out ? io_r_97_b : _GEN_3786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3788 = 9'h62 == r_count_12_io_out ? io_r_98_b : _GEN_3787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3789 = 9'h63 == r_count_12_io_out ? io_r_99_b : _GEN_3788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3790 = 9'h64 == r_count_12_io_out ? io_r_100_b : _GEN_3789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3791 = 9'h65 == r_count_12_io_out ? io_r_101_b : _GEN_3790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3792 = 9'h66 == r_count_12_io_out ? io_r_102_b : _GEN_3791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3793 = 9'h67 == r_count_12_io_out ? io_r_103_b : _GEN_3792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3794 = 9'h68 == r_count_12_io_out ? io_r_104_b : _GEN_3793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3795 = 9'h69 == r_count_12_io_out ? io_r_105_b : _GEN_3794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3796 = 9'h6a == r_count_12_io_out ? io_r_106_b : _GEN_3795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3797 = 9'h6b == r_count_12_io_out ? io_r_107_b : _GEN_3796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3798 = 9'h6c == r_count_12_io_out ? io_r_108_b : _GEN_3797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3799 = 9'h6d == r_count_12_io_out ? io_r_109_b : _GEN_3798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3800 = 9'h6e == r_count_12_io_out ? io_r_110_b : _GEN_3799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3801 = 9'h6f == r_count_12_io_out ? io_r_111_b : _GEN_3800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3802 = 9'h70 == r_count_12_io_out ? io_r_112_b : _GEN_3801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3803 = 9'h71 == r_count_12_io_out ? io_r_113_b : _GEN_3802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3804 = 9'h72 == r_count_12_io_out ? io_r_114_b : _GEN_3803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3805 = 9'h73 == r_count_12_io_out ? io_r_115_b : _GEN_3804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3806 = 9'h74 == r_count_12_io_out ? io_r_116_b : _GEN_3805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3807 = 9'h75 == r_count_12_io_out ? io_r_117_b : _GEN_3806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3808 = 9'h76 == r_count_12_io_out ? io_r_118_b : _GEN_3807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3809 = 9'h77 == r_count_12_io_out ? io_r_119_b : _GEN_3808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3810 = 9'h78 == r_count_12_io_out ? io_r_120_b : _GEN_3809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3811 = 9'h79 == r_count_12_io_out ? io_r_121_b : _GEN_3810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3812 = 9'h7a == r_count_12_io_out ? io_r_122_b : _GEN_3811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3813 = 9'h7b == r_count_12_io_out ? io_r_123_b : _GEN_3812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3814 = 9'h7c == r_count_12_io_out ? io_r_124_b : _GEN_3813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3815 = 9'h7d == r_count_12_io_out ? io_r_125_b : _GEN_3814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3816 = 9'h7e == r_count_12_io_out ? io_r_126_b : _GEN_3815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3817 = 9'h7f == r_count_12_io_out ? io_r_127_b : _GEN_3816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3818 = 9'h80 == r_count_12_io_out ? io_r_128_b : _GEN_3817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3819 = 9'h81 == r_count_12_io_out ? io_r_129_b : _GEN_3818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3820 = 9'h82 == r_count_12_io_out ? io_r_130_b : _GEN_3819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3821 = 9'h83 == r_count_12_io_out ? io_r_131_b : _GEN_3820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3822 = 9'h84 == r_count_12_io_out ? io_r_132_b : _GEN_3821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3823 = 9'h85 == r_count_12_io_out ? io_r_133_b : _GEN_3822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3824 = 9'h86 == r_count_12_io_out ? io_r_134_b : _GEN_3823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3825 = 9'h87 == r_count_12_io_out ? io_r_135_b : _GEN_3824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3826 = 9'h88 == r_count_12_io_out ? io_r_136_b : _GEN_3825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3827 = 9'h89 == r_count_12_io_out ? io_r_137_b : _GEN_3826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3828 = 9'h8a == r_count_12_io_out ? io_r_138_b : _GEN_3827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3829 = 9'h8b == r_count_12_io_out ? io_r_139_b : _GEN_3828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3830 = 9'h8c == r_count_12_io_out ? io_r_140_b : _GEN_3829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3831 = 9'h8d == r_count_12_io_out ? io_r_141_b : _GEN_3830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3832 = 9'h8e == r_count_12_io_out ? io_r_142_b : _GEN_3831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3833 = 9'h8f == r_count_12_io_out ? io_r_143_b : _GEN_3832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3834 = 9'h90 == r_count_12_io_out ? io_r_144_b : _GEN_3833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3835 = 9'h91 == r_count_12_io_out ? io_r_145_b : _GEN_3834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3836 = 9'h92 == r_count_12_io_out ? io_r_146_b : _GEN_3835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3837 = 9'h93 == r_count_12_io_out ? io_r_147_b : _GEN_3836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3838 = 9'h94 == r_count_12_io_out ? io_r_148_b : _GEN_3837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3839 = 9'h95 == r_count_12_io_out ? io_r_149_b : _GEN_3838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3840 = 9'h96 == r_count_12_io_out ? io_r_150_b : _GEN_3839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3841 = 9'h97 == r_count_12_io_out ? io_r_151_b : _GEN_3840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3842 = 9'h98 == r_count_12_io_out ? io_r_152_b : _GEN_3841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3843 = 9'h99 == r_count_12_io_out ? io_r_153_b : _GEN_3842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3844 = 9'h9a == r_count_12_io_out ? io_r_154_b : _GEN_3843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3845 = 9'h9b == r_count_12_io_out ? io_r_155_b : _GEN_3844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3846 = 9'h9c == r_count_12_io_out ? io_r_156_b : _GEN_3845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3847 = 9'h9d == r_count_12_io_out ? io_r_157_b : _GEN_3846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3848 = 9'h9e == r_count_12_io_out ? io_r_158_b : _GEN_3847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3849 = 9'h9f == r_count_12_io_out ? io_r_159_b : _GEN_3848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3850 = 9'ha0 == r_count_12_io_out ? io_r_160_b : _GEN_3849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3851 = 9'ha1 == r_count_12_io_out ? io_r_161_b : _GEN_3850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3852 = 9'ha2 == r_count_12_io_out ? io_r_162_b : _GEN_3851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3853 = 9'ha3 == r_count_12_io_out ? io_r_163_b : _GEN_3852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3854 = 9'ha4 == r_count_12_io_out ? io_r_164_b : _GEN_3853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3855 = 9'ha5 == r_count_12_io_out ? io_r_165_b : _GEN_3854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3856 = 9'ha6 == r_count_12_io_out ? io_r_166_b : _GEN_3855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3857 = 9'ha7 == r_count_12_io_out ? io_r_167_b : _GEN_3856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3858 = 9'ha8 == r_count_12_io_out ? io_r_168_b : _GEN_3857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3859 = 9'ha9 == r_count_12_io_out ? io_r_169_b : _GEN_3858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3860 = 9'haa == r_count_12_io_out ? io_r_170_b : _GEN_3859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3861 = 9'hab == r_count_12_io_out ? io_r_171_b : _GEN_3860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3862 = 9'hac == r_count_12_io_out ? io_r_172_b : _GEN_3861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3863 = 9'had == r_count_12_io_out ? io_r_173_b : _GEN_3862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3864 = 9'hae == r_count_12_io_out ? io_r_174_b : _GEN_3863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3865 = 9'haf == r_count_12_io_out ? io_r_175_b : _GEN_3864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3866 = 9'hb0 == r_count_12_io_out ? io_r_176_b : _GEN_3865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3867 = 9'hb1 == r_count_12_io_out ? io_r_177_b : _GEN_3866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3868 = 9'hb2 == r_count_12_io_out ? io_r_178_b : _GEN_3867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3869 = 9'hb3 == r_count_12_io_out ? io_r_179_b : _GEN_3868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3870 = 9'hb4 == r_count_12_io_out ? io_r_180_b : _GEN_3869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3871 = 9'hb5 == r_count_12_io_out ? io_r_181_b : _GEN_3870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3872 = 9'hb6 == r_count_12_io_out ? io_r_182_b : _GEN_3871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3873 = 9'hb7 == r_count_12_io_out ? io_r_183_b : _GEN_3872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3874 = 9'hb8 == r_count_12_io_out ? io_r_184_b : _GEN_3873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3875 = 9'hb9 == r_count_12_io_out ? io_r_185_b : _GEN_3874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3876 = 9'hba == r_count_12_io_out ? io_r_186_b : _GEN_3875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3877 = 9'hbb == r_count_12_io_out ? io_r_187_b : _GEN_3876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3878 = 9'hbc == r_count_12_io_out ? io_r_188_b : _GEN_3877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3879 = 9'hbd == r_count_12_io_out ? io_r_189_b : _GEN_3878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3880 = 9'hbe == r_count_12_io_out ? io_r_190_b : _GEN_3879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3881 = 9'hbf == r_count_12_io_out ? io_r_191_b : _GEN_3880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3882 = 9'hc0 == r_count_12_io_out ? io_r_192_b : _GEN_3881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3883 = 9'hc1 == r_count_12_io_out ? io_r_193_b : _GEN_3882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3884 = 9'hc2 == r_count_12_io_out ? io_r_194_b : _GEN_3883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3885 = 9'hc3 == r_count_12_io_out ? io_r_195_b : _GEN_3884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3886 = 9'hc4 == r_count_12_io_out ? io_r_196_b : _GEN_3885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3887 = 9'hc5 == r_count_12_io_out ? io_r_197_b : _GEN_3886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3888 = 9'hc6 == r_count_12_io_out ? io_r_198_b : _GEN_3887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3889 = 9'hc7 == r_count_12_io_out ? io_r_199_b : _GEN_3888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3890 = 9'hc8 == r_count_12_io_out ? io_r_200_b : _GEN_3889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3891 = 9'hc9 == r_count_12_io_out ? io_r_201_b : _GEN_3890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3892 = 9'hca == r_count_12_io_out ? io_r_202_b : _GEN_3891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3893 = 9'hcb == r_count_12_io_out ? io_r_203_b : _GEN_3892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3894 = 9'hcc == r_count_12_io_out ? io_r_204_b : _GEN_3893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3895 = 9'hcd == r_count_12_io_out ? io_r_205_b : _GEN_3894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3896 = 9'hce == r_count_12_io_out ? io_r_206_b : _GEN_3895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3897 = 9'hcf == r_count_12_io_out ? io_r_207_b : _GEN_3896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3898 = 9'hd0 == r_count_12_io_out ? io_r_208_b : _GEN_3897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3899 = 9'hd1 == r_count_12_io_out ? io_r_209_b : _GEN_3898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3900 = 9'hd2 == r_count_12_io_out ? io_r_210_b : _GEN_3899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3901 = 9'hd3 == r_count_12_io_out ? io_r_211_b : _GEN_3900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3902 = 9'hd4 == r_count_12_io_out ? io_r_212_b : _GEN_3901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3903 = 9'hd5 == r_count_12_io_out ? io_r_213_b : _GEN_3902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3904 = 9'hd6 == r_count_12_io_out ? io_r_214_b : _GEN_3903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3905 = 9'hd7 == r_count_12_io_out ? io_r_215_b : _GEN_3904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3906 = 9'hd8 == r_count_12_io_out ? io_r_216_b : _GEN_3905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3907 = 9'hd9 == r_count_12_io_out ? io_r_217_b : _GEN_3906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3908 = 9'hda == r_count_12_io_out ? io_r_218_b : _GEN_3907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3909 = 9'hdb == r_count_12_io_out ? io_r_219_b : _GEN_3908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3910 = 9'hdc == r_count_12_io_out ? io_r_220_b : _GEN_3909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3911 = 9'hdd == r_count_12_io_out ? io_r_221_b : _GEN_3910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3912 = 9'hde == r_count_12_io_out ? io_r_222_b : _GEN_3911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3913 = 9'hdf == r_count_12_io_out ? io_r_223_b : _GEN_3912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3914 = 9'he0 == r_count_12_io_out ? io_r_224_b : _GEN_3913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3915 = 9'he1 == r_count_12_io_out ? io_r_225_b : _GEN_3914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3916 = 9'he2 == r_count_12_io_out ? io_r_226_b : _GEN_3915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3917 = 9'he3 == r_count_12_io_out ? io_r_227_b : _GEN_3916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3918 = 9'he4 == r_count_12_io_out ? io_r_228_b : _GEN_3917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3919 = 9'he5 == r_count_12_io_out ? io_r_229_b : _GEN_3918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3920 = 9'he6 == r_count_12_io_out ? io_r_230_b : _GEN_3919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3921 = 9'he7 == r_count_12_io_out ? io_r_231_b : _GEN_3920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3922 = 9'he8 == r_count_12_io_out ? io_r_232_b : _GEN_3921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3923 = 9'he9 == r_count_12_io_out ? io_r_233_b : _GEN_3922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3924 = 9'hea == r_count_12_io_out ? io_r_234_b : _GEN_3923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3925 = 9'heb == r_count_12_io_out ? io_r_235_b : _GEN_3924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3926 = 9'hec == r_count_12_io_out ? io_r_236_b : _GEN_3925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3927 = 9'hed == r_count_12_io_out ? io_r_237_b : _GEN_3926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3928 = 9'hee == r_count_12_io_out ? io_r_238_b : _GEN_3927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3929 = 9'hef == r_count_12_io_out ? io_r_239_b : _GEN_3928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3930 = 9'hf0 == r_count_12_io_out ? io_r_240_b : _GEN_3929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3931 = 9'hf1 == r_count_12_io_out ? io_r_241_b : _GEN_3930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3932 = 9'hf2 == r_count_12_io_out ? io_r_242_b : _GEN_3931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3933 = 9'hf3 == r_count_12_io_out ? io_r_243_b : _GEN_3932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3934 = 9'hf4 == r_count_12_io_out ? io_r_244_b : _GEN_3933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3935 = 9'hf5 == r_count_12_io_out ? io_r_245_b : _GEN_3934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3936 = 9'hf6 == r_count_12_io_out ? io_r_246_b : _GEN_3935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3937 = 9'hf7 == r_count_12_io_out ? io_r_247_b : _GEN_3936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3938 = 9'hf8 == r_count_12_io_out ? io_r_248_b : _GEN_3937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3939 = 9'hf9 == r_count_12_io_out ? io_r_249_b : _GEN_3938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3940 = 9'hfa == r_count_12_io_out ? io_r_250_b : _GEN_3939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3941 = 9'hfb == r_count_12_io_out ? io_r_251_b : _GEN_3940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3942 = 9'hfc == r_count_12_io_out ? io_r_252_b : _GEN_3941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3943 = 9'hfd == r_count_12_io_out ? io_r_253_b : _GEN_3942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3944 = 9'hfe == r_count_12_io_out ? io_r_254_b : _GEN_3943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3945 = 9'hff == r_count_12_io_out ? io_r_255_b : _GEN_3944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3946 = 9'h100 == r_count_12_io_out ? io_r_256_b : _GEN_3945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3947 = 9'h101 == r_count_12_io_out ? io_r_257_b : _GEN_3946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3948 = 9'h102 == r_count_12_io_out ? io_r_258_b : _GEN_3947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3949 = 9'h103 == r_count_12_io_out ? io_r_259_b : _GEN_3948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3950 = 9'h104 == r_count_12_io_out ? io_r_260_b : _GEN_3949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3951 = 9'h105 == r_count_12_io_out ? io_r_261_b : _GEN_3950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3952 = 9'h106 == r_count_12_io_out ? io_r_262_b : _GEN_3951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3953 = 9'h107 == r_count_12_io_out ? io_r_263_b : _GEN_3952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3954 = 9'h108 == r_count_12_io_out ? io_r_264_b : _GEN_3953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3955 = 9'h109 == r_count_12_io_out ? io_r_265_b : _GEN_3954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3956 = 9'h10a == r_count_12_io_out ? io_r_266_b : _GEN_3955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3957 = 9'h10b == r_count_12_io_out ? io_r_267_b : _GEN_3956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3958 = 9'h10c == r_count_12_io_out ? io_r_268_b : _GEN_3957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3959 = 9'h10d == r_count_12_io_out ? io_r_269_b : _GEN_3958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3960 = 9'h10e == r_count_12_io_out ? io_r_270_b : _GEN_3959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3961 = 9'h10f == r_count_12_io_out ? io_r_271_b : _GEN_3960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3962 = 9'h110 == r_count_12_io_out ? io_r_272_b : _GEN_3961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3963 = 9'h111 == r_count_12_io_out ? io_r_273_b : _GEN_3962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3964 = 9'h112 == r_count_12_io_out ? io_r_274_b : _GEN_3963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3965 = 9'h113 == r_count_12_io_out ? io_r_275_b : _GEN_3964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3966 = 9'h114 == r_count_12_io_out ? io_r_276_b : _GEN_3965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3967 = 9'h115 == r_count_12_io_out ? io_r_277_b : _GEN_3966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3968 = 9'h116 == r_count_12_io_out ? io_r_278_b : _GEN_3967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3969 = 9'h117 == r_count_12_io_out ? io_r_279_b : _GEN_3968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3970 = 9'h118 == r_count_12_io_out ? io_r_280_b : _GEN_3969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3971 = 9'h119 == r_count_12_io_out ? io_r_281_b : _GEN_3970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3972 = 9'h11a == r_count_12_io_out ? io_r_282_b : _GEN_3971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3973 = 9'h11b == r_count_12_io_out ? io_r_283_b : _GEN_3972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3974 = 9'h11c == r_count_12_io_out ? io_r_284_b : _GEN_3973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3975 = 9'h11d == r_count_12_io_out ? io_r_285_b : _GEN_3974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3976 = 9'h11e == r_count_12_io_out ? io_r_286_b : _GEN_3975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3977 = 9'h11f == r_count_12_io_out ? io_r_287_b : _GEN_3976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3978 = 9'h120 == r_count_12_io_out ? io_r_288_b : _GEN_3977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3979 = 9'h121 == r_count_12_io_out ? io_r_289_b : _GEN_3978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3980 = 9'h122 == r_count_12_io_out ? io_r_290_b : _GEN_3979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3981 = 9'h123 == r_count_12_io_out ? io_r_291_b : _GEN_3980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3982 = 9'h124 == r_count_12_io_out ? io_r_292_b : _GEN_3981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3983 = 9'h125 == r_count_12_io_out ? io_r_293_b : _GEN_3982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3984 = 9'h126 == r_count_12_io_out ? io_r_294_b : _GEN_3983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3985 = 9'h127 == r_count_12_io_out ? io_r_295_b : _GEN_3984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3986 = 9'h128 == r_count_12_io_out ? io_r_296_b : _GEN_3985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3987 = 9'h129 == r_count_12_io_out ? io_r_297_b : _GEN_3986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3988 = 9'h12a == r_count_12_io_out ? io_r_298_b : _GEN_3987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3991 = 9'h1 == r_count_13_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3992 = 9'h2 == r_count_13_io_out ? io_r_2_b : _GEN_3991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3993 = 9'h3 == r_count_13_io_out ? io_r_3_b : _GEN_3992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3994 = 9'h4 == r_count_13_io_out ? io_r_4_b : _GEN_3993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3995 = 9'h5 == r_count_13_io_out ? io_r_5_b : _GEN_3994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3996 = 9'h6 == r_count_13_io_out ? io_r_6_b : _GEN_3995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3997 = 9'h7 == r_count_13_io_out ? io_r_7_b : _GEN_3996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3998 = 9'h8 == r_count_13_io_out ? io_r_8_b : _GEN_3997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3999 = 9'h9 == r_count_13_io_out ? io_r_9_b : _GEN_3998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4000 = 9'ha == r_count_13_io_out ? io_r_10_b : _GEN_3999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4001 = 9'hb == r_count_13_io_out ? io_r_11_b : _GEN_4000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4002 = 9'hc == r_count_13_io_out ? io_r_12_b : _GEN_4001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4003 = 9'hd == r_count_13_io_out ? io_r_13_b : _GEN_4002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4004 = 9'he == r_count_13_io_out ? io_r_14_b : _GEN_4003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4005 = 9'hf == r_count_13_io_out ? io_r_15_b : _GEN_4004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4006 = 9'h10 == r_count_13_io_out ? io_r_16_b : _GEN_4005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4007 = 9'h11 == r_count_13_io_out ? io_r_17_b : _GEN_4006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4008 = 9'h12 == r_count_13_io_out ? io_r_18_b : _GEN_4007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4009 = 9'h13 == r_count_13_io_out ? io_r_19_b : _GEN_4008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4010 = 9'h14 == r_count_13_io_out ? io_r_20_b : _GEN_4009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4011 = 9'h15 == r_count_13_io_out ? io_r_21_b : _GEN_4010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4012 = 9'h16 == r_count_13_io_out ? io_r_22_b : _GEN_4011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4013 = 9'h17 == r_count_13_io_out ? io_r_23_b : _GEN_4012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4014 = 9'h18 == r_count_13_io_out ? io_r_24_b : _GEN_4013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4015 = 9'h19 == r_count_13_io_out ? io_r_25_b : _GEN_4014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4016 = 9'h1a == r_count_13_io_out ? io_r_26_b : _GEN_4015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4017 = 9'h1b == r_count_13_io_out ? io_r_27_b : _GEN_4016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4018 = 9'h1c == r_count_13_io_out ? io_r_28_b : _GEN_4017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4019 = 9'h1d == r_count_13_io_out ? io_r_29_b : _GEN_4018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4020 = 9'h1e == r_count_13_io_out ? io_r_30_b : _GEN_4019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4021 = 9'h1f == r_count_13_io_out ? io_r_31_b : _GEN_4020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4022 = 9'h20 == r_count_13_io_out ? io_r_32_b : _GEN_4021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4023 = 9'h21 == r_count_13_io_out ? io_r_33_b : _GEN_4022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4024 = 9'h22 == r_count_13_io_out ? io_r_34_b : _GEN_4023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4025 = 9'h23 == r_count_13_io_out ? io_r_35_b : _GEN_4024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4026 = 9'h24 == r_count_13_io_out ? io_r_36_b : _GEN_4025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4027 = 9'h25 == r_count_13_io_out ? io_r_37_b : _GEN_4026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4028 = 9'h26 == r_count_13_io_out ? io_r_38_b : _GEN_4027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4029 = 9'h27 == r_count_13_io_out ? io_r_39_b : _GEN_4028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4030 = 9'h28 == r_count_13_io_out ? io_r_40_b : _GEN_4029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4031 = 9'h29 == r_count_13_io_out ? io_r_41_b : _GEN_4030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4032 = 9'h2a == r_count_13_io_out ? io_r_42_b : _GEN_4031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4033 = 9'h2b == r_count_13_io_out ? io_r_43_b : _GEN_4032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4034 = 9'h2c == r_count_13_io_out ? io_r_44_b : _GEN_4033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4035 = 9'h2d == r_count_13_io_out ? io_r_45_b : _GEN_4034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4036 = 9'h2e == r_count_13_io_out ? io_r_46_b : _GEN_4035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4037 = 9'h2f == r_count_13_io_out ? io_r_47_b : _GEN_4036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4038 = 9'h30 == r_count_13_io_out ? io_r_48_b : _GEN_4037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4039 = 9'h31 == r_count_13_io_out ? io_r_49_b : _GEN_4038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4040 = 9'h32 == r_count_13_io_out ? io_r_50_b : _GEN_4039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4041 = 9'h33 == r_count_13_io_out ? io_r_51_b : _GEN_4040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4042 = 9'h34 == r_count_13_io_out ? io_r_52_b : _GEN_4041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4043 = 9'h35 == r_count_13_io_out ? io_r_53_b : _GEN_4042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4044 = 9'h36 == r_count_13_io_out ? io_r_54_b : _GEN_4043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4045 = 9'h37 == r_count_13_io_out ? io_r_55_b : _GEN_4044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4046 = 9'h38 == r_count_13_io_out ? io_r_56_b : _GEN_4045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4047 = 9'h39 == r_count_13_io_out ? io_r_57_b : _GEN_4046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4048 = 9'h3a == r_count_13_io_out ? io_r_58_b : _GEN_4047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4049 = 9'h3b == r_count_13_io_out ? io_r_59_b : _GEN_4048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4050 = 9'h3c == r_count_13_io_out ? io_r_60_b : _GEN_4049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4051 = 9'h3d == r_count_13_io_out ? io_r_61_b : _GEN_4050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4052 = 9'h3e == r_count_13_io_out ? io_r_62_b : _GEN_4051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4053 = 9'h3f == r_count_13_io_out ? io_r_63_b : _GEN_4052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4054 = 9'h40 == r_count_13_io_out ? io_r_64_b : _GEN_4053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4055 = 9'h41 == r_count_13_io_out ? io_r_65_b : _GEN_4054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4056 = 9'h42 == r_count_13_io_out ? io_r_66_b : _GEN_4055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4057 = 9'h43 == r_count_13_io_out ? io_r_67_b : _GEN_4056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4058 = 9'h44 == r_count_13_io_out ? io_r_68_b : _GEN_4057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4059 = 9'h45 == r_count_13_io_out ? io_r_69_b : _GEN_4058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4060 = 9'h46 == r_count_13_io_out ? io_r_70_b : _GEN_4059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4061 = 9'h47 == r_count_13_io_out ? io_r_71_b : _GEN_4060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4062 = 9'h48 == r_count_13_io_out ? io_r_72_b : _GEN_4061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4063 = 9'h49 == r_count_13_io_out ? io_r_73_b : _GEN_4062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4064 = 9'h4a == r_count_13_io_out ? io_r_74_b : _GEN_4063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4065 = 9'h4b == r_count_13_io_out ? io_r_75_b : _GEN_4064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4066 = 9'h4c == r_count_13_io_out ? io_r_76_b : _GEN_4065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4067 = 9'h4d == r_count_13_io_out ? io_r_77_b : _GEN_4066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4068 = 9'h4e == r_count_13_io_out ? io_r_78_b : _GEN_4067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4069 = 9'h4f == r_count_13_io_out ? io_r_79_b : _GEN_4068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4070 = 9'h50 == r_count_13_io_out ? io_r_80_b : _GEN_4069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4071 = 9'h51 == r_count_13_io_out ? io_r_81_b : _GEN_4070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4072 = 9'h52 == r_count_13_io_out ? io_r_82_b : _GEN_4071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4073 = 9'h53 == r_count_13_io_out ? io_r_83_b : _GEN_4072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4074 = 9'h54 == r_count_13_io_out ? io_r_84_b : _GEN_4073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4075 = 9'h55 == r_count_13_io_out ? io_r_85_b : _GEN_4074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4076 = 9'h56 == r_count_13_io_out ? io_r_86_b : _GEN_4075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4077 = 9'h57 == r_count_13_io_out ? io_r_87_b : _GEN_4076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4078 = 9'h58 == r_count_13_io_out ? io_r_88_b : _GEN_4077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4079 = 9'h59 == r_count_13_io_out ? io_r_89_b : _GEN_4078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4080 = 9'h5a == r_count_13_io_out ? io_r_90_b : _GEN_4079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4081 = 9'h5b == r_count_13_io_out ? io_r_91_b : _GEN_4080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4082 = 9'h5c == r_count_13_io_out ? io_r_92_b : _GEN_4081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4083 = 9'h5d == r_count_13_io_out ? io_r_93_b : _GEN_4082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4084 = 9'h5e == r_count_13_io_out ? io_r_94_b : _GEN_4083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4085 = 9'h5f == r_count_13_io_out ? io_r_95_b : _GEN_4084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4086 = 9'h60 == r_count_13_io_out ? io_r_96_b : _GEN_4085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4087 = 9'h61 == r_count_13_io_out ? io_r_97_b : _GEN_4086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4088 = 9'h62 == r_count_13_io_out ? io_r_98_b : _GEN_4087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4089 = 9'h63 == r_count_13_io_out ? io_r_99_b : _GEN_4088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4090 = 9'h64 == r_count_13_io_out ? io_r_100_b : _GEN_4089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4091 = 9'h65 == r_count_13_io_out ? io_r_101_b : _GEN_4090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4092 = 9'h66 == r_count_13_io_out ? io_r_102_b : _GEN_4091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4093 = 9'h67 == r_count_13_io_out ? io_r_103_b : _GEN_4092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4094 = 9'h68 == r_count_13_io_out ? io_r_104_b : _GEN_4093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4095 = 9'h69 == r_count_13_io_out ? io_r_105_b : _GEN_4094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4096 = 9'h6a == r_count_13_io_out ? io_r_106_b : _GEN_4095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4097 = 9'h6b == r_count_13_io_out ? io_r_107_b : _GEN_4096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4098 = 9'h6c == r_count_13_io_out ? io_r_108_b : _GEN_4097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4099 = 9'h6d == r_count_13_io_out ? io_r_109_b : _GEN_4098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4100 = 9'h6e == r_count_13_io_out ? io_r_110_b : _GEN_4099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4101 = 9'h6f == r_count_13_io_out ? io_r_111_b : _GEN_4100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4102 = 9'h70 == r_count_13_io_out ? io_r_112_b : _GEN_4101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4103 = 9'h71 == r_count_13_io_out ? io_r_113_b : _GEN_4102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4104 = 9'h72 == r_count_13_io_out ? io_r_114_b : _GEN_4103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4105 = 9'h73 == r_count_13_io_out ? io_r_115_b : _GEN_4104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4106 = 9'h74 == r_count_13_io_out ? io_r_116_b : _GEN_4105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4107 = 9'h75 == r_count_13_io_out ? io_r_117_b : _GEN_4106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4108 = 9'h76 == r_count_13_io_out ? io_r_118_b : _GEN_4107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4109 = 9'h77 == r_count_13_io_out ? io_r_119_b : _GEN_4108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4110 = 9'h78 == r_count_13_io_out ? io_r_120_b : _GEN_4109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4111 = 9'h79 == r_count_13_io_out ? io_r_121_b : _GEN_4110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4112 = 9'h7a == r_count_13_io_out ? io_r_122_b : _GEN_4111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4113 = 9'h7b == r_count_13_io_out ? io_r_123_b : _GEN_4112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4114 = 9'h7c == r_count_13_io_out ? io_r_124_b : _GEN_4113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4115 = 9'h7d == r_count_13_io_out ? io_r_125_b : _GEN_4114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4116 = 9'h7e == r_count_13_io_out ? io_r_126_b : _GEN_4115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4117 = 9'h7f == r_count_13_io_out ? io_r_127_b : _GEN_4116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4118 = 9'h80 == r_count_13_io_out ? io_r_128_b : _GEN_4117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4119 = 9'h81 == r_count_13_io_out ? io_r_129_b : _GEN_4118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4120 = 9'h82 == r_count_13_io_out ? io_r_130_b : _GEN_4119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4121 = 9'h83 == r_count_13_io_out ? io_r_131_b : _GEN_4120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4122 = 9'h84 == r_count_13_io_out ? io_r_132_b : _GEN_4121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4123 = 9'h85 == r_count_13_io_out ? io_r_133_b : _GEN_4122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4124 = 9'h86 == r_count_13_io_out ? io_r_134_b : _GEN_4123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4125 = 9'h87 == r_count_13_io_out ? io_r_135_b : _GEN_4124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4126 = 9'h88 == r_count_13_io_out ? io_r_136_b : _GEN_4125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4127 = 9'h89 == r_count_13_io_out ? io_r_137_b : _GEN_4126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4128 = 9'h8a == r_count_13_io_out ? io_r_138_b : _GEN_4127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4129 = 9'h8b == r_count_13_io_out ? io_r_139_b : _GEN_4128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4130 = 9'h8c == r_count_13_io_out ? io_r_140_b : _GEN_4129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4131 = 9'h8d == r_count_13_io_out ? io_r_141_b : _GEN_4130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4132 = 9'h8e == r_count_13_io_out ? io_r_142_b : _GEN_4131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4133 = 9'h8f == r_count_13_io_out ? io_r_143_b : _GEN_4132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4134 = 9'h90 == r_count_13_io_out ? io_r_144_b : _GEN_4133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4135 = 9'h91 == r_count_13_io_out ? io_r_145_b : _GEN_4134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4136 = 9'h92 == r_count_13_io_out ? io_r_146_b : _GEN_4135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4137 = 9'h93 == r_count_13_io_out ? io_r_147_b : _GEN_4136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4138 = 9'h94 == r_count_13_io_out ? io_r_148_b : _GEN_4137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4139 = 9'h95 == r_count_13_io_out ? io_r_149_b : _GEN_4138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4140 = 9'h96 == r_count_13_io_out ? io_r_150_b : _GEN_4139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4141 = 9'h97 == r_count_13_io_out ? io_r_151_b : _GEN_4140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4142 = 9'h98 == r_count_13_io_out ? io_r_152_b : _GEN_4141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4143 = 9'h99 == r_count_13_io_out ? io_r_153_b : _GEN_4142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4144 = 9'h9a == r_count_13_io_out ? io_r_154_b : _GEN_4143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4145 = 9'h9b == r_count_13_io_out ? io_r_155_b : _GEN_4144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4146 = 9'h9c == r_count_13_io_out ? io_r_156_b : _GEN_4145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4147 = 9'h9d == r_count_13_io_out ? io_r_157_b : _GEN_4146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4148 = 9'h9e == r_count_13_io_out ? io_r_158_b : _GEN_4147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4149 = 9'h9f == r_count_13_io_out ? io_r_159_b : _GEN_4148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4150 = 9'ha0 == r_count_13_io_out ? io_r_160_b : _GEN_4149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4151 = 9'ha1 == r_count_13_io_out ? io_r_161_b : _GEN_4150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4152 = 9'ha2 == r_count_13_io_out ? io_r_162_b : _GEN_4151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4153 = 9'ha3 == r_count_13_io_out ? io_r_163_b : _GEN_4152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4154 = 9'ha4 == r_count_13_io_out ? io_r_164_b : _GEN_4153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4155 = 9'ha5 == r_count_13_io_out ? io_r_165_b : _GEN_4154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4156 = 9'ha6 == r_count_13_io_out ? io_r_166_b : _GEN_4155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4157 = 9'ha7 == r_count_13_io_out ? io_r_167_b : _GEN_4156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4158 = 9'ha8 == r_count_13_io_out ? io_r_168_b : _GEN_4157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4159 = 9'ha9 == r_count_13_io_out ? io_r_169_b : _GEN_4158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4160 = 9'haa == r_count_13_io_out ? io_r_170_b : _GEN_4159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4161 = 9'hab == r_count_13_io_out ? io_r_171_b : _GEN_4160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4162 = 9'hac == r_count_13_io_out ? io_r_172_b : _GEN_4161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4163 = 9'had == r_count_13_io_out ? io_r_173_b : _GEN_4162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4164 = 9'hae == r_count_13_io_out ? io_r_174_b : _GEN_4163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4165 = 9'haf == r_count_13_io_out ? io_r_175_b : _GEN_4164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4166 = 9'hb0 == r_count_13_io_out ? io_r_176_b : _GEN_4165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4167 = 9'hb1 == r_count_13_io_out ? io_r_177_b : _GEN_4166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4168 = 9'hb2 == r_count_13_io_out ? io_r_178_b : _GEN_4167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4169 = 9'hb3 == r_count_13_io_out ? io_r_179_b : _GEN_4168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4170 = 9'hb4 == r_count_13_io_out ? io_r_180_b : _GEN_4169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4171 = 9'hb5 == r_count_13_io_out ? io_r_181_b : _GEN_4170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4172 = 9'hb6 == r_count_13_io_out ? io_r_182_b : _GEN_4171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4173 = 9'hb7 == r_count_13_io_out ? io_r_183_b : _GEN_4172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4174 = 9'hb8 == r_count_13_io_out ? io_r_184_b : _GEN_4173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4175 = 9'hb9 == r_count_13_io_out ? io_r_185_b : _GEN_4174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4176 = 9'hba == r_count_13_io_out ? io_r_186_b : _GEN_4175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4177 = 9'hbb == r_count_13_io_out ? io_r_187_b : _GEN_4176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4178 = 9'hbc == r_count_13_io_out ? io_r_188_b : _GEN_4177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4179 = 9'hbd == r_count_13_io_out ? io_r_189_b : _GEN_4178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4180 = 9'hbe == r_count_13_io_out ? io_r_190_b : _GEN_4179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4181 = 9'hbf == r_count_13_io_out ? io_r_191_b : _GEN_4180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4182 = 9'hc0 == r_count_13_io_out ? io_r_192_b : _GEN_4181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4183 = 9'hc1 == r_count_13_io_out ? io_r_193_b : _GEN_4182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4184 = 9'hc2 == r_count_13_io_out ? io_r_194_b : _GEN_4183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4185 = 9'hc3 == r_count_13_io_out ? io_r_195_b : _GEN_4184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4186 = 9'hc4 == r_count_13_io_out ? io_r_196_b : _GEN_4185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4187 = 9'hc5 == r_count_13_io_out ? io_r_197_b : _GEN_4186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4188 = 9'hc6 == r_count_13_io_out ? io_r_198_b : _GEN_4187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4189 = 9'hc7 == r_count_13_io_out ? io_r_199_b : _GEN_4188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4190 = 9'hc8 == r_count_13_io_out ? io_r_200_b : _GEN_4189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4191 = 9'hc9 == r_count_13_io_out ? io_r_201_b : _GEN_4190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4192 = 9'hca == r_count_13_io_out ? io_r_202_b : _GEN_4191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4193 = 9'hcb == r_count_13_io_out ? io_r_203_b : _GEN_4192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4194 = 9'hcc == r_count_13_io_out ? io_r_204_b : _GEN_4193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4195 = 9'hcd == r_count_13_io_out ? io_r_205_b : _GEN_4194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4196 = 9'hce == r_count_13_io_out ? io_r_206_b : _GEN_4195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4197 = 9'hcf == r_count_13_io_out ? io_r_207_b : _GEN_4196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4198 = 9'hd0 == r_count_13_io_out ? io_r_208_b : _GEN_4197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4199 = 9'hd1 == r_count_13_io_out ? io_r_209_b : _GEN_4198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4200 = 9'hd2 == r_count_13_io_out ? io_r_210_b : _GEN_4199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4201 = 9'hd3 == r_count_13_io_out ? io_r_211_b : _GEN_4200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4202 = 9'hd4 == r_count_13_io_out ? io_r_212_b : _GEN_4201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4203 = 9'hd5 == r_count_13_io_out ? io_r_213_b : _GEN_4202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4204 = 9'hd6 == r_count_13_io_out ? io_r_214_b : _GEN_4203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4205 = 9'hd7 == r_count_13_io_out ? io_r_215_b : _GEN_4204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4206 = 9'hd8 == r_count_13_io_out ? io_r_216_b : _GEN_4205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4207 = 9'hd9 == r_count_13_io_out ? io_r_217_b : _GEN_4206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4208 = 9'hda == r_count_13_io_out ? io_r_218_b : _GEN_4207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4209 = 9'hdb == r_count_13_io_out ? io_r_219_b : _GEN_4208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4210 = 9'hdc == r_count_13_io_out ? io_r_220_b : _GEN_4209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4211 = 9'hdd == r_count_13_io_out ? io_r_221_b : _GEN_4210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4212 = 9'hde == r_count_13_io_out ? io_r_222_b : _GEN_4211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4213 = 9'hdf == r_count_13_io_out ? io_r_223_b : _GEN_4212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4214 = 9'he0 == r_count_13_io_out ? io_r_224_b : _GEN_4213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4215 = 9'he1 == r_count_13_io_out ? io_r_225_b : _GEN_4214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4216 = 9'he2 == r_count_13_io_out ? io_r_226_b : _GEN_4215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4217 = 9'he3 == r_count_13_io_out ? io_r_227_b : _GEN_4216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4218 = 9'he4 == r_count_13_io_out ? io_r_228_b : _GEN_4217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4219 = 9'he5 == r_count_13_io_out ? io_r_229_b : _GEN_4218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4220 = 9'he6 == r_count_13_io_out ? io_r_230_b : _GEN_4219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4221 = 9'he7 == r_count_13_io_out ? io_r_231_b : _GEN_4220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4222 = 9'he8 == r_count_13_io_out ? io_r_232_b : _GEN_4221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4223 = 9'he9 == r_count_13_io_out ? io_r_233_b : _GEN_4222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4224 = 9'hea == r_count_13_io_out ? io_r_234_b : _GEN_4223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4225 = 9'heb == r_count_13_io_out ? io_r_235_b : _GEN_4224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4226 = 9'hec == r_count_13_io_out ? io_r_236_b : _GEN_4225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4227 = 9'hed == r_count_13_io_out ? io_r_237_b : _GEN_4226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4228 = 9'hee == r_count_13_io_out ? io_r_238_b : _GEN_4227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4229 = 9'hef == r_count_13_io_out ? io_r_239_b : _GEN_4228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4230 = 9'hf0 == r_count_13_io_out ? io_r_240_b : _GEN_4229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4231 = 9'hf1 == r_count_13_io_out ? io_r_241_b : _GEN_4230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4232 = 9'hf2 == r_count_13_io_out ? io_r_242_b : _GEN_4231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4233 = 9'hf3 == r_count_13_io_out ? io_r_243_b : _GEN_4232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4234 = 9'hf4 == r_count_13_io_out ? io_r_244_b : _GEN_4233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4235 = 9'hf5 == r_count_13_io_out ? io_r_245_b : _GEN_4234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4236 = 9'hf6 == r_count_13_io_out ? io_r_246_b : _GEN_4235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4237 = 9'hf7 == r_count_13_io_out ? io_r_247_b : _GEN_4236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4238 = 9'hf8 == r_count_13_io_out ? io_r_248_b : _GEN_4237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4239 = 9'hf9 == r_count_13_io_out ? io_r_249_b : _GEN_4238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4240 = 9'hfa == r_count_13_io_out ? io_r_250_b : _GEN_4239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4241 = 9'hfb == r_count_13_io_out ? io_r_251_b : _GEN_4240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4242 = 9'hfc == r_count_13_io_out ? io_r_252_b : _GEN_4241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4243 = 9'hfd == r_count_13_io_out ? io_r_253_b : _GEN_4242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4244 = 9'hfe == r_count_13_io_out ? io_r_254_b : _GEN_4243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4245 = 9'hff == r_count_13_io_out ? io_r_255_b : _GEN_4244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4246 = 9'h100 == r_count_13_io_out ? io_r_256_b : _GEN_4245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4247 = 9'h101 == r_count_13_io_out ? io_r_257_b : _GEN_4246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4248 = 9'h102 == r_count_13_io_out ? io_r_258_b : _GEN_4247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4249 = 9'h103 == r_count_13_io_out ? io_r_259_b : _GEN_4248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4250 = 9'h104 == r_count_13_io_out ? io_r_260_b : _GEN_4249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4251 = 9'h105 == r_count_13_io_out ? io_r_261_b : _GEN_4250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4252 = 9'h106 == r_count_13_io_out ? io_r_262_b : _GEN_4251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4253 = 9'h107 == r_count_13_io_out ? io_r_263_b : _GEN_4252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4254 = 9'h108 == r_count_13_io_out ? io_r_264_b : _GEN_4253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4255 = 9'h109 == r_count_13_io_out ? io_r_265_b : _GEN_4254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4256 = 9'h10a == r_count_13_io_out ? io_r_266_b : _GEN_4255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4257 = 9'h10b == r_count_13_io_out ? io_r_267_b : _GEN_4256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4258 = 9'h10c == r_count_13_io_out ? io_r_268_b : _GEN_4257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4259 = 9'h10d == r_count_13_io_out ? io_r_269_b : _GEN_4258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4260 = 9'h10e == r_count_13_io_out ? io_r_270_b : _GEN_4259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4261 = 9'h10f == r_count_13_io_out ? io_r_271_b : _GEN_4260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4262 = 9'h110 == r_count_13_io_out ? io_r_272_b : _GEN_4261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4263 = 9'h111 == r_count_13_io_out ? io_r_273_b : _GEN_4262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4264 = 9'h112 == r_count_13_io_out ? io_r_274_b : _GEN_4263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4265 = 9'h113 == r_count_13_io_out ? io_r_275_b : _GEN_4264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4266 = 9'h114 == r_count_13_io_out ? io_r_276_b : _GEN_4265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4267 = 9'h115 == r_count_13_io_out ? io_r_277_b : _GEN_4266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4268 = 9'h116 == r_count_13_io_out ? io_r_278_b : _GEN_4267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4269 = 9'h117 == r_count_13_io_out ? io_r_279_b : _GEN_4268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4270 = 9'h118 == r_count_13_io_out ? io_r_280_b : _GEN_4269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4271 = 9'h119 == r_count_13_io_out ? io_r_281_b : _GEN_4270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4272 = 9'h11a == r_count_13_io_out ? io_r_282_b : _GEN_4271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4273 = 9'h11b == r_count_13_io_out ? io_r_283_b : _GEN_4272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4274 = 9'h11c == r_count_13_io_out ? io_r_284_b : _GEN_4273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4275 = 9'h11d == r_count_13_io_out ? io_r_285_b : _GEN_4274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4276 = 9'h11e == r_count_13_io_out ? io_r_286_b : _GEN_4275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4277 = 9'h11f == r_count_13_io_out ? io_r_287_b : _GEN_4276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4278 = 9'h120 == r_count_13_io_out ? io_r_288_b : _GEN_4277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4279 = 9'h121 == r_count_13_io_out ? io_r_289_b : _GEN_4278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4280 = 9'h122 == r_count_13_io_out ? io_r_290_b : _GEN_4279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4281 = 9'h123 == r_count_13_io_out ? io_r_291_b : _GEN_4280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4282 = 9'h124 == r_count_13_io_out ? io_r_292_b : _GEN_4281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4283 = 9'h125 == r_count_13_io_out ? io_r_293_b : _GEN_4282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4284 = 9'h126 == r_count_13_io_out ? io_r_294_b : _GEN_4283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4285 = 9'h127 == r_count_13_io_out ? io_r_295_b : _GEN_4284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4286 = 9'h128 == r_count_13_io_out ? io_r_296_b : _GEN_4285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4287 = 9'h129 == r_count_13_io_out ? io_r_297_b : _GEN_4286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4288 = 9'h12a == r_count_13_io_out ? io_r_298_b : _GEN_4287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4291 = 9'h1 == r_count_14_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4292 = 9'h2 == r_count_14_io_out ? io_r_2_b : _GEN_4291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4293 = 9'h3 == r_count_14_io_out ? io_r_3_b : _GEN_4292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4294 = 9'h4 == r_count_14_io_out ? io_r_4_b : _GEN_4293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4295 = 9'h5 == r_count_14_io_out ? io_r_5_b : _GEN_4294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4296 = 9'h6 == r_count_14_io_out ? io_r_6_b : _GEN_4295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4297 = 9'h7 == r_count_14_io_out ? io_r_7_b : _GEN_4296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4298 = 9'h8 == r_count_14_io_out ? io_r_8_b : _GEN_4297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4299 = 9'h9 == r_count_14_io_out ? io_r_9_b : _GEN_4298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4300 = 9'ha == r_count_14_io_out ? io_r_10_b : _GEN_4299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4301 = 9'hb == r_count_14_io_out ? io_r_11_b : _GEN_4300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4302 = 9'hc == r_count_14_io_out ? io_r_12_b : _GEN_4301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4303 = 9'hd == r_count_14_io_out ? io_r_13_b : _GEN_4302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4304 = 9'he == r_count_14_io_out ? io_r_14_b : _GEN_4303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4305 = 9'hf == r_count_14_io_out ? io_r_15_b : _GEN_4304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4306 = 9'h10 == r_count_14_io_out ? io_r_16_b : _GEN_4305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4307 = 9'h11 == r_count_14_io_out ? io_r_17_b : _GEN_4306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4308 = 9'h12 == r_count_14_io_out ? io_r_18_b : _GEN_4307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4309 = 9'h13 == r_count_14_io_out ? io_r_19_b : _GEN_4308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4310 = 9'h14 == r_count_14_io_out ? io_r_20_b : _GEN_4309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4311 = 9'h15 == r_count_14_io_out ? io_r_21_b : _GEN_4310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4312 = 9'h16 == r_count_14_io_out ? io_r_22_b : _GEN_4311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4313 = 9'h17 == r_count_14_io_out ? io_r_23_b : _GEN_4312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4314 = 9'h18 == r_count_14_io_out ? io_r_24_b : _GEN_4313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4315 = 9'h19 == r_count_14_io_out ? io_r_25_b : _GEN_4314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4316 = 9'h1a == r_count_14_io_out ? io_r_26_b : _GEN_4315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4317 = 9'h1b == r_count_14_io_out ? io_r_27_b : _GEN_4316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4318 = 9'h1c == r_count_14_io_out ? io_r_28_b : _GEN_4317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4319 = 9'h1d == r_count_14_io_out ? io_r_29_b : _GEN_4318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4320 = 9'h1e == r_count_14_io_out ? io_r_30_b : _GEN_4319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4321 = 9'h1f == r_count_14_io_out ? io_r_31_b : _GEN_4320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4322 = 9'h20 == r_count_14_io_out ? io_r_32_b : _GEN_4321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4323 = 9'h21 == r_count_14_io_out ? io_r_33_b : _GEN_4322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4324 = 9'h22 == r_count_14_io_out ? io_r_34_b : _GEN_4323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4325 = 9'h23 == r_count_14_io_out ? io_r_35_b : _GEN_4324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4326 = 9'h24 == r_count_14_io_out ? io_r_36_b : _GEN_4325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4327 = 9'h25 == r_count_14_io_out ? io_r_37_b : _GEN_4326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4328 = 9'h26 == r_count_14_io_out ? io_r_38_b : _GEN_4327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4329 = 9'h27 == r_count_14_io_out ? io_r_39_b : _GEN_4328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4330 = 9'h28 == r_count_14_io_out ? io_r_40_b : _GEN_4329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4331 = 9'h29 == r_count_14_io_out ? io_r_41_b : _GEN_4330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4332 = 9'h2a == r_count_14_io_out ? io_r_42_b : _GEN_4331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4333 = 9'h2b == r_count_14_io_out ? io_r_43_b : _GEN_4332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4334 = 9'h2c == r_count_14_io_out ? io_r_44_b : _GEN_4333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4335 = 9'h2d == r_count_14_io_out ? io_r_45_b : _GEN_4334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4336 = 9'h2e == r_count_14_io_out ? io_r_46_b : _GEN_4335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4337 = 9'h2f == r_count_14_io_out ? io_r_47_b : _GEN_4336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4338 = 9'h30 == r_count_14_io_out ? io_r_48_b : _GEN_4337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4339 = 9'h31 == r_count_14_io_out ? io_r_49_b : _GEN_4338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4340 = 9'h32 == r_count_14_io_out ? io_r_50_b : _GEN_4339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4341 = 9'h33 == r_count_14_io_out ? io_r_51_b : _GEN_4340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4342 = 9'h34 == r_count_14_io_out ? io_r_52_b : _GEN_4341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4343 = 9'h35 == r_count_14_io_out ? io_r_53_b : _GEN_4342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4344 = 9'h36 == r_count_14_io_out ? io_r_54_b : _GEN_4343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4345 = 9'h37 == r_count_14_io_out ? io_r_55_b : _GEN_4344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4346 = 9'h38 == r_count_14_io_out ? io_r_56_b : _GEN_4345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4347 = 9'h39 == r_count_14_io_out ? io_r_57_b : _GEN_4346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4348 = 9'h3a == r_count_14_io_out ? io_r_58_b : _GEN_4347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4349 = 9'h3b == r_count_14_io_out ? io_r_59_b : _GEN_4348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4350 = 9'h3c == r_count_14_io_out ? io_r_60_b : _GEN_4349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4351 = 9'h3d == r_count_14_io_out ? io_r_61_b : _GEN_4350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4352 = 9'h3e == r_count_14_io_out ? io_r_62_b : _GEN_4351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4353 = 9'h3f == r_count_14_io_out ? io_r_63_b : _GEN_4352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4354 = 9'h40 == r_count_14_io_out ? io_r_64_b : _GEN_4353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4355 = 9'h41 == r_count_14_io_out ? io_r_65_b : _GEN_4354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4356 = 9'h42 == r_count_14_io_out ? io_r_66_b : _GEN_4355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4357 = 9'h43 == r_count_14_io_out ? io_r_67_b : _GEN_4356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4358 = 9'h44 == r_count_14_io_out ? io_r_68_b : _GEN_4357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4359 = 9'h45 == r_count_14_io_out ? io_r_69_b : _GEN_4358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4360 = 9'h46 == r_count_14_io_out ? io_r_70_b : _GEN_4359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4361 = 9'h47 == r_count_14_io_out ? io_r_71_b : _GEN_4360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4362 = 9'h48 == r_count_14_io_out ? io_r_72_b : _GEN_4361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4363 = 9'h49 == r_count_14_io_out ? io_r_73_b : _GEN_4362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4364 = 9'h4a == r_count_14_io_out ? io_r_74_b : _GEN_4363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4365 = 9'h4b == r_count_14_io_out ? io_r_75_b : _GEN_4364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4366 = 9'h4c == r_count_14_io_out ? io_r_76_b : _GEN_4365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4367 = 9'h4d == r_count_14_io_out ? io_r_77_b : _GEN_4366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4368 = 9'h4e == r_count_14_io_out ? io_r_78_b : _GEN_4367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4369 = 9'h4f == r_count_14_io_out ? io_r_79_b : _GEN_4368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4370 = 9'h50 == r_count_14_io_out ? io_r_80_b : _GEN_4369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4371 = 9'h51 == r_count_14_io_out ? io_r_81_b : _GEN_4370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4372 = 9'h52 == r_count_14_io_out ? io_r_82_b : _GEN_4371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4373 = 9'h53 == r_count_14_io_out ? io_r_83_b : _GEN_4372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4374 = 9'h54 == r_count_14_io_out ? io_r_84_b : _GEN_4373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4375 = 9'h55 == r_count_14_io_out ? io_r_85_b : _GEN_4374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4376 = 9'h56 == r_count_14_io_out ? io_r_86_b : _GEN_4375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4377 = 9'h57 == r_count_14_io_out ? io_r_87_b : _GEN_4376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4378 = 9'h58 == r_count_14_io_out ? io_r_88_b : _GEN_4377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4379 = 9'h59 == r_count_14_io_out ? io_r_89_b : _GEN_4378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4380 = 9'h5a == r_count_14_io_out ? io_r_90_b : _GEN_4379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4381 = 9'h5b == r_count_14_io_out ? io_r_91_b : _GEN_4380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4382 = 9'h5c == r_count_14_io_out ? io_r_92_b : _GEN_4381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4383 = 9'h5d == r_count_14_io_out ? io_r_93_b : _GEN_4382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4384 = 9'h5e == r_count_14_io_out ? io_r_94_b : _GEN_4383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4385 = 9'h5f == r_count_14_io_out ? io_r_95_b : _GEN_4384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4386 = 9'h60 == r_count_14_io_out ? io_r_96_b : _GEN_4385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4387 = 9'h61 == r_count_14_io_out ? io_r_97_b : _GEN_4386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4388 = 9'h62 == r_count_14_io_out ? io_r_98_b : _GEN_4387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4389 = 9'h63 == r_count_14_io_out ? io_r_99_b : _GEN_4388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4390 = 9'h64 == r_count_14_io_out ? io_r_100_b : _GEN_4389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4391 = 9'h65 == r_count_14_io_out ? io_r_101_b : _GEN_4390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4392 = 9'h66 == r_count_14_io_out ? io_r_102_b : _GEN_4391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4393 = 9'h67 == r_count_14_io_out ? io_r_103_b : _GEN_4392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4394 = 9'h68 == r_count_14_io_out ? io_r_104_b : _GEN_4393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4395 = 9'h69 == r_count_14_io_out ? io_r_105_b : _GEN_4394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4396 = 9'h6a == r_count_14_io_out ? io_r_106_b : _GEN_4395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4397 = 9'h6b == r_count_14_io_out ? io_r_107_b : _GEN_4396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4398 = 9'h6c == r_count_14_io_out ? io_r_108_b : _GEN_4397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4399 = 9'h6d == r_count_14_io_out ? io_r_109_b : _GEN_4398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4400 = 9'h6e == r_count_14_io_out ? io_r_110_b : _GEN_4399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4401 = 9'h6f == r_count_14_io_out ? io_r_111_b : _GEN_4400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4402 = 9'h70 == r_count_14_io_out ? io_r_112_b : _GEN_4401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4403 = 9'h71 == r_count_14_io_out ? io_r_113_b : _GEN_4402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4404 = 9'h72 == r_count_14_io_out ? io_r_114_b : _GEN_4403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4405 = 9'h73 == r_count_14_io_out ? io_r_115_b : _GEN_4404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4406 = 9'h74 == r_count_14_io_out ? io_r_116_b : _GEN_4405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4407 = 9'h75 == r_count_14_io_out ? io_r_117_b : _GEN_4406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4408 = 9'h76 == r_count_14_io_out ? io_r_118_b : _GEN_4407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4409 = 9'h77 == r_count_14_io_out ? io_r_119_b : _GEN_4408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4410 = 9'h78 == r_count_14_io_out ? io_r_120_b : _GEN_4409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4411 = 9'h79 == r_count_14_io_out ? io_r_121_b : _GEN_4410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4412 = 9'h7a == r_count_14_io_out ? io_r_122_b : _GEN_4411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4413 = 9'h7b == r_count_14_io_out ? io_r_123_b : _GEN_4412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4414 = 9'h7c == r_count_14_io_out ? io_r_124_b : _GEN_4413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4415 = 9'h7d == r_count_14_io_out ? io_r_125_b : _GEN_4414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4416 = 9'h7e == r_count_14_io_out ? io_r_126_b : _GEN_4415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4417 = 9'h7f == r_count_14_io_out ? io_r_127_b : _GEN_4416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4418 = 9'h80 == r_count_14_io_out ? io_r_128_b : _GEN_4417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4419 = 9'h81 == r_count_14_io_out ? io_r_129_b : _GEN_4418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4420 = 9'h82 == r_count_14_io_out ? io_r_130_b : _GEN_4419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4421 = 9'h83 == r_count_14_io_out ? io_r_131_b : _GEN_4420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4422 = 9'h84 == r_count_14_io_out ? io_r_132_b : _GEN_4421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4423 = 9'h85 == r_count_14_io_out ? io_r_133_b : _GEN_4422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4424 = 9'h86 == r_count_14_io_out ? io_r_134_b : _GEN_4423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4425 = 9'h87 == r_count_14_io_out ? io_r_135_b : _GEN_4424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4426 = 9'h88 == r_count_14_io_out ? io_r_136_b : _GEN_4425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4427 = 9'h89 == r_count_14_io_out ? io_r_137_b : _GEN_4426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4428 = 9'h8a == r_count_14_io_out ? io_r_138_b : _GEN_4427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4429 = 9'h8b == r_count_14_io_out ? io_r_139_b : _GEN_4428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4430 = 9'h8c == r_count_14_io_out ? io_r_140_b : _GEN_4429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4431 = 9'h8d == r_count_14_io_out ? io_r_141_b : _GEN_4430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4432 = 9'h8e == r_count_14_io_out ? io_r_142_b : _GEN_4431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4433 = 9'h8f == r_count_14_io_out ? io_r_143_b : _GEN_4432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4434 = 9'h90 == r_count_14_io_out ? io_r_144_b : _GEN_4433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4435 = 9'h91 == r_count_14_io_out ? io_r_145_b : _GEN_4434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4436 = 9'h92 == r_count_14_io_out ? io_r_146_b : _GEN_4435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4437 = 9'h93 == r_count_14_io_out ? io_r_147_b : _GEN_4436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4438 = 9'h94 == r_count_14_io_out ? io_r_148_b : _GEN_4437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4439 = 9'h95 == r_count_14_io_out ? io_r_149_b : _GEN_4438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4440 = 9'h96 == r_count_14_io_out ? io_r_150_b : _GEN_4439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4441 = 9'h97 == r_count_14_io_out ? io_r_151_b : _GEN_4440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4442 = 9'h98 == r_count_14_io_out ? io_r_152_b : _GEN_4441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4443 = 9'h99 == r_count_14_io_out ? io_r_153_b : _GEN_4442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4444 = 9'h9a == r_count_14_io_out ? io_r_154_b : _GEN_4443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4445 = 9'h9b == r_count_14_io_out ? io_r_155_b : _GEN_4444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4446 = 9'h9c == r_count_14_io_out ? io_r_156_b : _GEN_4445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4447 = 9'h9d == r_count_14_io_out ? io_r_157_b : _GEN_4446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4448 = 9'h9e == r_count_14_io_out ? io_r_158_b : _GEN_4447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4449 = 9'h9f == r_count_14_io_out ? io_r_159_b : _GEN_4448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4450 = 9'ha0 == r_count_14_io_out ? io_r_160_b : _GEN_4449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4451 = 9'ha1 == r_count_14_io_out ? io_r_161_b : _GEN_4450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4452 = 9'ha2 == r_count_14_io_out ? io_r_162_b : _GEN_4451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4453 = 9'ha3 == r_count_14_io_out ? io_r_163_b : _GEN_4452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4454 = 9'ha4 == r_count_14_io_out ? io_r_164_b : _GEN_4453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4455 = 9'ha5 == r_count_14_io_out ? io_r_165_b : _GEN_4454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4456 = 9'ha6 == r_count_14_io_out ? io_r_166_b : _GEN_4455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4457 = 9'ha7 == r_count_14_io_out ? io_r_167_b : _GEN_4456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4458 = 9'ha8 == r_count_14_io_out ? io_r_168_b : _GEN_4457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4459 = 9'ha9 == r_count_14_io_out ? io_r_169_b : _GEN_4458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4460 = 9'haa == r_count_14_io_out ? io_r_170_b : _GEN_4459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4461 = 9'hab == r_count_14_io_out ? io_r_171_b : _GEN_4460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4462 = 9'hac == r_count_14_io_out ? io_r_172_b : _GEN_4461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4463 = 9'had == r_count_14_io_out ? io_r_173_b : _GEN_4462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4464 = 9'hae == r_count_14_io_out ? io_r_174_b : _GEN_4463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4465 = 9'haf == r_count_14_io_out ? io_r_175_b : _GEN_4464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4466 = 9'hb0 == r_count_14_io_out ? io_r_176_b : _GEN_4465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4467 = 9'hb1 == r_count_14_io_out ? io_r_177_b : _GEN_4466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4468 = 9'hb2 == r_count_14_io_out ? io_r_178_b : _GEN_4467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4469 = 9'hb3 == r_count_14_io_out ? io_r_179_b : _GEN_4468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4470 = 9'hb4 == r_count_14_io_out ? io_r_180_b : _GEN_4469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4471 = 9'hb5 == r_count_14_io_out ? io_r_181_b : _GEN_4470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4472 = 9'hb6 == r_count_14_io_out ? io_r_182_b : _GEN_4471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4473 = 9'hb7 == r_count_14_io_out ? io_r_183_b : _GEN_4472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4474 = 9'hb8 == r_count_14_io_out ? io_r_184_b : _GEN_4473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4475 = 9'hb9 == r_count_14_io_out ? io_r_185_b : _GEN_4474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4476 = 9'hba == r_count_14_io_out ? io_r_186_b : _GEN_4475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4477 = 9'hbb == r_count_14_io_out ? io_r_187_b : _GEN_4476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4478 = 9'hbc == r_count_14_io_out ? io_r_188_b : _GEN_4477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4479 = 9'hbd == r_count_14_io_out ? io_r_189_b : _GEN_4478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4480 = 9'hbe == r_count_14_io_out ? io_r_190_b : _GEN_4479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4481 = 9'hbf == r_count_14_io_out ? io_r_191_b : _GEN_4480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4482 = 9'hc0 == r_count_14_io_out ? io_r_192_b : _GEN_4481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4483 = 9'hc1 == r_count_14_io_out ? io_r_193_b : _GEN_4482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4484 = 9'hc2 == r_count_14_io_out ? io_r_194_b : _GEN_4483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4485 = 9'hc3 == r_count_14_io_out ? io_r_195_b : _GEN_4484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4486 = 9'hc4 == r_count_14_io_out ? io_r_196_b : _GEN_4485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4487 = 9'hc5 == r_count_14_io_out ? io_r_197_b : _GEN_4486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4488 = 9'hc6 == r_count_14_io_out ? io_r_198_b : _GEN_4487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4489 = 9'hc7 == r_count_14_io_out ? io_r_199_b : _GEN_4488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4490 = 9'hc8 == r_count_14_io_out ? io_r_200_b : _GEN_4489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4491 = 9'hc9 == r_count_14_io_out ? io_r_201_b : _GEN_4490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4492 = 9'hca == r_count_14_io_out ? io_r_202_b : _GEN_4491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4493 = 9'hcb == r_count_14_io_out ? io_r_203_b : _GEN_4492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4494 = 9'hcc == r_count_14_io_out ? io_r_204_b : _GEN_4493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4495 = 9'hcd == r_count_14_io_out ? io_r_205_b : _GEN_4494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4496 = 9'hce == r_count_14_io_out ? io_r_206_b : _GEN_4495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4497 = 9'hcf == r_count_14_io_out ? io_r_207_b : _GEN_4496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4498 = 9'hd0 == r_count_14_io_out ? io_r_208_b : _GEN_4497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4499 = 9'hd1 == r_count_14_io_out ? io_r_209_b : _GEN_4498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4500 = 9'hd2 == r_count_14_io_out ? io_r_210_b : _GEN_4499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4501 = 9'hd3 == r_count_14_io_out ? io_r_211_b : _GEN_4500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4502 = 9'hd4 == r_count_14_io_out ? io_r_212_b : _GEN_4501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4503 = 9'hd5 == r_count_14_io_out ? io_r_213_b : _GEN_4502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4504 = 9'hd6 == r_count_14_io_out ? io_r_214_b : _GEN_4503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4505 = 9'hd7 == r_count_14_io_out ? io_r_215_b : _GEN_4504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4506 = 9'hd8 == r_count_14_io_out ? io_r_216_b : _GEN_4505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4507 = 9'hd9 == r_count_14_io_out ? io_r_217_b : _GEN_4506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4508 = 9'hda == r_count_14_io_out ? io_r_218_b : _GEN_4507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4509 = 9'hdb == r_count_14_io_out ? io_r_219_b : _GEN_4508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4510 = 9'hdc == r_count_14_io_out ? io_r_220_b : _GEN_4509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4511 = 9'hdd == r_count_14_io_out ? io_r_221_b : _GEN_4510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4512 = 9'hde == r_count_14_io_out ? io_r_222_b : _GEN_4511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4513 = 9'hdf == r_count_14_io_out ? io_r_223_b : _GEN_4512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4514 = 9'he0 == r_count_14_io_out ? io_r_224_b : _GEN_4513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4515 = 9'he1 == r_count_14_io_out ? io_r_225_b : _GEN_4514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4516 = 9'he2 == r_count_14_io_out ? io_r_226_b : _GEN_4515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4517 = 9'he3 == r_count_14_io_out ? io_r_227_b : _GEN_4516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4518 = 9'he4 == r_count_14_io_out ? io_r_228_b : _GEN_4517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4519 = 9'he5 == r_count_14_io_out ? io_r_229_b : _GEN_4518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4520 = 9'he6 == r_count_14_io_out ? io_r_230_b : _GEN_4519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4521 = 9'he7 == r_count_14_io_out ? io_r_231_b : _GEN_4520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4522 = 9'he8 == r_count_14_io_out ? io_r_232_b : _GEN_4521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4523 = 9'he9 == r_count_14_io_out ? io_r_233_b : _GEN_4522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4524 = 9'hea == r_count_14_io_out ? io_r_234_b : _GEN_4523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4525 = 9'heb == r_count_14_io_out ? io_r_235_b : _GEN_4524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4526 = 9'hec == r_count_14_io_out ? io_r_236_b : _GEN_4525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4527 = 9'hed == r_count_14_io_out ? io_r_237_b : _GEN_4526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4528 = 9'hee == r_count_14_io_out ? io_r_238_b : _GEN_4527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4529 = 9'hef == r_count_14_io_out ? io_r_239_b : _GEN_4528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4530 = 9'hf0 == r_count_14_io_out ? io_r_240_b : _GEN_4529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4531 = 9'hf1 == r_count_14_io_out ? io_r_241_b : _GEN_4530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4532 = 9'hf2 == r_count_14_io_out ? io_r_242_b : _GEN_4531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4533 = 9'hf3 == r_count_14_io_out ? io_r_243_b : _GEN_4532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4534 = 9'hf4 == r_count_14_io_out ? io_r_244_b : _GEN_4533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4535 = 9'hf5 == r_count_14_io_out ? io_r_245_b : _GEN_4534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4536 = 9'hf6 == r_count_14_io_out ? io_r_246_b : _GEN_4535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4537 = 9'hf7 == r_count_14_io_out ? io_r_247_b : _GEN_4536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4538 = 9'hf8 == r_count_14_io_out ? io_r_248_b : _GEN_4537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4539 = 9'hf9 == r_count_14_io_out ? io_r_249_b : _GEN_4538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4540 = 9'hfa == r_count_14_io_out ? io_r_250_b : _GEN_4539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4541 = 9'hfb == r_count_14_io_out ? io_r_251_b : _GEN_4540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4542 = 9'hfc == r_count_14_io_out ? io_r_252_b : _GEN_4541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4543 = 9'hfd == r_count_14_io_out ? io_r_253_b : _GEN_4542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4544 = 9'hfe == r_count_14_io_out ? io_r_254_b : _GEN_4543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4545 = 9'hff == r_count_14_io_out ? io_r_255_b : _GEN_4544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4546 = 9'h100 == r_count_14_io_out ? io_r_256_b : _GEN_4545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4547 = 9'h101 == r_count_14_io_out ? io_r_257_b : _GEN_4546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4548 = 9'h102 == r_count_14_io_out ? io_r_258_b : _GEN_4547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4549 = 9'h103 == r_count_14_io_out ? io_r_259_b : _GEN_4548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4550 = 9'h104 == r_count_14_io_out ? io_r_260_b : _GEN_4549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4551 = 9'h105 == r_count_14_io_out ? io_r_261_b : _GEN_4550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4552 = 9'h106 == r_count_14_io_out ? io_r_262_b : _GEN_4551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4553 = 9'h107 == r_count_14_io_out ? io_r_263_b : _GEN_4552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4554 = 9'h108 == r_count_14_io_out ? io_r_264_b : _GEN_4553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4555 = 9'h109 == r_count_14_io_out ? io_r_265_b : _GEN_4554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4556 = 9'h10a == r_count_14_io_out ? io_r_266_b : _GEN_4555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4557 = 9'h10b == r_count_14_io_out ? io_r_267_b : _GEN_4556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4558 = 9'h10c == r_count_14_io_out ? io_r_268_b : _GEN_4557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4559 = 9'h10d == r_count_14_io_out ? io_r_269_b : _GEN_4558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4560 = 9'h10e == r_count_14_io_out ? io_r_270_b : _GEN_4559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4561 = 9'h10f == r_count_14_io_out ? io_r_271_b : _GEN_4560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4562 = 9'h110 == r_count_14_io_out ? io_r_272_b : _GEN_4561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4563 = 9'h111 == r_count_14_io_out ? io_r_273_b : _GEN_4562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4564 = 9'h112 == r_count_14_io_out ? io_r_274_b : _GEN_4563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4565 = 9'h113 == r_count_14_io_out ? io_r_275_b : _GEN_4564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4566 = 9'h114 == r_count_14_io_out ? io_r_276_b : _GEN_4565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4567 = 9'h115 == r_count_14_io_out ? io_r_277_b : _GEN_4566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4568 = 9'h116 == r_count_14_io_out ? io_r_278_b : _GEN_4567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4569 = 9'h117 == r_count_14_io_out ? io_r_279_b : _GEN_4568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4570 = 9'h118 == r_count_14_io_out ? io_r_280_b : _GEN_4569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4571 = 9'h119 == r_count_14_io_out ? io_r_281_b : _GEN_4570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4572 = 9'h11a == r_count_14_io_out ? io_r_282_b : _GEN_4571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4573 = 9'h11b == r_count_14_io_out ? io_r_283_b : _GEN_4572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4574 = 9'h11c == r_count_14_io_out ? io_r_284_b : _GEN_4573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4575 = 9'h11d == r_count_14_io_out ? io_r_285_b : _GEN_4574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4576 = 9'h11e == r_count_14_io_out ? io_r_286_b : _GEN_4575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4577 = 9'h11f == r_count_14_io_out ? io_r_287_b : _GEN_4576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4578 = 9'h120 == r_count_14_io_out ? io_r_288_b : _GEN_4577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4579 = 9'h121 == r_count_14_io_out ? io_r_289_b : _GEN_4578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4580 = 9'h122 == r_count_14_io_out ? io_r_290_b : _GEN_4579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4581 = 9'h123 == r_count_14_io_out ? io_r_291_b : _GEN_4580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4582 = 9'h124 == r_count_14_io_out ? io_r_292_b : _GEN_4581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4583 = 9'h125 == r_count_14_io_out ? io_r_293_b : _GEN_4582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4584 = 9'h126 == r_count_14_io_out ? io_r_294_b : _GEN_4583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4585 = 9'h127 == r_count_14_io_out ? io_r_295_b : _GEN_4584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4586 = 9'h128 == r_count_14_io_out ? io_r_296_b : _GEN_4585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4587 = 9'h129 == r_count_14_io_out ? io_r_297_b : _GEN_4586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4588 = 9'h12a == r_count_14_io_out ? io_r_298_b : _GEN_4587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4591 = 9'h1 == r_count_15_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4592 = 9'h2 == r_count_15_io_out ? io_r_2_b : _GEN_4591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4593 = 9'h3 == r_count_15_io_out ? io_r_3_b : _GEN_4592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4594 = 9'h4 == r_count_15_io_out ? io_r_4_b : _GEN_4593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4595 = 9'h5 == r_count_15_io_out ? io_r_5_b : _GEN_4594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4596 = 9'h6 == r_count_15_io_out ? io_r_6_b : _GEN_4595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4597 = 9'h7 == r_count_15_io_out ? io_r_7_b : _GEN_4596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4598 = 9'h8 == r_count_15_io_out ? io_r_8_b : _GEN_4597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4599 = 9'h9 == r_count_15_io_out ? io_r_9_b : _GEN_4598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4600 = 9'ha == r_count_15_io_out ? io_r_10_b : _GEN_4599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4601 = 9'hb == r_count_15_io_out ? io_r_11_b : _GEN_4600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4602 = 9'hc == r_count_15_io_out ? io_r_12_b : _GEN_4601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4603 = 9'hd == r_count_15_io_out ? io_r_13_b : _GEN_4602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4604 = 9'he == r_count_15_io_out ? io_r_14_b : _GEN_4603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4605 = 9'hf == r_count_15_io_out ? io_r_15_b : _GEN_4604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4606 = 9'h10 == r_count_15_io_out ? io_r_16_b : _GEN_4605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4607 = 9'h11 == r_count_15_io_out ? io_r_17_b : _GEN_4606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4608 = 9'h12 == r_count_15_io_out ? io_r_18_b : _GEN_4607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4609 = 9'h13 == r_count_15_io_out ? io_r_19_b : _GEN_4608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4610 = 9'h14 == r_count_15_io_out ? io_r_20_b : _GEN_4609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4611 = 9'h15 == r_count_15_io_out ? io_r_21_b : _GEN_4610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4612 = 9'h16 == r_count_15_io_out ? io_r_22_b : _GEN_4611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4613 = 9'h17 == r_count_15_io_out ? io_r_23_b : _GEN_4612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4614 = 9'h18 == r_count_15_io_out ? io_r_24_b : _GEN_4613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4615 = 9'h19 == r_count_15_io_out ? io_r_25_b : _GEN_4614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4616 = 9'h1a == r_count_15_io_out ? io_r_26_b : _GEN_4615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4617 = 9'h1b == r_count_15_io_out ? io_r_27_b : _GEN_4616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4618 = 9'h1c == r_count_15_io_out ? io_r_28_b : _GEN_4617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4619 = 9'h1d == r_count_15_io_out ? io_r_29_b : _GEN_4618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4620 = 9'h1e == r_count_15_io_out ? io_r_30_b : _GEN_4619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4621 = 9'h1f == r_count_15_io_out ? io_r_31_b : _GEN_4620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4622 = 9'h20 == r_count_15_io_out ? io_r_32_b : _GEN_4621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4623 = 9'h21 == r_count_15_io_out ? io_r_33_b : _GEN_4622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4624 = 9'h22 == r_count_15_io_out ? io_r_34_b : _GEN_4623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4625 = 9'h23 == r_count_15_io_out ? io_r_35_b : _GEN_4624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4626 = 9'h24 == r_count_15_io_out ? io_r_36_b : _GEN_4625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4627 = 9'h25 == r_count_15_io_out ? io_r_37_b : _GEN_4626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4628 = 9'h26 == r_count_15_io_out ? io_r_38_b : _GEN_4627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4629 = 9'h27 == r_count_15_io_out ? io_r_39_b : _GEN_4628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4630 = 9'h28 == r_count_15_io_out ? io_r_40_b : _GEN_4629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4631 = 9'h29 == r_count_15_io_out ? io_r_41_b : _GEN_4630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4632 = 9'h2a == r_count_15_io_out ? io_r_42_b : _GEN_4631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4633 = 9'h2b == r_count_15_io_out ? io_r_43_b : _GEN_4632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4634 = 9'h2c == r_count_15_io_out ? io_r_44_b : _GEN_4633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4635 = 9'h2d == r_count_15_io_out ? io_r_45_b : _GEN_4634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4636 = 9'h2e == r_count_15_io_out ? io_r_46_b : _GEN_4635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4637 = 9'h2f == r_count_15_io_out ? io_r_47_b : _GEN_4636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4638 = 9'h30 == r_count_15_io_out ? io_r_48_b : _GEN_4637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4639 = 9'h31 == r_count_15_io_out ? io_r_49_b : _GEN_4638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4640 = 9'h32 == r_count_15_io_out ? io_r_50_b : _GEN_4639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4641 = 9'h33 == r_count_15_io_out ? io_r_51_b : _GEN_4640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4642 = 9'h34 == r_count_15_io_out ? io_r_52_b : _GEN_4641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4643 = 9'h35 == r_count_15_io_out ? io_r_53_b : _GEN_4642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4644 = 9'h36 == r_count_15_io_out ? io_r_54_b : _GEN_4643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4645 = 9'h37 == r_count_15_io_out ? io_r_55_b : _GEN_4644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4646 = 9'h38 == r_count_15_io_out ? io_r_56_b : _GEN_4645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4647 = 9'h39 == r_count_15_io_out ? io_r_57_b : _GEN_4646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4648 = 9'h3a == r_count_15_io_out ? io_r_58_b : _GEN_4647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4649 = 9'h3b == r_count_15_io_out ? io_r_59_b : _GEN_4648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4650 = 9'h3c == r_count_15_io_out ? io_r_60_b : _GEN_4649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4651 = 9'h3d == r_count_15_io_out ? io_r_61_b : _GEN_4650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4652 = 9'h3e == r_count_15_io_out ? io_r_62_b : _GEN_4651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4653 = 9'h3f == r_count_15_io_out ? io_r_63_b : _GEN_4652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4654 = 9'h40 == r_count_15_io_out ? io_r_64_b : _GEN_4653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4655 = 9'h41 == r_count_15_io_out ? io_r_65_b : _GEN_4654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4656 = 9'h42 == r_count_15_io_out ? io_r_66_b : _GEN_4655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4657 = 9'h43 == r_count_15_io_out ? io_r_67_b : _GEN_4656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4658 = 9'h44 == r_count_15_io_out ? io_r_68_b : _GEN_4657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4659 = 9'h45 == r_count_15_io_out ? io_r_69_b : _GEN_4658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4660 = 9'h46 == r_count_15_io_out ? io_r_70_b : _GEN_4659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4661 = 9'h47 == r_count_15_io_out ? io_r_71_b : _GEN_4660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4662 = 9'h48 == r_count_15_io_out ? io_r_72_b : _GEN_4661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4663 = 9'h49 == r_count_15_io_out ? io_r_73_b : _GEN_4662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4664 = 9'h4a == r_count_15_io_out ? io_r_74_b : _GEN_4663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4665 = 9'h4b == r_count_15_io_out ? io_r_75_b : _GEN_4664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4666 = 9'h4c == r_count_15_io_out ? io_r_76_b : _GEN_4665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4667 = 9'h4d == r_count_15_io_out ? io_r_77_b : _GEN_4666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4668 = 9'h4e == r_count_15_io_out ? io_r_78_b : _GEN_4667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4669 = 9'h4f == r_count_15_io_out ? io_r_79_b : _GEN_4668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4670 = 9'h50 == r_count_15_io_out ? io_r_80_b : _GEN_4669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4671 = 9'h51 == r_count_15_io_out ? io_r_81_b : _GEN_4670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4672 = 9'h52 == r_count_15_io_out ? io_r_82_b : _GEN_4671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4673 = 9'h53 == r_count_15_io_out ? io_r_83_b : _GEN_4672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4674 = 9'h54 == r_count_15_io_out ? io_r_84_b : _GEN_4673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4675 = 9'h55 == r_count_15_io_out ? io_r_85_b : _GEN_4674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4676 = 9'h56 == r_count_15_io_out ? io_r_86_b : _GEN_4675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4677 = 9'h57 == r_count_15_io_out ? io_r_87_b : _GEN_4676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4678 = 9'h58 == r_count_15_io_out ? io_r_88_b : _GEN_4677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4679 = 9'h59 == r_count_15_io_out ? io_r_89_b : _GEN_4678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4680 = 9'h5a == r_count_15_io_out ? io_r_90_b : _GEN_4679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4681 = 9'h5b == r_count_15_io_out ? io_r_91_b : _GEN_4680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4682 = 9'h5c == r_count_15_io_out ? io_r_92_b : _GEN_4681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4683 = 9'h5d == r_count_15_io_out ? io_r_93_b : _GEN_4682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4684 = 9'h5e == r_count_15_io_out ? io_r_94_b : _GEN_4683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4685 = 9'h5f == r_count_15_io_out ? io_r_95_b : _GEN_4684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4686 = 9'h60 == r_count_15_io_out ? io_r_96_b : _GEN_4685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4687 = 9'h61 == r_count_15_io_out ? io_r_97_b : _GEN_4686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4688 = 9'h62 == r_count_15_io_out ? io_r_98_b : _GEN_4687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4689 = 9'h63 == r_count_15_io_out ? io_r_99_b : _GEN_4688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4690 = 9'h64 == r_count_15_io_out ? io_r_100_b : _GEN_4689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4691 = 9'h65 == r_count_15_io_out ? io_r_101_b : _GEN_4690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4692 = 9'h66 == r_count_15_io_out ? io_r_102_b : _GEN_4691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4693 = 9'h67 == r_count_15_io_out ? io_r_103_b : _GEN_4692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4694 = 9'h68 == r_count_15_io_out ? io_r_104_b : _GEN_4693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4695 = 9'h69 == r_count_15_io_out ? io_r_105_b : _GEN_4694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4696 = 9'h6a == r_count_15_io_out ? io_r_106_b : _GEN_4695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4697 = 9'h6b == r_count_15_io_out ? io_r_107_b : _GEN_4696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4698 = 9'h6c == r_count_15_io_out ? io_r_108_b : _GEN_4697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4699 = 9'h6d == r_count_15_io_out ? io_r_109_b : _GEN_4698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4700 = 9'h6e == r_count_15_io_out ? io_r_110_b : _GEN_4699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4701 = 9'h6f == r_count_15_io_out ? io_r_111_b : _GEN_4700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4702 = 9'h70 == r_count_15_io_out ? io_r_112_b : _GEN_4701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4703 = 9'h71 == r_count_15_io_out ? io_r_113_b : _GEN_4702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4704 = 9'h72 == r_count_15_io_out ? io_r_114_b : _GEN_4703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4705 = 9'h73 == r_count_15_io_out ? io_r_115_b : _GEN_4704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4706 = 9'h74 == r_count_15_io_out ? io_r_116_b : _GEN_4705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4707 = 9'h75 == r_count_15_io_out ? io_r_117_b : _GEN_4706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4708 = 9'h76 == r_count_15_io_out ? io_r_118_b : _GEN_4707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4709 = 9'h77 == r_count_15_io_out ? io_r_119_b : _GEN_4708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4710 = 9'h78 == r_count_15_io_out ? io_r_120_b : _GEN_4709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4711 = 9'h79 == r_count_15_io_out ? io_r_121_b : _GEN_4710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4712 = 9'h7a == r_count_15_io_out ? io_r_122_b : _GEN_4711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4713 = 9'h7b == r_count_15_io_out ? io_r_123_b : _GEN_4712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4714 = 9'h7c == r_count_15_io_out ? io_r_124_b : _GEN_4713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4715 = 9'h7d == r_count_15_io_out ? io_r_125_b : _GEN_4714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4716 = 9'h7e == r_count_15_io_out ? io_r_126_b : _GEN_4715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4717 = 9'h7f == r_count_15_io_out ? io_r_127_b : _GEN_4716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4718 = 9'h80 == r_count_15_io_out ? io_r_128_b : _GEN_4717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4719 = 9'h81 == r_count_15_io_out ? io_r_129_b : _GEN_4718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4720 = 9'h82 == r_count_15_io_out ? io_r_130_b : _GEN_4719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4721 = 9'h83 == r_count_15_io_out ? io_r_131_b : _GEN_4720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4722 = 9'h84 == r_count_15_io_out ? io_r_132_b : _GEN_4721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4723 = 9'h85 == r_count_15_io_out ? io_r_133_b : _GEN_4722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4724 = 9'h86 == r_count_15_io_out ? io_r_134_b : _GEN_4723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4725 = 9'h87 == r_count_15_io_out ? io_r_135_b : _GEN_4724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4726 = 9'h88 == r_count_15_io_out ? io_r_136_b : _GEN_4725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4727 = 9'h89 == r_count_15_io_out ? io_r_137_b : _GEN_4726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4728 = 9'h8a == r_count_15_io_out ? io_r_138_b : _GEN_4727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4729 = 9'h8b == r_count_15_io_out ? io_r_139_b : _GEN_4728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4730 = 9'h8c == r_count_15_io_out ? io_r_140_b : _GEN_4729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4731 = 9'h8d == r_count_15_io_out ? io_r_141_b : _GEN_4730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4732 = 9'h8e == r_count_15_io_out ? io_r_142_b : _GEN_4731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4733 = 9'h8f == r_count_15_io_out ? io_r_143_b : _GEN_4732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4734 = 9'h90 == r_count_15_io_out ? io_r_144_b : _GEN_4733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4735 = 9'h91 == r_count_15_io_out ? io_r_145_b : _GEN_4734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4736 = 9'h92 == r_count_15_io_out ? io_r_146_b : _GEN_4735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4737 = 9'h93 == r_count_15_io_out ? io_r_147_b : _GEN_4736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4738 = 9'h94 == r_count_15_io_out ? io_r_148_b : _GEN_4737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4739 = 9'h95 == r_count_15_io_out ? io_r_149_b : _GEN_4738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4740 = 9'h96 == r_count_15_io_out ? io_r_150_b : _GEN_4739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4741 = 9'h97 == r_count_15_io_out ? io_r_151_b : _GEN_4740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4742 = 9'h98 == r_count_15_io_out ? io_r_152_b : _GEN_4741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4743 = 9'h99 == r_count_15_io_out ? io_r_153_b : _GEN_4742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4744 = 9'h9a == r_count_15_io_out ? io_r_154_b : _GEN_4743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4745 = 9'h9b == r_count_15_io_out ? io_r_155_b : _GEN_4744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4746 = 9'h9c == r_count_15_io_out ? io_r_156_b : _GEN_4745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4747 = 9'h9d == r_count_15_io_out ? io_r_157_b : _GEN_4746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4748 = 9'h9e == r_count_15_io_out ? io_r_158_b : _GEN_4747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4749 = 9'h9f == r_count_15_io_out ? io_r_159_b : _GEN_4748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4750 = 9'ha0 == r_count_15_io_out ? io_r_160_b : _GEN_4749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4751 = 9'ha1 == r_count_15_io_out ? io_r_161_b : _GEN_4750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4752 = 9'ha2 == r_count_15_io_out ? io_r_162_b : _GEN_4751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4753 = 9'ha3 == r_count_15_io_out ? io_r_163_b : _GEN_4752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4754 = 9'ha4 == r_count_15_io_out ? io_r_164_b : _GEN_4753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4755 = 9'ha5 == r_count_15_io_out ? io_r_165_b : _GEN_4754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4756 = 9'ha6 == r_count_15_io_out ? io_r_166_b : _GEN_4755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4757 = 9'ha7 == r_count_15_io_out ? io_r_167_b : _GEN_4756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4758 = 9'ha8 == r_count_15_io_out ? io_r_168_b : _GEN_4757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4759 = 9'ha9 == r_count_15_io_out ? io_r_169_b : _GEN_4758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4760 = 9'haa == r_count_15_io_out ? io_r_170_b : _GEN_4759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4761 = 9'hab == r_count_15_io_out ? io_r_171_b : _GEN_4760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4762 = 9'hac == r_count_15_io_out ? io_r_172_b : _GEN_4761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4763 = 9'had == r_count_15_io_out ? io_r_173_b : _GEN_4762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4764 = 9'hae == r_count_15_io_out ? io_r_174_b : _GEN_4763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4765 = 9'haf == r_count_15_io_out ? io_r_175_b : _GEN_4764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4766 = 9'hb0 == r_count_15_io_out ? io_r_176_b : _GEN_4765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4767 = 9'hb1 == r_count_15_io_out ? io_r_177_b : _GEN_4766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4768 = 9'hb2 == r_count_15_io_out ? io_r_178_b : _GEN_4767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4769 = 9'hb3 == r_count_15_io_out ? io_r_179_b : _GEN_4768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4770 = 9'hb4 == r_count_15_io_out ? io_r_180_b : _GEN_4769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4771 = 9'hb5 == r_count_15_io_out ? io_r_181_b : _GEN_4770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4772 = 9'hb6 == r_count_15_io_out ? io_r_182_b : _GEN_4771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4773 = 9'hb7 == r_count_15_io_out ? io_r_183_b : _GEN_4772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4774 = 9'hb8 == r_count_15_io_out ? io_r_184_b : _GEN_4773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4775 = 9'hb9 == r_count_15_io_out ? io_r_185_b : _GEN_4774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4776 = 9'hba == r_count_15_io_out ? io_r_186_b : _GEN_4775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4777 = 9'hbb == r_count_15_io_out ? io_r_187_b : _GEN_4776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4778 = 9'hbc == r_count_15_io_out ? io_r_188_b : _GEN_4777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4779 = 9'hbd == r_count_15_io_out ? io_r_189_b : _GEN_4778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4780 = 9'hbe == r_count_15_io_out ? io_r_190_b : _GEN_4779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4781 = 9'hbf == r_count_15_io_out ? io_r_191_b : _GEN_4780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4782 = 9'hc0 == r_count_15_io_out ? io_r_192_b : _GEN_4781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4783 = 9'hc1 == r_count_15_io_out ? io_r_193_b : _GEN_4782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4784 = 9'hc2 == r_count_15_io_out ? io_r_194_b : _GEN_4783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4785 = 9'hc3 == r_count_15_io_out ? io_r_195_b : _GEN_4784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4786 = 9'hc4 == r_count_15_io_out ? io_r_196_b : _GEN_4785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4787 = 9'hc5 == r_count_15_io_out ? io_r_197_b : _GEN_4786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4788 = 9'hc6 == r_count_15_io_out ? io_r_198_b : _GEN_4787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4789 = 9'hc7 == r_count_15_io_out ? io_r_199_b : _GEN_4788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4790 = 9'hc8 == r_count_15_io_out ? io_r_200_b : _GEN_4789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4791 = 9'hc9 == r_count_15_io_out ? io_r_201_b : _GEN_4790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4792 = 9'hca == r_count_15_io_out ? io_r_202_b : _GEN_4791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4793 = 9'hcb == r_count_15_io_out ? io_r_203_b : _GEN_4792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4794 = 9'hcc == r_count_15_io_out ? io_r_204_b : _GEN_4793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4795 = 9'hcd == r_count_15_io_out ? io_r_205_b : _GEN_4794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4796 = 9'hce == r_count_15_io_out ? io_r_206_b : _GEN_4795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4797 = 9'hcf == r_count_15_io_out ? io_r_207_b : _GEN_4796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4798 = 9'hd0 == r_count_15_io_out ? io_r_208_b : _GEN_4797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4799 = 9'hd1 == r_count_15_io_out ? io_r_209_b : _GEN_4798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4800 = 9'hd2 == r_count_15_io_out ? io_r_210_b : _GEN_4799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4801 = 9'hd3 == r_count_15_io_out ? io_r_211_b : _GEN_4800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4802 = 9'hd4 == r_count_15_io_out ? io_r_212_b : _GEN_4801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4803 = 9'hd5 == r_count_15_io_out ? io_r_213_b : _GEN_4802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4804 = 9'hd6 == r_count_15_io_out ? io_r_214_b : _GEN_4803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4805 = 9'hd7 == r_count_15_io_out ? io_r_215_b : _GEN_4804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4806 = 9'hd8 == r_count_15_io_out ? io_r_216_b : _GEN_4805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4807 = 9'hd9 == r_count_15_io_out ? io_r_217_b : _GEN_4806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4808 = 9'hda == r_count_15_io_out ? io_r_218_b : _GEN_4807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4809 = 9'hdb == r_count_15_io_out ? io_r_219_b : _GEN_4808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4810 = 9'hdc == r_count_15_io_out ? io_r_220_b : _GEN_4809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4811 = 9'hdd == r_count_15_io_out ? io_r_221_b : _GEN_4810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4812 = 9'hde == r_count_15_io_out ? io_r_222_b : _GEN_4811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4813 = 9'hdf == r_count_15_io_out ? io_r_223_b : _GEN_4812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4814 = 9'he0 == r_count_15_io_out ? io_r_224_b : _GEN_4813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4815 = 9'he1 == r_count_15_io_out ? io_r_225_b : _GEN_4814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4816 = 9'he2 == r_count_15_io_out ? io_r_226_b : _GEN_4815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4817 = 9'he3 == r_count_15_io_out ? io_r_227_b : _GEN_4816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4818 = 9'he4 == r_count_15_io_out ? io_r_228_b : _GEN_4817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4819 = 9'he5 == r_count_15_io_out ? io_r_229_b : _GEN_4818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4820 = 9'he6 == r_count_15_io_out ? io_r_230_b : _GEN_4819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4821 = 9'he7 == r_count_15_io_out ? io_r_231_b : _GEN_4820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4822 = 9'he8 == r_count_15_io_out ? io_r_232_b : _GEN_4821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4823 = 9'he9 == r_count_15_io_out ? io_r_233_b : _GEN_4822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4824 = 9'hea == r_count_15_io_out ? io_r_234_b : _GEN_4823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4825 = 9'heb == r_count_15_io_out ? io_r_235_b : _GEN_4824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4826 = 9'hec == r_count_15_io_out ? io_r_236_b : _GEN_4825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4827 = 9'hed == r_count_15_io_out ? io_r_237_b : _GEN_4826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4828 = 9'hee == r_count_15_io_out ? io_r_238_b : _GEN_4827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4829 = 9'hef == r_count_15_io_out ? io_r_239_b : _GEN_4828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4830 = 9'hf0 == r_count_15_io_out ? io_r_240_b : _GEN_4829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4831 = 9'hf1 == r_count_15_io_out ? io_r_241_b : _GEN_4830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4832 = 9'hf2 == r_count_15_io_out ? io_r_242_b : _GEN_4831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4833 = 9'hf3 == r_count_15_io_out ? io_r_243_b : _GEN_4832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4834 = 9'hf4 == r_count_15_io_out ? io_r_244_b : _GEN_4833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4835 = 9'hf5 == r_count_15_io_out ? io_r_245_b : _GEN_4834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4836 = 9'hf6 == r_count_15_io_out ? io_r_246_b : _GEN_4835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4837 = 9'hf7 == r_count_15_io_out ? io_r_247_b : _GEN_4836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4838 = 9'hf8 == r_count_15_io_out ? io_r_248_b : _GEN_4837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4839 = 9'hf9 == r_count_15_io_out ? io_r_249_b : _GEN_4838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4840 = 9'hfa == r_count_15_io_out ? io_r_250_b : _GEN_4839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4841 = 9'hfb == r_count_15_io_out ? io_r_251_b : _GEN_4840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4842 = 9'hfc == r_count_15_io_out ? io_r_252_b : _GEN_4841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4843 = 9'hfd == r_count_15_io_out ? io_r_253_b : _GEN_4842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4844 = 9'hfe == r_count_15_io_out ? io_r_254_b : _GEN_4843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4845 = 9'hff == r_count_15_io_out ? io_r_255_b : _GEN_4844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4846 = 9'h100 == r_count_15_io_out ? io_r_256_b : _GEN_4845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4847 = 9'h101 == r_count_15_io_out ? io_r_257_b : _GEN_4846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4848 = 9'h102 == r_count_15_io_out ? io_r_258_b : _GEN_4847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4849 = 9'h103 == r_count_15_io_out ? io_r_259_b : _GEN_4848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4850 = 9'h104 == r_count_15_io_out ? io_r_260_b : _GEN_4849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4851 = 9'h105 == r_count_15_io_out ? io_r_261_b : _GEN_4850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4852 = 9'h106 == r_count_15_io_out ? io_r_262_b : _GEN_4851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4853 = 9'h107 == r_count_15_io_out ? io_r_263_b : _GEN_4852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4854 = 9'h108 == r_count_15_io_out ? io_r_264_b : _GEN_4853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4855 = 9'h109 == r_count_15_io_out ? io_r_265_b : _GEN_4854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4856 = 9'h10a == r_count_15_io_out ? io_r_266_b : _GEN_4855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4857 = 9'h10b == r_count_15_io_out ? io_r_267_b : _GEN_4856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4858 = 9'h10c == r_count_15_io_out ? io_r_268_b : _GEN_4857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4859 = 9'h10d == r_count_15_io_out ? io_r_269_b : _GEN_4858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4860 = 9'h10e == r_count_15_io_out ? io_r_270_b : _GEN_4859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4861 = 9'h10f == r_count_15_io_out ? io_r_271_b : _GEN_4860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4862 = 9'h110 == r_count_15_io_out ? io_r_272_b : _GEN_4861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4863 = 9'h111 == r_count_15_io_out ? io_r_273_b : _GEN_4862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4864 = 9'h112 == r_count_15_io_out ? io_r_274_b : _GEN_4863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4865 = 9'h113 == r_count_15_io_out ? io_r_275_b : _GEN_4864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4866 = 9'h114 == r_count_15_io_out ? io_r_276_b : _GEN_4865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4867 = 9'h115 == r_count_15_io_out ? io_r_277_b : _GEN_4866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4868 = 9'h116 == r_count_15_io_out ? io_r_278_b : _GEN_4867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4869 = 9'h117 == r_count_15_io_out ? io_r_279_b : _GEN_4868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4870 = 9'h118 == r_count_15_io_out ? io_r_280_b : _GEN_4869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4871 = 9'h119 == r_count_15_io_out ? io_r_281_b : _GEN_4870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4872 = 9'h11a == r_count_15_io_out ? io_r_282_b : _GEN_4871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4873 = 9'h11b == r_count_15_io_out ? io_r_283_b : _GEN_4872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4874 = 9'h11c == r_count_15_io_out ? io_r_284_b : _GEN_4873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4875 = 9'h11d == r_count_15_io_out ? io_r_285_b : _GEN_4874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4876 = 9'h11e == r_count_15_io_out ? io_r_286_b : _GEN_4875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4877 = 9'h11f == r_count_15_io_out ? io_r_287_b : _GEN_4876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4878 = 9'h120 == r_count_15_io_out ? io_r_288_b : _GEN_4877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4879 = 9'h121 == r_count_15_io_out ? io_r_289_b : _GEN_4878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4880 = 9'h122 == r_count_15_io_out ? io_r_290_b : _GEN_4879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4881 = 9'h123 == r_count_15_io_out ? io_r_291_b : _GEN_4880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4882 = 9'h124 == r_count_15_io_out ? io_r_292_b : _GEN_4881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4883 = 9'h125 == r_count_15_io_out ? io_r_293_b : _GEN_4882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4884 = 9'h126 == r_count_15_io_out ? io_r_294_b : _GEN_4883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4885 = 9'h127 == r_count_15_io_out ? io_r_295_b : _GEN_4884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4886 = 9'h128 == r_count_15_io_out ? io_r_296_b : _GEN_4885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4887 = 9'h129 == r_count_15_io_out ? io_r_297_b : _GEN_4886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4888 = 9'h12a == r_count_15_io_out ? io_r_298_b : _GEN_4887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4891 = 9'h1 == r_count_16_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4892 = 9'h2 == r_count_16_io_out ? io_r_2_b : _GEN_4891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4893 = 9'h3 == r_count_16_io_out ? io_r_3_b : _GEN_4892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4894 = 9'h4 == r_count_16_io_out ? io_r_4_b : _GEN_4893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4895 = 9'h5 == r_count_16_io_out ? io_r_5_b : _GEN_4894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4896 = 9'h6 == r_count_16_io_out ? io_r_6_b : _GEN_4895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4897 = 9'h7 == r_count_16_io_out ? io_r_7_b : _GEN_4896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4898 = 9'h8 == r_count_16_io_out ? io_r_8_b : _GEN_4897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4899 = 9'h9 == r_count_16_io_out ? io_r_9_b : _GEN_4898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4900 = 9'ha == r_count_16_io_out ? io_r_10_b : _GEN_4899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4901 = 9'hb == r_count_16_io_out ? io_r_11_b : _GEN_4900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4902 = 9'hc == r_count_16_io_out ? io_r_12_b : _GEN_4901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4903 = 9'hd == r_count_16_io_out ? io_r_13_b : _GEN_4902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4904 = 9'he == r_count_16_io_out ? io_r_14_b : _GEN_4903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4905 = 9'hf == r_count_16_io_out ? io_r_15_b : _GEN_4904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4906 = 9'h10 == r_count_16_io_out ? io_r_16_b : _GEN_4905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4907 = 9'h11 == r_count_16_io_out ? io_r_17_b : _GEN_4906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4908 = 9'h12 == r_count_16_io_out ? io_r_18_b : _GEN_4907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4909 = 9'h13 == r_count_16_io_out ? io_r_19_b : _GEN_4908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4910 = 9'h14 == r_count_16_io_out ? io_r_20_b : _GEN_4909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4911 = 9'h15 == r_count_16_io_out ? io_r_21_b : _GEN_4910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4912 = 9'h16 == r_count_16_io_out ? io_r_22_b : _GEN_4911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4913 = 9'h17 == r_count_16_io_out ? io_r_23_b : _GEN_4912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4914 = 9'h18 == r_count_16_io_out ? io_r_24_b : _GEN_4913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4915 = 9'h19 == r_count_16_io_out ? io_r_25_b : _GEN_4914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4916 = 9'h1a == r_count_16_io_out ? io_r_26_b : _GEN_4915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4917 = 9'h1b == r_count_16_io_out ? io_r_27_b : _GEN_4916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4918 = 9'h1c == r_count_16_io_out ? io_r_28_b : _GEN_4917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4919 = 9'h1d == r_count_16_io_out ? io_r_29_b : _GEN_4918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4920 = 9'h1e == r_count_16_io_out ? io_r_30_b : _GEN_4919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4921 = 9'h1f == r_count_16_io_out ? io_r_31_b : _GEN_4920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4922 = 9'h20 == r_count_16_io_out ? io_r_32_b : _GEN_4921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4923 = 9'h21 == r_count_16_io_out ? io_r_33_b : _GEN_4922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4924 = 9'h22 == r_count_16_io_out ? io_r_34_b : _GEN_4923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4925 = 9'h23 == r_count_16_io_out ? io_r_35_b : _GEN_4924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4926 = 9'h24 == r_count_16_io_out ? io_r_36_b : _GEN_4925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4927 = 9'h25 == r_count_16_io_out ? io_r_37_b : _GEN_4926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4928 = 9'h26 == r_count_16_io_out ? io_r_38_b : _GEN_4927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4929 = 9'h27 == r_count_16_io_out ? io_r_39_b : _GEN_4928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4930 = 9'h28 == r_count_16_io_out ? io_r_40_b : _GEN_4929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4931 = 9'h29 == r_count_16_io_out ? io_r_41_b : _GEN_4930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4932 = 9'h2a == r_count_16_io_out ? io_r_42_b : _GEN_4931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4933 = 9'h2b == r_count_16_io_out ? io_r_43_b : _GEN_4932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4934 = 9'h2c == r_count_16_io_out ? io_r_44_b : _GEN_4933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4935 = 9'h2d == r_count_16_io_out ? io_r_45_b : _GEN_4934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4936 = 9'h2e == r_count_16_io_out ? io_r_46_b : _GEN_4935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4937 = 9'h2f == r_count_16_io_out ? io_r_47_b : _GEN_4936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4938 = 9'h30 == r_count_16_io_out ? io_r_48_b : _GEN_4937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4939 = 9'h31 == r_count_16_io_out ? io_r_49_b : _GEN_4938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4940 = 9'h32 == r_count_16_io_out ? io_r_50_b : _GEN_4939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4941 = 9'h33 == r_count_16_io_out ? io_r_51_b : _GEN_4940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4942 = 9'h34 == r_count_16_io_out ? io_r_52_b : _GEN_4941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4943 = 9'h35 == r_count_16_io_out ? io_r_53_b : _GEN_4942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4944 = 9'h36 == r_count_16_io_out ? io_r_54_b : _GEN_4943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4945 = 9'h37 == r_count_16_io_out ? io_r_55_b : _GEN_4944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4946 = 9'h38 == r_count_16_io_out ? io_r_56_b : _GEN_4945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4947 = 9'h39 == r_count_16_io_out ? io_r_57_b : _GEN_4946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4948 = 9'h3a == r_count_16_io_out ? io_r_58_b : _GEN_4947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4949 = 9'h3b == r_count_16_io_out ? io_r_59_b : _GEN_4948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4950 = 9'h3c == r_count_16_io_out ? io_r_60_b : _GEN_4949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4951 = 9'h3d == r_count_16_io_out ? io_r_61_b : _GEN_4950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4952 = 9'h3e == r_count_16_io_out ? io_r_62_b : _GEN_4951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4953 = 9'h3f == r_count_16_io_out ? io_r_63_b : _GEN_4952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4954 = 9'h40 == r_count_16_io_out ? io_r_64_b : _GEN_4953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4955 = 9'h41 == r_count_16_io_out ? io_r_65_b : _GEN_4954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4956 = 9'h42 == r_count_16_io_out ? io_r_66_b : _GEN_4955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4957 = 9'h43 == r_count_16_io_out ? io_r_67_b : _GEN_4956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4958 = 9'h44 == r_count_16_io_out ? io_r_68_b : _GEN_4957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4959 = 9'h45 == r_count_16_io_out ? io_r_69_b : _GEN_4958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4960 = 9'h46 == r_count_16_io_out ? io_r_70_b : _GEN_4959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4961 = 9'h47 == r_count_16_io_out ? io_r_71_b : _GEN_4960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4962 = 9'h48 == r_count_16_io_out ? io_r_72_b : _GEN_4961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4963 = 9'h49 == r_count_16_io_out ? io_r_73_b : _GEN_4962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4964 = 9'h4a == r_count_16_io_out ? io_r_74_b : _GEN_4963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4965 = 9'h4b == r_count_16_io_out ? io_r_75_b : _GEN_4964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4966 = 9'h4c == r_count_16_io_out ? io_r_76_b : _GEN_4965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4967 = 9'h4d == r_count_16_io_out ? io_r_77_b : _GEN_4966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4968 = 9'h4e == r_count_16_io_out ? io_r_78_b : _GEN_4967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4969 = 9'h4f == r_count_16_io_out ? io_r_79_b : _GEN_4968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4970 = 9'h50 == r_count_16_io_out ? io_r_80_b : _GEN_4969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4971 = 9'h51 == r_count_16_io_out ? io_r_81_b : _GEN_4970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4972 = 9'h52 == r_count_16_io_out ? io_r_82_b : _GEN_4971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4973 = 9'h53 == r_count_16_io_out ? io_r_83_b : _GEN_4972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4974 = 9'h54 == r_count_16_io_out ? io_r_84_b : _GEN_4973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4975 = 9'h55 == r_count_16_io_out ? io_r_85_b : _GEN_4974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4976 = 9'h56 == r_count_16_io_out ? io_r_86_b : _GEN_4975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4977 = 9'h57 == r_count_16_io_out ? io_r_87_b : _GEN_4976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4978 = 9'h58 == r_count_16_io_out ? io_r_88_b : _GEN_4977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4979 = 9'h59 == r_count_16_io_out ? io_r_89_b : _GEN_4978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4980 = 9'h5a == r_count_16_io_out ? io_r_90_b : _GEN_4979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4981 = 9'h5b == r_count_16_io_out ? io_r_91_b : _GEN_4980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4982 = 9'h5c == r_count_16_io_out ? io_r_92_b : _GEN_4981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4983 = 9'h5d == r_count_16_io_out ? io_r_93_b : _GEN_4982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4984 = 9'h5e == r_count_16_io_out ? io_r_94_b : _GEN_4983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4985 = 9'h5f == r_count_16_io_out ? io_r_95_b : _GEN_4984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4986 = 9'h60 == r_count_16_io_out ? io_r_96_b : _GEN_4985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4987 = 9'h61 == r_count_16_io_out ? io_r_97_b : _GEN_4986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4988 = 9'h62 == r_count_16_io_out ? io_r_98_b : _GEN_4987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4989 = 9'h63 == r_count_16_io_out ? io_r_99_b : _GEN_4988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4990 = 9'h64 == r_count_16_io_out ? io_r_100_b : _GEN_4989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4991 = 9'h65 == r_count_16_io_out ? io_r_101_b : _GEN_4990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4992 = 9'h66 == r_count_16_io_out ? io_r_102_b : _GEN_4991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4993 = 9'h67 == r_count_16_io_out ? io_r_103_b : _GEN_4992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4994 = 9'h68 == r_count_16_io_out ? io_r_104_b : _GEN_4993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4995 = 9'h69 == r_count_16_io_out ? io_r_105_b : _GEN_4994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4996 = 9'h6a == r_count_16_io_out ? io_r_106_b : _GEN_4995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4997 = 9'h6b == r_count_16_io_out ? io_r_107_b : _GEN_4996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4998 = 9'h6c == r_count_16_io_out ? io_r_108_b : _GEN_4997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4999 = 9'h6d == r_count_16_io_out ? io_r_109_b : _GEN_4998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5000 = 9'h6e == r_count_16_io_out ? io_r_110_b : _GEN_4999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5001 = 9'h6f == r_count_16_io_out ? io_r_111_b : _GEN_5000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5002 = 9'h70 == r_count_16_io_out ? io_r_112_b : _GEN_5001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5003 = 9'h71 == r_count_16_io_out ? io_r_113_b : _GEN_5002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5004 = 9'h72 == r_count_16_io_out ? io_r_114_b : _GEN_5003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5005 = 9'h73 == r_count_16_io_out ? io_r_115_b : _GEN_5004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5006 = 9'h74 == r_count_16_io_out ? io_r_116_b : _GEN_5005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5007 = 9'h75 == r_count_16_io_out ? io_r_117_b : _GEN_5006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5008 = 9'h76 == r_count_16_io_out ? io_r_118_b : _GEN_5007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5009 = 9'h77 == r_count_16_io_out ? io_r_119_b : _GEN_5008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5010 = 9'h78 == r_count_16_io_out ? io_r_120_b : _GEN_5009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5011 = 9'h79 == r_count_16_io_out ? io_r_121_b : _GEN_5010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5012 = 9'h7a == r_count_16_io_out ? io_r_122_b : _GEN_5011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5013 = 9'h7b == r_count_16_io_out ? io_r_123_b : _GEN_5012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5014 = 9'h7c == r_count_16_io_out ? io_r_124_b : _GEN_5013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5015 = 9'h7d == r_count_16_io_out ? io_r_125_b : _GEN_5014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5016 = 9'h7e == r_count_16_io_out ? io_r_126_b : _GEN_5015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5017 = 9'h7f == r_count_16_io_out ? io_r_127_b : _GEN_5016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5018 = 9'h80 == r_count_16_io_out ? io_r_128_b : _GEN_5017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5019 = 9'h81 == r_count_16_io_out ? io_r_129_b : _GEN_5018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5020 = 9'h82 == r_count_16_io_out ? io_r_130_b : _GEN_5019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5021 = 9'h83 == r_count_16_io_out ? io_r_131_b : _GEN_5020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5022 = 9'h84 == r_count_16_io_out ? io_r_132_b : _GEN_5021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5023 = 9'h85 == r_count_16_io_out ? io_r_133_b : _GEN_5022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5024 = 9'h86 == r_count_16_io_out ? io_r_134_b : _GEN_5023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5025 = 9'h87 == r_count_16_io_out ? io_r_135_b : _GEN_5024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5026 = 9'h88 == r_count_16_io_out ? io_r_136_b : _GEN_5025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5027 = 9'h89 == r_count_16_io_out ? io_r_137_b : _GEN_5026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5028 = 9'h8a == r_count_16_io_out ? io_r_138_b : _GEN_5027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5029 = 9'h8b == r_count_16_io_out ? io_r_139_b : _GEN_5028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5030 = 9'h8c == r_count_16_io_out ? io_r_140_b : _GEN_5029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5031 = 9'h8d == r_count_16_io_out ? io_r_141_b : _GEN_5030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5032 = 9'h8e == r_count_16_io_out ? io_r_142_b : _GEN_5031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5033 = 9'h8f == r_count_16_io_out ? io_r_143_b : _GEN_5032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5034 = 9'h90 == r_count_16_io_out ? io_r_144_b : _GEN_5033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5035 = 9'h91 == r_count_16_io_out ? io_r_145_b : _GEN_5034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5036 = 9'h92 == r_count_16_io_out ? io_r_146_b : _GEN_5035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5037 = 9'h93 == r_count_16_io_out ? io_r_147_b : _GEN_5036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5038 = 9'h94 == r_count_16_io_out ? io_r_148_b : _GEN_5037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5039 = 9'h95 == r_count_16_io_out ? io_r_149_b : _GEN_5038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5040 = 9'h96 == r_count_16_io_out ? io_r_150_b : _GEN_5039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5041 = 9'h97 == r_count_16_io_out ? io_r_151_b : _GEN_5040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5042 = 9'h98 == r_count_16_io_out ? io_r_152_b : _GEN_5041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5043 = 9'h99 == r_count_16_io_out ? io_r_153_b : _GEN_5042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5044 = 9'h9a == r_count_16_io_out ? io_r_154_b : _GEN_5043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5045 = 9'h9b == r_count_16_io_out ? io_r_155_b : _GEN_5044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5046 = 9'h9c == r_count_16_io_out ? io_r_156_b : _GEN_5045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5047 = 9'h9d == r_count_16_io_out ? io_r_157_b : _GEN_5046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5048 = 9'h9e == r_count_16_io_out ? io_r_158_b : _GEN_5047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5049 = 9'h9f == r_count_16_io_out ? io_r_159_b : _GEN_5048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5050 = 9'ha0 == r_count_16_io_out ? io_r_160_b : _GEN_5049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5051 = 9'ha1 == r_count_16_io_out ? io_r_161_b : _GEN_5050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5052 = 9'ha2 == r_count_16_io_out ? io_r_162_b : _GEN_5051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5053 = 9'ha3 == r_count_16_io_out ? io_r_163_b : _GEN_5052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5054 = 9'ha4 == r_count_16_io_out ? io_r_164_b : _GEN_5053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5055 = 9'ha5 == r_count_16_io_out ? io_r_165_b : _GEN_5054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5056 = 9'ha6 == r_count_16_io_out ? io_r_166_b : _GEN_5055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5057 = 9'ha7 == r_count_16_io_out ? io_r_167_b : _GEN_5056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5058 = 9'ha8 == r_count_16_io_out ? io_r_168_b : _GEN_5057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5059 = 9'ha9 == r_count_16_io_out ? io_r_169_b : _GEN_5058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5060 = 9'haa == r_count_16_io_out ? io_r_170_b : _GEN_5059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5061 = 9'hab == r_count_16_io_out ? io_r_171_b : _GEN_5060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5062 = 9'hac == r_count_16_io_out ? io_r_172_b : _GEN_5061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5063 = 9'had == r_count_16_io_out ? io_r_173_b : _GEN_5062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5064 = 9'hae == r_count_16_io_out ? io_r_174_b : _GEN_5063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5065 = 9'haf == r_count_16_io_out ? io_r_175_b : _GEN_5064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5066 = 9'hb0 == r_count_16_io_out ? io_r_176_b : _GEN_5065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5067 = 9'hb1 == r_count_16_io_out ? io_r_177_b : _GEN_5066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5068 = 9'hb2 == r_count_16_io_out ? io_r_178_b : _GEN_5067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5069 = 9'hb3 == r_count_16_io_out ? io_r_179_b : _GEN_5068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5070 = 9'hb4 == r_count_16_io_out ? io_r_180_b : _GEN_5069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5071 = 9'hb5 == r_count_16_io_out ? io_r_181_b : _GEN_5070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5072 = 9'hb6 == r_count_16_io_out ? io_r_182_b : _GEN_5071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5073 = 9'hb7 == r_count_16_io_out ? io_r_183_b : _GEN_5072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5074 = 9'hb8 == r_count_16_io_out ? io_r_184_b : _GEN_5073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5075 = 9'hb9 == r_count_16_io_out ? io_r_185_b : _GEN_5074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5076 = 9'hba == r_count_16_io_out ? io_r_186_b : _GEN_5075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5077 = 9'hbb == r_count_16_io_out ? io_r_187_b : _GEN_5076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5078 = 9'hbc == r_count_16_io_out ? io_r_188_b : _GEN_5077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5079 = 9'hbd == r_count_16_io_out ? io_r_189_b : _GEN_5078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5080 = 9'hbe == r_count_16_io_out ? io_r_190_b : _GEN_5079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5081 = 9'hbf == r_count_16_io_out ? io_r_191_b : _GEN_5080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5082 = 9'hc0 == r_count_16_io_out ? io_r_192_b : _GEN_5081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5083 = 9'hc1 == r_count_16_io_out ? io_r_193_b : _GEN_5082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5084 = 9'hc2 == r_count_16_io_out ? io_r_194_b : _GEN_5083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5085 = 9'hc3 == r_count_16_io_out ? io_r_195_b : _GEN_5084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5086 = 9'hc4 == r_count_16_io_out ? io_r_196_b : _GEN_5085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5087 = 9'hc5 == r_count_16_io_out ? io_r_197_b : _GEN_5086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5088 = 9'hc6 == r_count_16_io_out ? io_r_198_b : _GEN_5087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5089 = 9'hc7 == r_count_16_io_out ? io_r_199_b : _GEN_5088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5090 = 9'hc8 == r_count_16_io_out ? io_r_200_b : _GEN_5089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5091 = 9'hc9 == r_count_16_io_out ? io_r_201_b : _GEN_5090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5092 = 9'hca == r_count_16_io_out ? io_r_202_b : _GEN_5091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5093 = 9'hcb == r_count_16_io_out ? io_r_203_b : _GEN_5092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5094 = 9'hcc == r_count_16_io_out ? io_r_204_b : _GEN_5093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5095 = 9'hcd == r_count_16_io_out ? io_r_205_b : _GEN_5094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5096 = 9'hce == r_count_16_io_out ? io_r_206_b : _GEN_5095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5097 = 9'hcf == r_count_16_io_out ? io_r_207_b : _GEN_5096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5098 = 9'hd0 == r_count_16_io_out ? io_r_208_b : _GEN_5097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5099 = 9'hd1 == r_count_16_io_out ? io_r_209_b : _GEN_5098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5100 = 9'hd2 == r_count_16_io_out ? io_r_210_b : _GEN_5099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5101 = 9'hd3 == r_count_16_io_out ? io_r_211_b : _GEN_5100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5102 = 9'hd4 == r_count_16_io_out ? io_r_212_b : _GEN_5101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5103 = 9'hd5 == r_count_16_io_out ? io_r_213_b : _GEN_5102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5104 = 9'hd6 == r_count_16_io_out ? io_r_214_b : _GEN_5103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5105 = 9'hd7 == r_count_16_io_out ? io_r_215_b : _GEN_5104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5106 = 9'hd8 == r_count_16_io_out ? io_r_216_b : _GEN_5105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5107 = 9'hd9 == r_count_16_io_out ? io_r_217_b : _GEN_5106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5108 = 9'hda == r_count_16_io_out ? io_r_218_b : _GEN_5107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5109 = 9'hdb == r_count_16_io_out ? io_r_219_b : _GEN_5108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5110 = 9'hdc == r_count_16_io_out ? io_r_220_b : _GEN_5109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5111 = 9'hdd == r_count_16_io_out ? io_r_221_b : _GEN_5110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5112 = 9'hde == r_count_16_io_out ? io_r_222_b : _GEN_5111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5113 = 9'hdf == r_count_16_io_out ? io_r_223_b : _GEN_5112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5114 = 9'he0 == r_count_16_io_out ? io_r_224_b : _GEN_5113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5115 = 9'he1 == r_count_16_io_out ? io_r_225_b : _GEN_5114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5116 = 9'he2 == r_count_16_io_out ? io_r_226_b : _GEN_5115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5117 = 9'he3 == r_count_16_io_out ? io_r_227_b : _GEN_5116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5118 = 9'he4 == r_count_16_io_out ? io_r_228_b : _GEN_5117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5119 = 9'he5 == r_count_16_io_out ? io_r_229_b : _GEN_5118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5120 = 9'he6 == r_count_16_io_out ? io_r_230_b : _GEN_5119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5121 = 9'he7 == r_count_16_io_out ? io_r_231_b : _GEN_5120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5122 = 9'he8 == r_count_16_io_out ? io_r_232_b : _GEN_5121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5123 = 9'he9 == r_count_16_io_out ? io_r_233_b : _GEN_5122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5124 = 9'hea == r_count_16_io_out ? io_r_234_b : _GEN_5123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5125 = 9'heb == r_count_16_io_out ? io_r_235_b : _GEN_5124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5126 = 9'hec == r_count_16_io_out ? io_r_236_b : _GEN_5125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5127 = 9'hed == r_count_16_io_out ? io_r_237_b : _GEN_5126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5128 = 9'hee == r_count_16_io_out ? io_r_238_b : _GEN_5127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5129 = 9'hef == r_count_16_io_out ? io_r_239_b : _GEN_5128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5130 = 9'hf0 == r_count_16_io_out ? io_r_240_b : _GEN_5129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5131 = 9'hf1 == r_count_16_io_out ? io_r_241_b : _GEN_5130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5132 = 9'hf2 == r_count_16_io_out ? io_r_242_b : _GEN_5131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5133 = 9'hf3 == r_count_16_io_out ? io_r_243_b : _GEN_5132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5134 = 9'hf4 == r_count_16_io_out ? io_r_244_b : _GEN_5133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5135 = 9'hf5 == r_count_16_io_out ? io_r_245_b : _GEN_5134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5136 = 9'hf6 == r_count_16_io_out ? io_r_246_b : _GEN_5135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5137 = 9'hf7 == r_count_16_io_out ? io_r_247_b : _GEN_5136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5138 = 9'hf8 == r_count_16_io_out ? io_r_248_b : _GEN_5137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5139 = 9'hf9 == r_count_16_io_out ? io_r_249_b : _GEN_5138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5140 = 9'hfa == r_count_16_io_out ? io_r_250_b : _GEN_5139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5141 = 9'hfb == r_count_16_io_out ? io_r_251_b : _GEN_5140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5142 = 9'hfc == r_count_16_io_out ? io_r_252_b : _GEN_5141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5143 = 9'hfd == r_count_16_io_out ? io_r_253_b : _GEN_5142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5144 = 9'hfe == r_count_16_io_out ? io_r_254_b : _GEN_5143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5145 = 9'hff == r_count_16_io_out ? io_r_255_b : _GEN_5144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5146 = 9'h100 == r_count_16_io_out ? io_r_256_b : _GEN_5145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5147 = 9'h101 == r_count_16_io_out ? io_r_257_b : _GEN_5146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5148 = 9'h102 == r_count_16_io_out ? io_r_258_b : _GEN_5147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5149 = 9'h103 == r_count_16_io_out ? io_r_259_b : _GEN_5148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5150 = 9'h104 == r_count_16_io_out ? io_r_260_b : _GEN_5149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5151 = 9'h105 == r_count_16_io_out ? io_r_261_b : _GEN_5150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5152 = 9'h106 == r_count_16_io_out ? io_r_262_b : _GEN_5151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5153 = 9'h107 == r_count_16_io_out ? io_r_263_b : _GEN_5152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5154 = 9'h108 == r_count_16_io_out ? io_r_264_b : _GEN_5153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5155 = 9'h109 == r_count_16_io_out ? io_r_265_b : _GEN_5154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5156 = 9'h10a == r_count_16_io_out ? io_r_266_b : _GEN_5155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5157 = 9'h10b == r_count_16_io_out ? io_r_267_b : _GEN_5156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5158 = 9'h10c == r_count_16_io_out ? io_r_268_b : _GEN_5157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5159 = 9'h10d == r_count_16_io_out ? io_r_269_b : _GEN_5158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5160 = 9'h10e == r_count_16_io_out ? io_r_270_b : _GEN_5159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5161 = 9'h10f == r_count_16_io_out ? io_r_271_b : _GEN_5160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5162 = 9'h110 == r_count_16_io_out ? io_r_272_b : _GEN_5161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5163 = 9'h111 == r_count_16_io_out ? io_r_273_b : _GEN_5162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5164 = 9'h112 == r_count_16_io_out ? io_r_274_b : _GEN_5163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5165 = 9'h113 == r_count_16_io_out ? io_r_275_b : _GEN_5164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5166 = 9'h114 == r_count_16_io_out ? io_r_276_b : _GEN_5165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5167 = 9'h115 == r_count_16_io_out ? io_r_277_b : _GEN_5166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5168 = 9'h116 == r_count_16_io_out ? io_r_278_b : _GEN_5167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5169 = 9'h117 == r_count_16_io_out ? io_r_279_b : _GEN_5168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5170 = 9'h118 == r_count_16_io_out ? io_r_280_b : _GEN_5169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5171 = 9'h119 == r_count_16_io_out ? io_r_281_b : _GEN_5170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5172 = 9'h11a == r_count_16_io_out ? io_r_282_b : _GEN_5171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5173 = 9'h11b == r_count_16_io_out ? io_r_283_b : _GEN_5172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5174 = 9'h11c == r_count_16_io_out ? io_r_284_b : _GEN_5173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5175 = 9'h11d == r_count_16_io_out ? io_r_285_b : _GEN_5174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5176 = 9'h11e == r_count_16_io_out ? io_r_286_b : _GEN_5175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5177 = 9'h11f == r_count_16_io_out ? io_r_287_b : _GEN_5176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5178 = 9'h120 == r_count_16_io_out ? io_r_288_b : _GEN_5177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5179 = 9'h121 == r_count_16_io_out ? io_r_289_b : _GEN_5178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5180 = 9'h122 == r_count_16_io_out ? io_r_290_b : _GEN_5179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5181 = 9'h123 == r_count_16_io_out ? io_r_291_b : _GEN_5180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5182 = 9'h124 == r_count_16_io_out ? io_r_292_b : _GEN_5181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5183 = 9'h125 == r_count_16_io_out ? io_r_293_b : _GEN_5182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5184 = 9'h126 == r_count_16_io_out ? io_r_294_b : _GEN_5183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5185 = 9'h127 == r_count_16_io_out ? io_r_295_b : _GEN_5184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5186 = 9'h128 == r_count_16_io_out ? io_r_296_b : _GEN_5185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5187 = 9'h129 == r_count_16_io_out ? io_r_297_b : _GEN_5186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5188 = 9'h12a == r_count_16_io_out ? io_r_298_b : _GEN_5187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5191 = 9'h1 == r_count_17_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5192 = 9'h2 == r_count_17_io_out ? io_r_2_b : _GEN_5191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5193 = 9'h3 == r_count_17_io_out ? io_r_3_b : _GEN_5192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5194 = 9'h4 == r_count_17_io_out ? io_r_4_b : _GEN_5193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5195 = 9'h5 == r_count_17_io_out ? io_r_5_b : _GEN_5194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5196 = 9'h6 == r_count_17_io_out ? io_r_6_b : _GEN_5195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5197 = 9'h7 == r_count_17_io_out ? io_r_7_b : _GEN_5196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5198 = 9'h8 == r_count_17_io_out ? io_r_8_b : _GEN_5197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5199 = 9'h9 == r_count_17_io_out ? io_r_9_b : _GEN_5198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5200 = 9'ha == r_count_17_io_out ? io_r_10_b : _GEN_5199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5201 = 9'hb == r_count_17_io_out ? io_r_11_b : _GEN_5200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5202 = 9'hc == r_count_17_io_out ? io_r_12_b : _GEN_5201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5203 = 9'hd == r_count_17_io_out ? io_r_13_b : _GEN_5202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5204 = 9'he == r_count_17_io_out ? io_r_14_b : _GEN_5203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5205 = 9'hf == r_count_17_io_out ? io_r_15_b : _GEN_5204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5206 = 9'h10 == r_count_17_io_out ? io_r_16_b : _GEN_5205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5207 = 9'h11 == r_count_17_io_out ? io_r_17_b : _GEN_5206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5208 = 9'h12 == r_count_17_io_out ? io_r_18_b : _GEN_5207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5209 = 9'h13 == r_count_17_io_out ? io_r_19_b : _GEN_5208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5210 = 9'h14 == r_count_17_io_out ? io_r_20_b : _GEN_5209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5211 = 9'h15 == r_count_17_io_out ? io_r_21_b : _GEN_5210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5212 = 9'h16 == r_count_17_io_out ? io_r_22_b : _GEN_5211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5213 = 9'h17 == r_count_17_io_out ? io_r_23_b : _GEN_5212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5214 = 9'h18 == r_count_17_io_out ? io_r_24_b : _GEN_5213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5215 = 9'h19 == r_count_17_io_out ? io_r_25_b : _GEN_5214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5216 = 9'h1a == r_count_17_io_out ? io_r_26_b : _GEN_5215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5217 = 9'h1b == r_count_17_io_out ? io_r_27_b : _GEN_5216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5218 = 9'h1c == r_count_17_io_out ? io_r_28_b : _GEN_5217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5219 = 9'h1d == r_count_17_io_out ? io_r_29_b : _GEN_5218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5220 = 9'h1e == r_count_17_io_out ? io_r_30_b : _GEN_5219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5221 = 9'h1f == r_count_17_io_out ? io_r_31_b : _GEN_5220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5222 = 9'h20 == r_count_17_io_out ? io_r_32_b : _GEN_5221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5223 = 9'h21 == r_count_17_io_out ? io_r_33_b : _GEN_5222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5224 = 9'h22 == r_count_17_io_out ? io_r_34_b : _GEN_5223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5225 = 9'h23 == r_count_17_io_out ? io_r_35_b : _GEN_5224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5226 = 9'h24 == r_count_17_io_out ? io_r_36_b : _GEN_5225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5227 = 9'h25 == r_count_17_io_out ? io_r_37_b : _GEN_5226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5228 = 9'h26 == r_count_17_io_out ? io_r_38_b : _GEN_5227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5229 = 9'h27 == r_count_17_io_out ? io_r_39_b : _GEN_5228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5230 = 9'h28 == r_count_17_io_out ? io_r_40_b : _GEN_5229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5231 = 9'h29 == r_count_17_io_out ? io_r_41_b : _GEN_5230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5232 = 9'h2a == r_count_17_io_out ? io_r_42_b : _GEN_5231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5233 = 9'h2b == r_count_17_io_out ? io_r_43_b : _GEN_5232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5234 = 9'h2c == r_count_17_io_out ? io_r_44_b : _GEN_5233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5235 = 9'h2d == r_count_17_io_out ? io_r_45_b : _GEN_5234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5236 = 9'h2e == r_count_17_io_out ? io_r_46_b : _GEN_5235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5237 = 9'h2f == r_count_17_io_out ? io_r_47_b : _GEN_5236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5238 = 9'h30 == r_count_17_io_out ? io_r_48_b : _GEN_5237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5239 = 9'h31 == r_count_17_io_out ? io_r_49_b : _GEN_5238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5240 = 9'h32 == r_count_17_io_out ? io_r_50_b : _GEN_5239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5241 = 9'h33 == r_count_17_io_out ? io_r_51_b : _GEN_5240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5242 = 9'h34 == r_count_17_io_out ? io_r_52_b : _GEN_5241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5243 = 9'h35 == r_count_17_io_out ? io_r_53_b : _GEN_5242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5244 = 9'h36 == r_count_17_io_out ? io_r_54_b : _GEN_5243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5245 = 9'h37 == r_count_17_io_out ? io_r_55_b : _GEN_5244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5246 = 9'h38 == r_count_17_io_out ? io_r_56_b : _GEN_5245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5247 = 9'h39 == r_count_17_io_out ? io_r_57_b : _GEN_5246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5248 = 9'h3a == r_count_17_io_out ? io_r_58_b : _GEN_5247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5249 = 9'h3b == r_count_17_io_out ? io_r_59_b : _GEN_5248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5250 = 9'h3c == r_count_17_io_out ? io_r_60_b : _GEN_5249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5251 = 9'h3d == r_count_17_io_out ? io_r_61_b : _GEN_5250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5252 = 9'h3e == r_count_17_io_out ? io_r_62_b : _GEN_5251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5253 = 9'h3f == r_count_17_io_out ? io_r_63_b : _GEN_5252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5254 = 9'h40 == r_count_17_io_out ? io_r_64_b : _GEN_5253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5255 = 9'h41 == r_count_17_io_out ? io_r_65_b : _GEN_5254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5256 = 9'h42 == r_count_17_io_out ? io_r_66_b : _GEN_5255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5257 = 9'h43 == r_count_17_io_out ? io_r_67_b : _GEN_5256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5258 = 9'h44 == r_count_17_io_out ? io_r_68_b : _GEN_5257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5259 = 9'h45 == r_count_17_io_out ? io_r_69_b : _GEN_5258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5260 = 9'h46 == r_count_17_io_out ? io_r_70_b : _GEN_5259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5261 = 9'h47 == r_count_17_io_out ? io_r_71_b : _GEN_5260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5262 = 9'h48 == r_count_17_io_out ? io_r_72_b : _GEN_5261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5263 = 9'h49 == r_count_17_io_out ? io_r_73_b : _GEN_5262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5264 = 9'h4a == r_count_17_io_out ? io_r_74_b : _GEN_5263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5265 = 9'h4b == r_count_17_io_out ? io_r_75_b : _GEN_5264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5266 = 9'h4c == r_count_17_io_out ? io_r_76_b : _GEN_5265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5267 = 9'h4d == r_count_17_io_out ? io_r_77_b : _GEN_5266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5268 = 9'h4e == r_count_17_io_out ? io_r_78_b : _GEN_5267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5269 = 9'h4f == r_count_17_io_out ? io_r_79_b : _GEN_5268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5270 = 9'h50 == r_count_17_io_out ? io_r_80_b : _GEN_5269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5271 = 9'h51 == r_count_17_io_out ? io_r_81_b : _GEN_5270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5272 = 9'h52 == r_count_17_io_out ? io_r_82_b : _GEN_5271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5273 = 9'h53 == r_count_17_io_out ? io_r_83_b : _GEN_5272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5274 = 9'h54 == r_count_17_io_out ? io_r_84_b : _GEN_5273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5275 = 9'h55 == r_count_17_io_out ? io_r_85_b : _GEN_5274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5276 = 9'h56 == r_count_17_io_out ? io_r_86_b : _GEN_5275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5277 = 9'h57 == r_count_17_io_out ? io_r_87_b : _GEN_5276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5278 = 9'h58 == r_count_17_io_out ? io_r_88_b : _GEN_5277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5279 = 9'h59 == r_count_17_io_out ? io_r_89_b : _GEN_5278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5280 = 9'h5a == r_count_17_io_out ? io_r_90_b : _GEN_5279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5281 = 9'h5b == r_count_17_io_out ? io_r_91_b : _GEN_5280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5282 = 9'h5c == r_count_17_io_out ? io_r_92_b : _GEN_5281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5283 = 9'h5d == r_count_17_io_out ? io_r_93_b : _GEN_5282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5284 = 9'h5e == r_count_17_io_out ? io_r_94_b : _GEN_5283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5285 = 9'h5f == r_count_17_io_out ? io_r_95_b : _GEN_5284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5286 = 9'h60 == r_count_17_io_out ? io_r_96_b : _GEN_5285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5287 = 9'h61 == r_count_17_io_out ? io_r_97_b : _GEN_5286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5288 = 9'h62 == r_count_17_io_out ? io_r_98_b : _GEN_5287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5289 = 9'h63 == r_count_17_io_out ? io_r_99_b : _GEN_5288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5290 = 9'h64 == r_count_17_io_out ? io_r_100_b : _GEN_5289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5291 = 9'h65 == r_count_17_io_out ? io_r_101_b : _GEN_5290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5292 = 9'h66 == r_count_17_io_out ? io_r_102_b : _GEN_5291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5293 = 9'h67 == r_count_17_io_out ? io_r_103_b : _GEN_5292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5294 = 9'h68 == r_count_17_io_out ? io_r_104_b : _GEN_5293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5295 = 9'h69 == r_count_17_io_out ? io_r_105_b : _GEN_5294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5296 = 9'h6a == r_count_17_io_out ? io_r_106_b : _GEN_5295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5297 = 9'h6b == r_count_17_io_out ? io_r_107_b : _GEN_5296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5298 = 9'h6c == r_count_17_io_out ? io_r_108_b : _GEN_5297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5299 = 9'h6d == r_count_17_io_out ? io_r_109_b : _GEN_5298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5300 = 9'h6e == r_count_17_io_out ? io_r_110_b : _GEN_5299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5301 = 9'h6f == r_count_17_io_out ? io_r_111_b : _GEN_5300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5302 = 9'h70 == r_count_17_io_out ? io_r_112_b : _GEN_5301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5303 = 9'h71 == r_count_17_io_out ? io_r_113_b : _GEN_5302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5304 = 9'h72 == r_count_17_io_out ? io_r_114_b : _GEN_5303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5305 = 9'h73 == r_count_17_io_out ? io_r_115_b : _GEN_5304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5306 = 9'h74 == r_count_17_io_out ? io_r_116_b : _GEN_5305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5307 = 9'h75 == r_count_17_io_out ? io_r_117_b : _GEN_5306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5308 = 9'h76 == r_count_17_io_out ? io_r_118_b : _GEN_5307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5309 = 9'h77 == r_count_17_io_out ? io_r_119_b : _GEN_5308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5310 = 9'h78 == r_count_17_io_out ? io_r_120_b : _GEN_5309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5311 = 9'h79 == r_count_17_io_out ? io_r_121_b : _GEN_5310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5312 = 9'h7a == r_count_17_io_out ? io_r_122_b : _GEN_5311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5313 = 9'h7b == r_count_17_io_out ? io_r_123_b : _GEN_5312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5314 = 9'h7c == r_count_17_io_out ? io_r_124_b : _GEN_5313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5315 = 9'h7d == r_count_17_io_out ? io_r_125_b : _GEN_5314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5316 = 9'h7e == r_count_17_io_out ? io_r_126_b : _GEN_5315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5317 = 9'h7f == r_count_17_io_out ? io_r_127_b : _GEN_5316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5318 = 9'h80 == r_count_17_io_out ? io_r_128_b : _GEN_5317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5319 = 9'h81 == r_count_17_io_out ? io_r_129_b : _GEN_5318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5320 = 9'h82 == r_count_17_io_out ? io_r_130_b : _GEN_5319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5321 = 9'h83 == r_count_17_io_out ? io_r_131_b : _GEN_5320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5322 = 9'h84 == r_count_17_io_out ? io_r_132_b : _GEN_5321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5323 = 9'h85 == r_count_17_io_out ? io_r_133_b : _GEN_5322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5324 = 9'h86 == r_count_17_io_out ? io_r_134_b : _GEN_5323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5325 = 9'h87 == r_count_17_io_out ? io_r_135_b : _GEN_5324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5326 = 9'h88 == r_count_17_io_out ? io_r_136_b : _GEN_5325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5327 = 9'h89 == r_count_17_io_out ? io_r_137_b : _GEN_5326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5328 = 9'h8a == r_count_17_io_out ? io_r_138_b : _GEN_5327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5329 = 9'h8b == r_count_17_io_out ? io_r_139_b : _GEN_5328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5330 = 9'h8c == r_count_17_io_out ? io_r_140_b : _GEN_5329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5331 = 9'h8d == r_count_17_io_out ? io_r_141_b : _GEN_5330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5332 = 9'h8e == r_count_17_io_out ? io_r_142_b : _GEN_5331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5333 = 9'h8f == r_count_17_io_out ? io_r_143_b : _GEN_5332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5334 = 9'h90 == r_count_17_io_out ? io_r_144_b : _GEN_5333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5335 = 9'h91 == r_count_17_io_out ? io_r_145_b : _GEN_5334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5336 = 9'h92 == r_count_17_io_out ? io_r_146_b : _GEN_5335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5337 = 9'h93 == r_count_17_io_out ? io_r_147_b : _GEN_5336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5338 = 9'h94 == r_count_17_io_out ? io_r_148_b : _GEN_5337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5339 = 9'h95 == r_count_17_io_out ? io_r_149_b : _GEN_5338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5340 = 9'h96 == r_count_17_io_out ? io_r_150_b : _GEN_5339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5341 = 9'h97 == r_count_17_io_out ? io_r_151_b : _GEN_5340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5342 = 9'h98 == r_count_17_io_out ? io_r_152_b : _GEN_5341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5343 = 9'h99 == r_count_17_io_out ? io_r_153_b : _GEN_5342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5344 = 9'h9a == r_count_17_io_out ? io_r_154_b : _GEN_5343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5345 = 9'h9b == r_count_17_io_out ? io_r_155_b : _GEN_5344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5346 = 9'h9c == r_count_17_io_out ? io_r_156_b : _GEN_5345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5347 = 9'h9d == r_count_17_io_out ? io_r_157_b : _GEN_5346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5348 = 9'h9e == r_count_17_io_out ? io_r_158_b : _GEN_5347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5349 = 9'h9f == r_count_17_io_out ? io_r_159_b : _GEN_5348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5350 = 9'ha0 == r_count_17_io_out ? io_r_160_b : _GEN_5349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5351 = 9'ha1 == r_count_17_io_out ? io_r_161_b : _GEN_5350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5352 = 9'ha2 == r_count_17_io_out ? io_r_162_b : _GEN_5351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5353 = 9'ha3 == r_count_17_io_out ? io_r_163_b : _GEN_5352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5354 = 9'ha4 == r_count_17_io_out ? io_r_164_b : _GEN_5353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5355 = 9'ha5 == r_count_17_io_out ? io_r_165_b : _GEN_5354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5356 = 9'ha6 == r_count_17_io_out ? io_r_166_b : _GEN_5355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5357 = 9'ha7 == r_count_17_io_out ? io_r_167_b : _GEN_5356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5358 = 9'ha8 == r_count_17_io_out ? io_r_168_b : _GEN_5357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5359 = 9'ha9 == r_count_17_io_out ? io_r_169_b : _GEN_5358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5360 = 9'haa == r_count_17_io_out ? io_r_170_b : _GEN_5359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5361 = 9'hab == r_count_17_io_out ? io_r_171_b : _GEN_5360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5362 = 9'hac == r_count_17_io_out ? io_r_172_b : _GEN_5361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5363 = 9'had == r_count_17_io_out ? io_r_173_b : _GEN_5362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5364 = 9'hae == r_count_17_io_out ? io_r_174_b : _GEN_5363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5365 = 9'haf == r_count_17_io_out ? io_r_175_b : _GEN_5364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5366 = 9'hb0 == r_count_17_io_out ? io_r_176_b : _GEN_5365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5367 = 9'hb1 == r_count_17_io_out ? io_r_177_b : _GEN_5366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5368 = 9'hb2 == r_count_17_io_out ? io_r_178_b : _GEN_5367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5369 = 9'hb3 == r_count_17_io_out ? io_r_179_b : _GEN_5368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5370 = 9'hb4 == r_count_17_io_out ? io_r_180_b : _GEN_5369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5371 = 9'hb5 == r_count_17_io_out ? io_r_181_b : _GEN_5370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5372 = 9'hb6 == r_count_17_io_out ? io_r_182_b : _GEN_5371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5373 = 9'hb7 == r_count_17_io_out ? io_r_183_b : _GEN_5372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5374 = 9'hb8 == r_count_17_io_out ? io_r_184_b : _GEN_5373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5375 = 9'hb9 == r_count_17_io_out ? io_r_185_b : _GEN_5374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5376 = 9'hba == r_count_17_io_out ? io_r_186_b : _GEN_5375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5377 = 9'hbb == r_count_17_io_out ? io_r_187_b : _GEN_5376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5378 = 9'hbc == r_count_17_io_out ? io_r_188_b : _GEN_5377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5379 = 9'hbd == r_count_17_io_out ? io_r_189_b : _GEN_5378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5380 = 9'hbe == r_count_17_io_out ? io_r_190_b : _GEN_5379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5381 = 9'hbf == r_count_17_io_out ? io_r_191_b : _GEN_5380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5382 = 9'hc0 == r_count_17_io_out ? io_r_192_b : _GEN_5381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5383 = 9'hc1 == r_count_17_io_out ? io_r_193_b : _GEN_5382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5384 = 9'hc2 == r_count_17_io_out ? io_r_194_b : _GEN_5383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5385 = 9'hc3 == r_count_17_io_out ? io_r_195_b : _GEN_5384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5386 = 9'hc4 == r_count_17_io_out ? io_r_196_b : _GEN_5385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5387 = 9'hc5 == r_count_17_io_out ? io_r_197_b : _GEN_5386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5388 = 9'hc6 == r_count_17_io_out ? io_r_198_b : _GEN_5387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5389 = 9'hc7 == r_count_17_io_out ? io_r_199_b : _GEN_5388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5390 = 9'hc8 == r_count_17_io_out ? io_r_200_b : _GEN_5389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5391 = 9'hc9 == r_count_17_io_out ? io_r_201_b : _GEN_5390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5392 = 9'hca == r_count_17_io_out ? io_r_202_b : _GEN_5391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5393 = 9'hcb == r_count_17_io_out ? io_r_203_b : _GEN_5392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5394 = 9'hcc == r_count_17_io_out ? io_r_204_b : _GEN_5393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5395 = 9'hcd == r_count_17_io_out ? io_r_205_b : _GEN_5394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5396 = 9'hce == r_count_17_io_out ? io_r_206_b : _GEN_5395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5397 = 9'hcf == r_count_17_io_out ? io_r_207_b : _GEN_5396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5398 = 9'hd0 == r_count_17_io_out ? io_r_208_b : _GEN_5397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5399 = 9'hd1 == r_count_17_io_out ? io_r_209_b : _GEN_5398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5400 = 9'hd2 == r_count_17_io_out ? io_r_210_b : _GEN_5399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5401 = 9'hd3 == r_count_17_io_out ? io_r_211_b : _GEN_5400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5402 = 9'hd4 == r_count_17_io_out ? io_r_212_b : _GEN_5401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5403 = 9'hd5 == r_count_17_io_out ? io_r_213_b : _GEN_5402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5404 = 9'hd6 == r_count_17_io_out ? io_r_214_b : _GEN_5403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5405 = 9'hd7 == r_count_17_io_out ? io_r_215_b : _GEN_5404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5406 = 9'hd8 == r_count_17_io_out ? io_r_216_b : _GEN_5405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5407 = 9'hd9 == r_count_17_io_out ? io_r_217_b : _GEN_5406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5408 = 9'hda == r_count_17_io_out ? io_r_218_b : _GEN_5407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5409 = 9'hdb == r_count_17_io_out ? io_r_219_b : _GEN_5408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5410 = 9'hdc == r_count_17_io_out ? io_r_220_b : _GEN_5409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5411 = 9'hdd == r_count_17_io_out ? io_r_221_b : _GEN_5410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5412 = 9'hde == r_count_17_io_out ? io_r_222_b : _GEN_5411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5413 = 9'hdf == r_count_17_io_out ? io_r_223_b : _GEN_5412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5414 = 9'he0 == r_count_17_io_out ? io_r_224_b : _GEN_5413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5415 = 9'he1 == r_count_17_io_out ? io_r_225_b : _GEN_5414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5416 = 9'he2 == r_count_17_io_out ? io_r_226_b : _GEN_5415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5417 = 9'he3 == r_count_17_io_out ? io_r_227_b : _GEN_5416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5418 = 9'he4 == r_count_17_io_out ? io_r_228_b : _GEN_5417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5419 = 9'he5 == r_count_17_io_out ? io_r_229_b : _GEN_5418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5420 = 9'he6 == r_count_17_io_out ? io_r_230_b : _GEN_5419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5421 = 9'he7 == r_count_17_io_out ? io_r_231_b : _GEN_5420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5422 = 9'he8 == r_count_17_io_out ? io_r_232_b : _GEN_5421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5423 = 9'he9 == r_count_17_io_out ? io_r_233_b : _GEN_5422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5424 = 9'hea == r_count_17_io_out ? io_r_234_b : _GEN_5423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5425 = 9'heb == r_count_17_io_out ? io_r_235_b : _GEN_5424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5426 = 9'hec == r_count_17_io_out ? io_r_236_b : _GEN_5425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5427 = 9'hed == r_count_17_io_out ? io_r_237_b : _GEN_5426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5428 = 9'hee == r_count_17_io_out ? io_r_238_b : _GEN_5427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5429 = 9'hef == r_count_17_io_out ? io_r_239_b : _GEN_5428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5430 = 9'hf0 == r_count_17_io_out ? io_r_240_b : _GEN_5429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5431 = 9'hf1 == r_count_17_io_out ? io_r_241_b : _GEN_5430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5432 = 9'hf2 == r_count_17_io_out ? io_r_242_b : _GEN_5431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5433 = 9'hf3 == r_count_17_io_out ? io_r_243_b : _GEN_5432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5434 = 9'hf4 == r_count_17_io_out ? io_r_244_b : _GEN_5433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5435 = 9'hf5 == r_count_17_io_out ? io_r_245_b : _GEN_5434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5436 = 9'hf6 == r_count_17_io_out ? io_r_246_b : _GEN_5435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5437 = 9'hf7 == r_count_17_io_out ? io_r_247_b : _GEN_5436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5438 = 9'hf8 == r_count_17_io_out ? io_r_248_b : _GEN_5437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5439 = 9'hf9 == r_count_17_io_out ? io_r_249_b : _GEN_5438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5440 = 9'hfa == r_count_17_io_out ? io_r_250_b : _GEN_5439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5441 = 9'hfb == r_count_17_io_out ? io_r_251_b : _GEN_5440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5442 = 9'hfc == r_count_17_io_out ? io_r_252_b : _GEN_5441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5443 = 9'hfd == r_count_17_io_out ? io_r_253_b : _GEN_5442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5444 = 9'hfe == r_count_17_io_out ? io_r_254_b : _GEN_5443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5445 = 9'hff == r_count_17_io_out ? io_r_255_b : _GEN_5444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5446 = 9'h100 == r_count_17_io_out ? io_r_256_b : _GEN_5445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5447 = 9'h101 == r_count_17_io_out ? io_r_257_b : _GEN_5446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5448 = 9'h102 == r_count_17_io_out ? io_r_258_b : _GEN_5447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5449 = 9'h103 == r_count_17_io_out ? io_r_259_b : _GEN_5448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5450 = 9'h104 == r_count_17_io_out ? io_r_260_b : _GEN_5449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5451 = 9'h105 == r_count_17_io_out ? io_r_261_b : _GEN_5450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5452 = 9'h106 == r_count_17_io_out ? io_r_262_b : _GEN_5451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5453 = 9'h107 == r_count_17_io_out ? io_r_263_b : _GEN_5452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5454 = 9'h108 == r_count_17_io_out ? io_r_264_b : _GEN_5453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5455 = 9'h109 == r_count_17_io_out ? io_r_265_b : _GEN_5454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5456 = 9'h10a == r_count_17_io_out ? io_r_266_b : _GEN_5455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5457 = 9'h10b == r_count_17_io_out ? io_r_267_b : _GEN_5456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5458 = 9'h10c == r_count_17_io_out ? io_r_268_b : _GEN_5457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5459 = 9'h10d == r_count_17_io_out ? io_r_269_b : _GEN_5458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5460 = 9'h10e == r_count_17_io_out ? io_r_270_b : _GEN_5459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5461 = 9'h10f == r_count_17_io_out ? io_r_271_b : _GEN_5460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5462 = 9'h110 == r_count_17_io_out ? io_r_272_b : _GEN_5461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5463 = 9'h111 == r_count_17_io_out ? io_r_273_b : _GEN_5462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5464 = 9'h112 == r_count_17_io_out ? io_r_274_b : _GEN_5463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5465 = 9'h113 == r_count_17_io_out ? io_r_275_b : _GEN_5464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5466 = 9'h114 == r_count_17_io_out ? io_r_276_b : _GEN_5465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5467 = 9'h115 == r_count_17_io_out ? io_r_277_b : _GEN_5466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5468 = 9'h116 == r_count_17_io_out ? io_r_278_b : _GEN_5467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5469 = 9'h117 == r_count_17_io_out ? io_r_279_b : _GEN_5468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5470 = 9'h118 == r_count_17_io_out ? io_r_280_b : _GEN_5469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5471 = 9'h119 == r_count_17_io_out ? io_r_281_b : _GEN_5470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5472 = 9'h11a == r_count_17_io_out ? io_r_282_b : _GEN_5471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5473 = 9'h11b == r_count_17_io_out ? io_r_283_b : _GEN_5472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5474 = 9'h11c == r_count_17_io_out ? io_r_284_b : _GEN_5473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5475 = 9'h11d == r_count_17_io_out ? io_r_285_b : _GEN_5474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5476 = 9'h11e == r_count_17_io_out ? io_r_286_b : _GEN_5475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5477 = 9'h11f == r_count_17_io_out ? io_r_287_b : _GEN_5476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5478 = 9'h120 == r_count_17_io_out ? io_r_288_b : _GEN_5477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5479 = 9'h121 == r_count_17_io_out ? io_r_289_b : _GEN_5478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5480 = 9'h122 == r_count_17_io_out ? io_r_290_b : _GEN_5479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5481 = 9'h123 == r_count_17_io_out ? io_r_291_b : _GEN_5480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5482 = 9'h124 == r_count_17_io_out ? io_r_292_b : _GEN_5481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5483 = 9'h125 == r_count_17_io_out ? io_r_293_b : _GEN_5482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5484 = 9'h126 == r_count_17_io_out ? io_r_294_b : _GEN_5483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5485 = 9'h127 == r_count_17_io_out ? io_r_295_b : _GEN_5484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5486 = 9'h128 == r_count_17_io_out ? io_r_296_b : _GEN_5485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5487 = 9'h129 == r_count_17_io_out ? io_r_297_b : _GEN_5486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5488 = 9'h12a == r_count_17_io_out ? io_r_298_b : _GEN_5487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5491 = 9'h1 == r_count_18_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5492 = 9'h2 == r_count_18_io_out ? io_r_2_b : _GEN_5491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5493 = 9'h3 == r_count_18_io_out ? io_r_3_b : _GEN_5492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5494 = 9'h4 == r_count_18_io_out ? io_r_4_b : _GEN_5493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5495 = 9'h5 == r_count_18_io_out ? io_r_5_b : _GEN_5494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5496 = 9'h6 == r_count_18_io_out ? io_r_6_b : _GEN_5495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5497 = 9'h7 == r_count_18_io_out ? io_r_7_b : _GEN_5496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5498 = 9'h8 == r_count_18_io_out ? io_r_8_b : _GEN_5497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5499 = 9'h9 == r_count_18_io_out ? io_r_9_b : _GEN_5498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5500 = 9'ha == r_count_18_io_out ? io_r_10_b : _GEN_5499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5501 = 9'hb == r_count_18_io_out ? io_r_11_b : _GEN_5500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5502 = 9'hc == r_count_18_io_out ? io_r_12_b : _GEN_5501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5503 = 9'hd == r_count_18_io_out ? io_r_13_b : _GEN_5502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5504 = 9'he == r_count_18_io_out ? io_r_14_b : _GEN_5503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5505 = 9'hf == r_count_18_io_out ? io_r_15_b : _GEN_5504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5506 = 9'h10 == r_count_18_io_out ? io_r_16_b : _GEN_5505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5507 = 9'h11 == r_count_18_io_out ? io_r_17_b : _GEN_5506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5508 = 9'h12 == r_count_18_io_out ? io_r_18_b : _GEN_5507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5509 = 9'h13 == r_count_18_io_out ? io_r_19_b : _GEN_5508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5510 = 9'h14 == r_count_18_io_out ? io_r_20_b : _GEN_5509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5511 = 9'h15 == r_count_18_io_out ? io_r_21_b : _GEN_5510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5512 = 9'h16 == r_count_18_io_out ? io_r_22_b : _GEN_5511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5513 = 9'h17 == r_count_18_io_out ? io_r_23_b : _GEN_5512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5514 = 9'h18 == r_count_18_io_out ? io_r_24_b : _GEN_5513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5515 = 9'h19 == r_count_18_io_out ? io_r_25_b : _GEN_5514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5516 = 9'h1a == r_count_18_io_out ? io_r_26_b : _GEN_5515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5517 = 9'h1b == r_count_18_io_out ? io_r_27_b : _GEN_5516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5518 = 9'h1c == r_count_18_io_out ? io_r_28_b : _GEN_5517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5519 = 9'h1d == r_count_18_io_out ? io_r_29_b : _GEN_5518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5520 = 9'h1e == r_count_18_io_out ? io_r_30_b : _GEN_5519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5521 = 9'h1f == r_count_18_io_out ? io_r_31_b : _GEN_5520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5522 = 9'h20 == r_count_18_io_out ? io_r_32_b : _GEN_5521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5523 = 9'h21 == r_count_18_io_out ? io_r_33_b : _GEN_5522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5524 = 9'h22 == r_count_18_io_out ? io_r_34_b : _GEN_5523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5525 = 9'h23 == r_count_18_io_out ? io_r_35_b : _GEN_5524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5526 = 9'h24 == r_count_18_io_out ? io_r_36_b : _GEN_5525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5527 = 9'h25 == r_count_18_io_out ? io_r_37_b : _GEN_5526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5528 = 9'h26 == r_count_18_io_out ? io_r_38_b : _GEN_5527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5529 = 9'h27 == r_count_18_io_out ? io_r_39_b : _GEN_5528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5530 = 9'h28 == r_count_18_io_out ? io_r_40_b : _GEN_5529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5531 = 9'h29 == r_count_18_io_out ? io_r_41_b : _GEN_5530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5532 = 9'h2a == r_count_18_io_out ? io_r_42_b : _GEN_5531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5533 = 9'h2b == r_count_18_io_out ? io_r_43_b : _GEN_5532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5534 = 9'h2c == r_count_18_io_out ? io_r_44_b : _GEN_5533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5535 = 9'h2d == r_count_18_io_out ? io_r_45_b : _GEN_5534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5536 = 9'h2e == r_count_18_io_out ? io_r_46_b : _GEN_5535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5537 = 9'h2f == r_count_18_io_out ? io_r_47_b : _GEN_5536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5538 = 9'h30 == r_count_18_io_out ? io_r_48_b : _GEN_5537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5539 = 9'h31 == r_count_18_io_out ? io_r_49_b : _GEN_5538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5540 = 9'h32 == r_count_18_io_out ? io_r_50_b : _GEN_5539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5541 = 9'h33 == r_count_18_io_out ? io_r_51_b : _GEN_5540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5542 = 9'h34 == r_count_18_io_out ? io_r_52_b : _GEN_5541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5543 = 9'h35 == r_count_18_io_out ? io_r_53_b : _GEN_5542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5544 = 9'h36 == r_count_18_io_out ? io_r_54_b : _GEN_5543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5545 = 9'h37 == r_count_18_io_out ? io_r_55_b : _GEN_5544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5546 = 9'h38 == r_count_18_io_out ? io_r_56_b : _GEN_5545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5547 = 9'h39 == r_count_18_io_out ? io_r_57_b : _GEN_5546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5548 = 9'h3a == r_count_18_io_out ? io_r_58_b : _GEN_5547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5549 = 9'h3b == r_count_18_io_out ? io_r_59_b : _GEN_5548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5550 = 9'h3c == r_count_18_io_out ? io_r_60_b : _GEN_5549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5551 = 9'h3d == r_count_18_io_out ? io_r_61_b : _GEN_5550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5552 = 9'h3e == r_count_18_io_out ? io_r_62_b : _GEN_5551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5553 = 9'h3f == r_count_18_io_out ? io_r_63_b : _GEN_5552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5554 = 9'h40 == r_count_18_io_out ? io_r_64_b : _GEN_5553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5555 = 9'h41 == r_count_18_io_out ? io_r_65_b : _GEN_5554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5556 = 9'h42 == r_count_18_io_out ? io_r_66_b : _GEN_5555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5557 = 9'h43 == r_count_18_io_out ? io_r_67_b : _GEN_5556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5558 = 9'h44 == r_count_18_io_out ? io_r_68_b : _GEN_5557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5559 = 9'h45 == r_count_18_io_out ? io_r_69_b : _GEN_5558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5560 = 9'h46 == r_count_18_io_out ? io_r_70_b : _GEN_5559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5561 = 9'h47 == r_count_18_io_out ? io_r_71_b : _GEN_5560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5562 = 9'h48 == r_count_18_io_out ? io_r_72_b : _GEN_5561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5563 = 9'h49 == r_count_18_io_out ? io_r_73_b : _GEN_5562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5564 = 9'h4a == r_count_18_io_out ? io_r_74_b : _GEN_5563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5565 = 9'h4b == r_count_18_io_out ? io_r_75_b : _GEN_5564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5566 = 9'h4c == r_count_18_io_out ? io_r_76_b : _GEN_5565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5567 = 9'h4d == r_count_18_io_out ? io_r_77_b : _GEN_5566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5568 = 9'h4e == r_count_18_io_out ? io_r_78_b : _GEN_5567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5569 = 9'h4f == r_count_18_io_out ? io_r_79_b : _GEN_5568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5570 = 9'h50 == r_count_18_io_out ? io_r_80_b : _GEN_5569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5571 = 9'h51 == r_count_18_io_out ? io_r_81_b : _GEN_5570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5572 = 9'h52 == r_count_18_io_out ? io_r_82_b : _GEN_5571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5573 = 9'h53 == r_count_18_io_out ? io_r_83_b : _GEN_5572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5574 = 9'h54 == r_count_18_io_out ? io_r_84_b : _GEN_5573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5575 = 9'h55 == r_count_18_io_out ? io_r_85_b : _GEN_5574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5576 = 9'h56 == r_count_18_io_out ? io_r_86_b : _GEN_5575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5577 = 9'h57 == r_count_18_io_out ? io_r_87_b : _GEN_5576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5578 = 9'h58 == r_count_18_io_out ? io_r_88_b : _GEN_5577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5579 = 9'h59 == r_count_18_io_out ? io_r_89_b : _GEN_5578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5580 = 9'h5a == r_count_18_io_out ? io_r_90_b : _GEN_5579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5581 = 9'h5b == r_count_18_io_out ? io_r_91_b : _GEN_5580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5582 = 9'h5c == r_count_18_io_out ? io_r_92_b : _GEN_5581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5583 = 9'h5d == r_count_18_io_out ? io_r_93_b : _GEN_5582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5584 = 9'h5e == r_count_18_io_out ? io_r_94_b : _GEN_5583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5585 = 9'h5f == r_count_18_io_out ? io_r_95_b : _GEN_5584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5586 = 9'h60 == r_count_18_io_out ? io_r_96_b : _GEN_5585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5587 = 9'h61 == r_count_18_io_out ? io_r_97_b : _GEN_5586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5588 = 9'h62 == r_count_18_io_out ? io_r_98_b : _GEN_5587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5589 = 9'h63 == r_count_18_io_out ? io_r_99_b : _GEN_5588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5590 = 9'h64 == r_count_18_io_out ? io_r_100_b : _GEN_5589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5591 = 9'h65 == r_count_18_io_out ? io_r_101_b : _GEN_5590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5592 = 9'h66 == r_count_18_io_out ? io_r_102_b : _GEN_5591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5593 = 9'h67 == r_count_18_io_out ? io_r_103_b : _GEN_5592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5594 = 9'h68 == r_count_18_io_out ? io_r_104_b : _GEN_5593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5595 = 9'h69 == r_count_18_io_out ? io_r_105_b : _GEN_5594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5596 = 9'h6a == r_count_18_io_out ? io_r_106_b : _GEN_5595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5597 = 9'h6b == r_count_18_io_out ? io_r_107_b : _GEN_5596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5598 = 9'h6c == r_count_18_io_out ? io_r_108_b : _GEN_5597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5599 = 9'h6d == r_count_18_io_out ? io_r_109_b : _GEN_5598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5600 = 9'h6e == r_count_18_io_out ? io_r_110_b : _GEN_5599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5601 = 9'h6f == r_count_18_io_out ? io_r_111_b : _GEN_5600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5602 = 9'h70 == r_count_18_io_out ? io_r_112_b : _GEN_5601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5603 = 9'h71 == r_count_18_io_out ? io_r_113_b : _GEN_5602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5604 = 9'h72 == r_count_18_io_out ? io_r_114_b : _GEN_5603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5605 = 9'h73 == r_count_18_io_out ? io_r_115_b : _GEN_5604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5606 = 9'h74 == r_count_18_io_out ? io_r_116_b : _GEN_5605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5607 = 9'h75 == r_count_18_io_out ? io_r_117_b : _GEN_5606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5608 = 9'h76 == r_count_18_io_out ? io_r_118_b : _GEN_5607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5609 = 9'h77 == r_count_18_io_out ? io_r_119_b : _GEN_5608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5610 = 9'h78 == r_count_18_io_out ? io_r_120_b : _GEN_5609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5611 = 9'h79 == r_count_18_io_out ? io_r_121_b : _GEN_5610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5612 = 9'h7a == r_count_18_io_out ? io_r_122_b : _GEN_5611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5613 = 9'h7b == r_count_18_io_out ? io_r_123_b : _GEN_5612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5614 = 9'h7c == r_count_18_io_out ? io_r_124_b : _GEN_5613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5615 = 9'h7d == r_count_18_io_out ? io_r_125_b : _GEN_5614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5616 = 9'h7e == r_count_18_io_out ? io_r_126_b : _GEN_5615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5617 = 9'h7f == r_count_18_io_out ? io_r_127_b : _GEN_5616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5618 = 9'h80 == r_count_18_io_out ? io_r_128_b : _GEN_5617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5619 = 9'h81 == r_count_18_io_out ? io_r_129_b : _GEN_5618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5620 = 9'h82 == r_count_18_io_out ? io_r_130_b : _GEN_5619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5621 = 9'h83 == r_count_18_io_out ? io_r_131_b : _GEN_5620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5622 = 9'h84 == r_count_18_io_out ? io_r_132_b : _GEN_5621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5623 = 9'h85 == r_count_18_io_out ? io_r_133_b : _GEN_5622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5624 = 9'h86 == r_count_18_io_out ? io_r_134_b : _GEN_5623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5625 = 9'h87 == r_count_18_io_out ? io_r_135_b : _GEN_5624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5626 = 9'h88 == r_count_18_io_out ? io_r_136_b : _GEN_5625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5627 = 9'h89 == r_count_18_io_out ? io_r_137_b : _GEN_5626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5628 = 9'h8a == r_count_18_io_out ? io_r_138_b : _GEN_5627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5629 = 9'h8b == r_count_18_io_out ? io_r_139_b : _GEN_5628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5630 = 9'h8c == r_count_18_io_out ? io_r_140_b : _GEN_5629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5631 = 9'h8d == r_count_18_io_out ? io_r_141_b : _GEN_5630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5632 = 9'h8e == r_count_18_io_out ? io_r_142_b : _GEN_5631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5633 = 9'h8f == r_count_18_io_out ? io_r_143_b : _GEN_5632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5634 = 9'h90 == r_count_18_io_out ? io_r_144_b : _GEN_5633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5635 = 9'h91 == r_count_18_io_out ? io_r_145_b : _GEN_5634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5636 = 9'h92 == r_count_18_io_out ? io_r_146_b : _GEN_5635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5637 = 9'h93 == r_count_18_io_out ? io_r_147_b : _GEN_5636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5638 = 9'h94 == r_count_18_io_out ? io_r_148_b : _GEN_5637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5639 = 9'h95 == r_count_18_io_out ? io_r_149_b : _GEN_5638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5640 = 9'h96 == r_count_18_io_out ? io_r_150_b : _GEN_5639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5641 = 9'h97 == r_count_18_io_out ? io_r_151_b : _GEN_5640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5642 = 9'h98 == r_count_18_io_out ? io_r_152_b : _GEN_5641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5643 = 9'h99 == r_count_18_io_out ? io_r_153_b : _GEN_5642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5644 = 9'h9a == r_count_18_io_out ? io_r_154_b : _GEN_5643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5645 = 9'h9b == r_count_18_io_out ? io_r_155_b : _GEN_5644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5646 = 9'h9c == r_count_18_io_out ? io_r_156_b : _GEN_5645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5647 = 9'h9d == r_count_18_io_out ? io_r_157_b : _GEN_5646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5648 = 9'h9e == r_count_18_io_out ? io_r_158_b : _GEN_5647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5649 = 9'h9f == r_count_18_io_out ? io_r_159_b : _GEN_5648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5650 = 9'ha0 == r_count_18_io_out ? io_r_160_b : _GEN_5649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5651 = 9'ha1 == r_count_18_io_out ? io_r_161_b : _GEN_5650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5652 = 9'ha2 == r_count_18_io_out ? io_r_162_b : _GEN_5651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5653 = 9'ha3 == r_count_18_io_out ? io_r_163_b : _GEN_5652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5654 = 9'ha4 == r_count_18_io_out ? io_r_164_b : _GEN_5653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5655 = 9'ha5 == r_count_18_io_out ? io_r_165_b : _GEN_5654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5656 = 9'ha6 == r_count_18_io_out ? io_r_166_b : _GEN_5655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5657 = 9'ha7 == r_count_18_io_out ? io_r_167_b : _GEN_5656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5658 = 9'ha8 == r_count_18_io_out ? io_r_168_b : _GEN_5657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5659 = 9'ha9 == r_count_18_io_out ? io_r_169_b : _GEN_5658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5660 = 9'haa == r_count_18_io_out ? io_r_170_b : _GEN_5659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5661 = 9'hab == r_count_18_io_out ? io_r_171_b : _GEN_5660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5662 = 9'hac == r_count_18_io_out ? io_r_172_b : _GEN_5661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5663 = 9'had == r_count_18_io_out ? io_r_173_b : _GEN_5662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5664 = 9'hae == r_count_18_io_out ? io_r_174_b : _GEN_5663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5665 = 9'haf == r_count_18_io_out ? io_r_175_b : _GEN_5664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5666 = 9'hb0 == r_count_18_io_out ? io_r_176_b : _GEN_5665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5667 = 9'hb1 == r_count_18_io_out ? io_r_177_b : _GEN_5666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5668 = 9'hb2 == r_count_18_io_out ? io_r_178_b : _GEN_5667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5669 = 9'hb3 == r_count_18_io_out ? io_r_179_b : _GEN_5668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5670 = 9'hb4 == r_count_18_io_out ? io_r_180_b : _GEN_5669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5671 = 9'hb5 == r_count_18_io_out ? io_r_181_b : _GEN_5670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5672 = 9'hb6 == r_count_18_io_out ? io_r_182_b : _GEN_5671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5673 = 9'hb7 == r_count_18_io_out ? io_r_183_b : _GEN_5672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5674 = 9'hb8 == r_count_18_io_out ? io_r_184_b : _GEN_5673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5675 = 9'hb9 == r_count_18_io_out ? io_r_185_b : _GEN_5674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5676 = 9'hba == r_count_18_io_out ? io_r_186_b : _GEN_5675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5677 = 9'hbb == r_count_18_io_out ? io_r_187_b : _GEN_5676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5678 = 9'hbc == r_count_18_io_out ? io_r_188_b : _GEN_5677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5679 = 9'hbd == r_count_18_io_out ? io_r_189_b : _GEN_5678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5680 = 9'hbe == r_count_18_io_out ? io_r_190_b : _GEN_5679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5681 = 9'hbf == r_count_18_io_out ? io_r_191_b : _GEN_5680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5682 = 9'hc0 == r_count_18_io_out ? io_r_192_b : _GEN_5681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5683 = 9'hc1 == r_count_18_io_out ? io_r_193_b : _GEN_5682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5684 = 9'hc2 == r_count_18_io_out ? io_r_194_b : _GEN_5683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5685 = 9'hc3 == r_count_18_io_out ? io_r_195_b : _GEN_5684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5686 = 9'hc4 == r_count_18_io_out ? io_r_196_b : _GEN_5685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5687 = 9'hc5 == r_count_18_io_out ? io_r_197_b : _GEN_5686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5688 = 9'hc6 == r_count_18_io_out ? io_r_198_b : _GEN_5687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5689 = 9'hc7 == r_count_18_io_out ? io_r_199_b : _GEN_5688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5690 = 9'hc8 == r_count_18_io_out ? io_r_200_b : _GEN_5689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5691 = 9'hc9 == r_count_18_io_out ? io_r_201_b : _GEN_5690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5692 = 9'hca == r_count_18_io_out ? io_r_202_b : _GEN_5691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5693 = 9'hcb == r_count_18_io_out ? io_r_203_b : _GEN_5692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5694 = 9'hcc == r_count_18_io_out ? io_r_204_b : _GEN_5693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5695 = 9'hcd == r_count_18_io_out ? io_r_205_b : _GEN_5694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5696 = 9'hce == r_count_18_io_out ? io_r_206_b : _GEN_5695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5697 = 9'hcf == r_count_18_io_out ? io_r_207_b : _GEN_5696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5698 = 9'hd0 == r_count_18_io_out ? io_r_208_b : _GEN_5697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5699 = 9'hd1 == r_count_18_io_out ? io_r_209_b : _GEN_5698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5700 = 9'hd2 == r_count_18_io_out ? io_r_210_b : _GEN_5699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5701 = 9'hd3 == r_count_18_io_out ? io_r_211_b : _GEN_5700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5702 = 9'hd4 == r_count_18_io_out ? io_r_212_b : _GEN_5701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5703 = 9'hd5 == r_count_18_io_out ? io_r_213_b : _GEN_5702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5704 = 9'hd6 == r_count_18_io_out ? io_r_214_b : _GEN_5703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5705 = 9'hd7 == r_count_18_io_out ? io_r_215_b : _GEN_5704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5706 = 9'hd8 == r_count_18_io_out ? io_r_216_b : _GEN_5705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5707 = 9'hd9 == r_count_18_io_out ? io_r_217_b : _GEN_5706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5708 = 9'hda == r_count_18_io_out ? io_r_218_b : _GEN_5707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5709 = 9'hdb == r_count_18_io_out ? io_r_219_b : _GEN_5708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5710 = 9'hdc == r_count_18_io_out ? io_r_220_b : _GEN_5709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5711 = 9'hdd == r_count_18_io_out ? io_r_221_b : _GEN_5710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5712 = 9'hde == r_count_18_io_out ? io_r_222_b : _GEN_5711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5713 = 9'hdf == r_count_18_io_out ? io_r_223_b : _GEN_5712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5714 = 9'he0 == r_count_18_io_out ? io_r_224_b : _GEN_5713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5715 = 9'he1 == r_count_18_io_out ? io_r_225_b : _GEN_5714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5716 = 9'he2 == r_count_18_io_out ? io_r_226_b : _GEN_5715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5717 = 9'he3 == r_count_18_io_out ? io_r_227_b : _GEN_5716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5718 = 9'he4 == r_count_18_io_out ? io_r_228_b : _GEN_5717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5719 = 9'he5 == r_count_18_io_out ? io_r_229_b : _GEN_5718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5720 = 9'he6 == r_count_18_io_out ? io_r_230_b : _GEN_5719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5721 = 9'he7 == r_count_18_io_out ? io_r_231_b : _GEN_5720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5722 = 9'he8 == r_count_18_io_out ? io_r_232_b : _GEN_5721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5723 = 9'he9 == r_count_18_io_out ? io_r_233_b : _GEN_5722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5724 = 9'hea == r_count_18_io_out ? io_r_234_b : _GEN_5723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5725 = 9'heb == r_count_18_io_out ? io_r_235_b : _GEN_5724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5726 = 9'hec == r_count_18_io_out ? io_r_236_b : _GEN_5725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5727 = 9'hed == r_count_18_io_out ? io_r_237_b : _GEN_5726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5728 = 9'hee == r_count_18_io_out ? io_r_238_b : _GEN_5727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5729 = 9'hef == r_count_18_io_out ? io_r_239_b : _GEN_5728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5730 = 9'hf0 == r_count_18_io_out ? io_r_240_b : _GEN_5729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5731 = 9'hf1 == r_count_18_io_out ? io_r_241_b : _GEN_5730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5732 = 9'hf2 == r_count_18_io_out ? io_r_242_b : _GEN_5731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5733 = 9'hf3 == r_count_18_io_out ? io_r_243_b : _GEN_5732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5734 = 9'hf4 == r_count_18_io_out ? io_r_244_b : _GEN_5733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5735 = 9'hf5 == r_count_18_io_out ? io_r_245_b : _GEN_5734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5736 = 9'hf6 == r_count_18_io_out ? io_r_246_b : _GEN_5735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5737 = 9'hf7 == r_count_18_io_out ? io_r_247_b : _GEN_5736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5738 = 9'hf8 == r_count_18_io_out ? io_r_248_b : _GEN_5737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5739 = 9'hf9 == r_count_18_io_out ? io_r_249_b : _GEN_5738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5740 = 9'hfa == r_count_18_io_out ? io_r_250_b : _GEN_5739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5741 = 9'hfb == r_count_18_io_out ? io_r_251_b : _GEN_5740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5742 = 9'hfc == r_count_18_io_out ? io_r_252_b : _GEN_5741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5743 = 9'hfd == r_count_18_io_out ? io_r_253_b : _GEN_5742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5744 = 9'hfe == r_count_18_io_out ? io_r_254_b : _GEN_5743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5745 = 9'hff == r_count_18_io_out ? io_r_255_b : _GEN_5744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5746 = 9'h100 == r_count_18_io_out ? io_r_256_b : _GEN_5745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5747 = 9'h101 == r_count_18_io_out ? io_r_257_b : _GEN_5746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5748 = 9'h102 == r_count_18_io_out ? io_r_258_b : _GEN_5747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5749 = 9'h103 == r_count_18_io_out ? io_r_259_b : _GEN_5748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5750 = 9'h104 == r_count_18_io_out ? io_r_260_b : _GEN_5749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5751 = 9'h105 == r_count_18_io_out ? io_r_261_b : _GEN_5750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5752 = 9'h106 == r_count_18_io_out ? io_r_262_b : _GEN_5751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5753 = 9'h107 == r_count_18_io_out ? io_r_263_b : _GEN_5752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5754 = 9'h108 == r_count_18_io_out ? io_r_264_b : _GEN_5753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5755 = 9'h109 == r_count_18_io_out ? io_r_265_b : _GEN_5754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5756 = 9'h10a == r_count_18_io_out ? io_r_266_b : _GEN_5755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5757 = 9'h10b == r_count_18_io_out ? io_r_267_b : _GEN_5756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5758 = 9'h10c == r_count_18_io_out ? io_r_268_b : _GEN_5757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5759 = 9'h10d == r_count_18_io_out ? io_r_269_b : _GEN_5758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5760 = 9'h10e == r_count_18_io_out ? io_r_270_b : _GEN_5759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5761 = 9'h10f == r_count_18_io_out ? io_r_271_b : _GEN_5760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5762 = 9'h110 == r_count_18_io_out ? io_r_272_b : _GEN_5761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5763 = 9'h111 == r_count_18_io_out ? io_r_273_b : _GEN_5762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5764 = 9'h112 == r_count_18_io_out ? io_r_274_b : _GEN_5763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5765 = 9'h113 == r_count_18_io_out ? io_r_275_b : _GEN_5764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5766 = 9'h114 == r_count_18_io_out ? io_r_276_b : _GEN_5765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5767 = 9'h115 == r_count_18_io_out ? io_r_277_b : _GEN_5766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5768 = 9'h116 == r_count_18_io_out ? io_r_278_b : _GEN_5767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5769 = 9'h117 == r_count_18_io_out ? io_r_279_b : _GEN_5768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5770 = 9'h118 == r_count_18_io_out ? io_r_280_b : _GEN_5769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5771 = 9'h119 == r_count_18_io_out ? io_r_281_b : _GEN_5770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5772 = 9'h11a == r_count_18_io_out ? io_r_282_b : _GEN_5771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5773 = 9'h11b == r_count_18_io_out ? io_r_283_b : _GEN_5772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5774 = 9'h11c == r_count_18_io_out ? io_r_284_b : _GEN_5773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5775 = 9'h11d == r_count_18_io_out ? io_r_285_b : _GEN_5774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5776 = 9'h11e == r_count_18_io_out ? io_r_286_b : _GEN_5775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5777 = 9'h11f == r_count_18_io_out ? io_r_287_b : _GEN_5776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5778 = 9'h120 == r_count_18_io_out ? io_r_288_b : _GEN_5777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5779 = 9'h121 == r_count_18_io_out ? io_r_289_b : _GEN_5778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5780 = 9'h122 == r_count_18_io_out ? io_r_290_b : _GEN_5779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5781 = 9'h123 == r_count_18_io_out ? io_r_291_b : _GEN_5780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5782 = 9'h124 == r_count_18_io_out ? io_r_292_b : _GEN_5781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5783 = 9'h125 == r_count_18_io_out ? io_r_293_b : _GEN_5782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5784 = 9'h126 == r_count_18_io_out ? io_r_294_b : _GEN_5783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5785 = 9'h127 == r_count_18_io_out ? io_r_295_b : _GEN_5784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5786 = 9'h128 == r_count_18_io_out ? io_r_296_b : _GEN_5785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5787 = 9'h129 == r_count_18_io_out ? io_r_297_b : _GEN_5786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5788 = 9'h12a == r_count_18_io_out ? io_r_298_b : _GEN_5787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5791 = 9'h1 == r_count_19_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5792 = 9'h2 == r_count_19_io_out ? io_r_2_b : _GEN_5791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5793 = 9'h3 == r_count_19_io_out ? io_r_3_b : _GEN_5792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5794 = 9'h4 == r_count_19_io_out ? io_r_4_b : _GEN_5793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5795 = 9'h5 == r_count_19_io_out ? io_r_5_b : _GEN_5794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5796 = 9'h6 == r_count_19_io_out ? io_r_6_b : _GEN_5795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5797 = 9'h7 == r_count_19_io_out ? io_r_7_b : _GEN_5796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5798 = 9'h8 == r_count_19_io_out ? io_r_8_b : _GEN_5797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5799 = 9'h9 == r_count_19_io_out ? io_r_9_b : _GEN_5798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5800 = 9'ha == r_count_19_io_out ? io_r_10_b : _GEN_5799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5801 = 9'hb == r_count_19_io_out ? io_r_11_b : _GEN_5800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5802 = 9'hc == r_count_19_io_out ? io_r_12_b : _GEN_5801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5803 = 9'hd == r_count_19_io_out ? io_r_13_b : _GEN_5802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5804 = 9'he == r_count_19_io_out ? io_r_14_b : _GEN_5803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5805 = 9'hf == r_count_19_io_out ? io_r_15_b : _GEN_5804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5806 = 9'h10 == r_count_19_io_out ? io_r_16_b : _GEN_5805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5807 = 9'h11 == r_count_19_io_out ? io_r_17_b : _GEN_5806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5808 = 9'h12 == r_count_19_io_out ? io_r_18_b : _GEN_5807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5809 = 9'h13 == r_count_19_io_out ? io_r_19_b : _GEN_5808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5810 = 9'h14 == r_count_19_io_out ? io_r_20_b : _GEN_5809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5811 = 9'h15 == r_count_19_io_out ? io_r_21_b : _GEN_5810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5812 = 9'h16 == r_count_19_io_out ? io_r_22_b : _GEN_5811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5813 = 9'h17 == r_count_19_io_out ? io_r_23_b : _GEN_5812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5814 = 9'h18 == r_count_19_io_out ? io_r_24_b : _GEN_5813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5815 = 9'h19 == r_count_19_io_out ? io_r_25_b : _GEN_5814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5816 = 9'h1a == r_count_19_io_out ? io_r_26_b : _GEN_5815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5817 = 9'h1b == r_count_19_io_out ? io_r_27_b : _GEN_5816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5818 = 9'h1c == r_count_19_io_out ? io_r_28_b : _GEN_5817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5819 = 9'h1d == r_count_19_io_out ? io_r_29_b : _GEN_5818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5820 = 9'h1e == r_count_19_io_out ? io_r_30_b : _GEN_5819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5821 = 9'h1f == r_count_19_io_out ? io_r_31_b : _GEN_5820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5822 = 9'h20 == r_count_19_io_out ? io_r_32_b : _GEN_5821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5823 = 9'h21 == r_count_19_io_out ? io_r_33_b : _GEN_5822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5824 = 9'h22 == r_count_19_io_out ? io_r_34_b : _GEN_5823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5825 = 9'h23 == r_count_19_io_out ? io_r_35_b : _GEN_5824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5826 = 9'h24 == r_count_19_io_out ? io_r_36_b : _GEN_5825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5827 = 9'h25 == r_count_19_io_out ? io_r_37_b : _GEN_5826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5828 = 9'h26 == r_count_19_io_out ? io_r_38_b : _GEN_5827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5829 = 9'h27 == r_count_19_io_out ? io_r_39_b : _GEN_5828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5830 = 9'h28 == r_count_19_io_out ? io_r_40_b : _GEN_5829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5831 = 9'h29 == r_count_19_io_out ? io_r_41_b : _GEN_5830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5832 = 9'h2a == r_count_19_io_out ? io_r_42_b : _GEN_5831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5833 = 9'h2b == r_count_19_io_out ? io_r_43_b : _GEN_5832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5834 = 9'h2c == r_count_19_io_out ? io_r_44_b : _GEN_5833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5835 = 9'h2d == r_count_19_io_out ? io_r_45_b : _GEN_5834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5836 = 9'h2e == r_count_19_io_out ? io_r_46_b : _GEN_5835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5837 = 9'h2f == r_count_19_io_out ? io_r_47_b : _GEN_5836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5838 = 9'h30 == r_count_19_io_out ? io_r_48_b : _GEN_5837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5839 = 9'h31 == r_count_19_io_out ? io_r_49_b : _GEN_5838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5840 = 9'h32 == r_count_19_io_out ? io_r_50_b : _GEN_5839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5841 = 9'h33 == r_count_19_io_out ? io_r_51_b : _GEN_5840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5842 = 9'h34 == r_count_19_io_out ? io_r_52_b : _GEN_5841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5843 = 9'h35 == r_count_19_io_out ? io_r_53_b : _GEN_5842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5844 = 9'h36 == r_count_19_io_out ? io_r_54_b : _GEN_5843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5845 = 9'h37 == r_count_19_io_out ? io_r_55_b : _GEN_5844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5846 = 9'h38 == r_count_19_io_out ? io_r_56_b : _GEN_5845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5847 = 9'h39 == r_count_19_io_out ? io_r_57_b : _GEN_5846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5848 = 9'h3a == r_count_19_io_out ? io_r_58_b : _GEN_5847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5849 = 9'h3b == r_count_19_io_out ? io_r_59_b : _GEN_5848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5850 = 9'h3c == r_count_19_io_out ? io_r_60_b : _GEN_5849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5851 = 9'h3d == r_count_19_io_out ? io_r_61_b : _GEN_5850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5852 = 9'h3e == r_count_19_io_out ? io_r_62_b : _GEN_5851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5853 = 9'h3f == r_count_19_io_out ? io_r_63_b : _GEN_5852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5854 = 9'h40 == r_count_19_io_out ? io_r_64_b : _GEN_5853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5855 = 9'h41 == r_count_19_io_out ? io_r_65_b : _GEN_5854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5856 = 9'h42 == r_count_19_io_out ? io_r_66_b : _GEN_5855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5857 = 9'h43 == r_count_19_io_out ? io_r_67_b : _GEN_5856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5858 = 9'h44 == r_count_19_io_out ? io_r_68_b : _GEN_5857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5859 = 9'h45 == r_count_19_io_out ? io_r_69_b : _GEN_5858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5860 = 9'h46 == r_count_19_io_out ? io_r_70_b : _GEN_5859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5861 = 9'h47 == r_count_19_io_out ? io_r_71_b : _GEN_5860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5862 = 9'h48 == r_count_19_io_out ? io_r_72_b : _GEN_5861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5863 = 9'h49 == r_count_19_io_out ? io_r_73_b : _GEN_5862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5864 = 9'h4a == r_count_19_io_out ? io_r_74_b : _GEN_5863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5865 = 9'h4b == r_count_19_io_out ? io_r_75_b : _GEN_5864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5866 = 9'h4c == r_count_19_io_out ? io_r_76_b : _GEN_5865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5867 = 9'h4d == r_count_19_io_out ? io_r_77_b : _GEN_5866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5868 = 9'h4e == r_count_19_io_out ? io_r_78_b : _GEN_5867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5869 = 9'h4f == r_count_19_io_out ? io_r_79_b : _GEN_5868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5870 = 9'h50 == r_count_19_io_out ? io_r_80_b : _GEN_5869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5871 = 9'h51 == r_count_19_io_out ? io_r_81_b : _GEN_5870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5872 = 9'h52 == r_count_19_io_out ? io_r_82_b : _GEN_5871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5873 = 9'h53 == r_count_19_io_out ? io_r_83_b : _GEN_5872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5874 = 9'h54 == r_count_19_io_out ? io_r_84_b : _GEN_5873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5875 = 9'h55 == r_count_19_io_out ? io_r_85_b : _GEN_5874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5876 = 9'h56 == r_count_19_io_out ? io_r_86_b : _GEN_5875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5877 = 9'h57 == r_count_19_io_out ? io_r_87_b : _GEN_5876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5878 = 9'h58 == r_count_19_io_out ? io_r_88_b : _GEN_5877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5879 = 9'h59 == r_count_19_io_out ? io_r_89_b : _GEN_5878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5880 = 9'h5a == r_count_19_io_out ? io_r_90_b : _GEN_5879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5881 = 9'h5b == r_count_19_io_out ? io_r_91_b : _GEN_5880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5882 = 9'h5c == r_count_19_io_out ? io_r_92_b : _GEN_5881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5883 = 9'h5d == r_count_19_io_out ? io_r_93_b : _GEN_5882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5884 = 9'h5e == r_count_19_io_out ? io_r_94_b : _GEN_5883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5885 = 9'h5f == r_count_19_io_out ? io_r_95_b : _GEN_5884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5886 = 9'h60 == r_count_19_io_out ? io_r_96_b : _GEN_5885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5887 = 9'h61 == r_count_19_io_out ? io_r_97_b : _GEN_5886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5888 = 9'h62 == r_count_19_io_out ? io_r_98_b : _GEN_5887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5889 = 9'h63 == r_count_19_io_out ? io_r_99_b : _GEN_5888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5890 = 9'h64 == r_count_19_io_out ? io_r_100_b : _GEN_5889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5891 = 9'h65 == r_count_19_io_out ? io_r_101_b : _GEN_5890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5892 = 9'h66 == r_count_19_io_out ? io_r_102_b : _GEN_5891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5893 = 9'h67 == r_count_19_io_out ? io_r_103_b : _GEN_5892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5894 = 9'h68 == r_count_19_io_out ? io_r_104_b : _GEN_5893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5895 = 9'h69 == r_count_19_io_out ? io_r_105_b : _GEN_5894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5896 = 9'h6a == r_count_19_io_out ? io_r_106_b : _GEN_5895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5897 = 9'h6b == r_count_19_io_out ? io_r_107_b : _GEN_5896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5898 = 9'h6c == r_count_19_io_out ? io_r_108_b : _GEN_5897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5899 = 9'h6d == r_count_19_io_out ? io_r_109_b : _GEN_5898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5900 = 9'h6e == r_count_19_io_out ? io_r_110_b : _GEN_5899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5901 = 9'h6f == r_count_19_io_out ? io_r_111_b : _GEN_5900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5902 = 9'h70 == r_count_19_io_out ? io_r_112_b : _GEN_5901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5903 = 9'h71 == r_count_19_io_out ? io_r_113_b : _GEN_5902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5904 = 9'h72 == r_count_19_io_out ? io_r_114_b : _GEN_5903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5905 = 9'h73 == r_count_19_io_out ? io_r_115_b : _GEN_5904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5906 = 9'h74 == r_count_19_io_out ? io_r_116_b : _GEN_5905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5907 = 9'h75 == r_count_19_io_out ? io_r_117_b : _GEN_5906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5908 = 9'h76 == r_count_19_io_out ? io_r_118_b : _GEN_5907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5909 = 9'h77 == r_count_19_io_out ? io_r_119_b : _GEN_5908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5910 = 9'h78 == r_count_19_io_out ? io_r_120_b : _GEN_5909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5911 = 9'h79 == r_count_19_io_out ? io_r_121_b : _GEN_5910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5912 = 9'h7a == r_count_19_io_out ? io_r_122_b : _GEN_5911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5913 = 9'h7b == r_count_19_io_out ? io_r_123_b : _GEN_5912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5914 = 9'h7c == r_count_19_io_out ? io_r_124_b : _GEN_5913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5915 = 9'h7d == r_count_19_io_out ? io_r_125_b : _GEN_5914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5916 = 9'h7e == r_count_19_io_out ? io_r_126_b : _GEN_5915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5917 = 9'h7f == r_count_19_io_out ? io_r_127_b : _GEN_5916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5918 = 9'h80 == r_count_19_io_out ? io_r_128_b : _GEN_5917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5919 = 9'h81 == r_count_19_io_out ? io_r_129_b : _GEN_5918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5920 = 9'h82 == r_count_19_io_out ? io_r_130_b : _GEN_5919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5921 = 9'h83 == r_count_19_io_out ? io_r_131_b : _GEN_5920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5922 = 9'h84 == r_count_19_io_out ? io_r_132_b : _GEN_5921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5923 = 9'h85 == r_count_19_io_out ? io_r_133_b : _GEN_5922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5924 = 9'h86 == r_count_19_io_out ? io_r_134_b : _GEN_5923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5925 = 9'h87 == r_count_19_io_out ? io_r_135_b : _GEN_5924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5926 = 9'h88 == r_count_19_io_out ? io_r_136_b : _GEN_5925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5927 = 9'h89 == r_count_19_io_out ? io_r_137_b : _GEN_5926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5928 = 9'h8a == r_count_19_io_out ? io_r_138_b : _GEN_5927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5929 = 9'h8b == r_count_19_io_out ? io_r_139_b : _GEN_5928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5930 = 9'h8c == r_count_19_io_out ? io_r_140_b : _GEN_5929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5931 = 9'h8d == r_count_19_io_out ? io_r_141_b : _GEN_5930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5932 = 9'h8e == r_count_19_io_out ? io_r_142_b : _GEN_5931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5933 = 9'h8f == r_count_19_io_out ? io_r_143_b : _GEN_5932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5934 = 9'h90 == r_count_19_io_out ? io_r_144_b : _GEN_5933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5935 = 9'h91 == r_count_19_io_out ? io_r_145_b : _GEN_5934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5936 = 9'h92 == r_count_19_io_out ? io_r_146_b : _GEN_5935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5937 = 9'h93 == r_count_19_io_out ? io_r_147_b : _GEN_5936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5938 = 9'h94 == r_count_19_io_out ? io_r_148_b : _GEN_5937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5939 = 9'h95 == r_count_19_io_out ? io_r_149_b : _GEN_5938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5940 = 9'h96 == r_count_19_io_out ? io_r_150_b : _GEN_5939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5941 = 9'h97 == r_count_19_io_out ? io_r_151_b : _GEN_5940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5942 = 9'h98 == r_count_19_io_out ? io_r_152_b : _GEN_5941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5943 = 9'h99 == r_count_19_io_out ? io_r_153_b : _GEN_5942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5944 = 9'h9a == r_count_19_io_out ? io_r_154_b : _GEN_5943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5945 = 9'h9b == r_count_19_io_out ? io_r_155_b : _GEN_5944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5946 = 9'h9c == r_count_19_io_out ? io_r_156_b : _GEN_5945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5947 = 9'h9d == r_count_19_io_out ? io_r_157_b : _GEN_5946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5948 = 9'h9e == r_count_19_io_out ? io_r_158_b : _GEN_5947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5949 = 9'h9f == r_count_19_io_out ? io_r_159_b : _GEN_5948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5950 = 9'ha0 == r_count_19_io_out ? io_r_160_b : _GEN_5949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5951 = 9'ha1 == r_count_19_io_out ? io_r_161_b : _GEN_5950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5952 = 9'ha2 == r_count_19_io_out ? io_r_162_b : _GEN_5951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5953 = 9'ha3 == r_count_19_io_out ? io_r_163_b : _GEN_5952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5954 = 9'ha4 == r_count_19_io_out ? io_r_164_b : _GEN_5953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5955 = 9'ha5 == r_count_19_io_out ? io_r_165_b : _GEN_5954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5956 = 9'ha6 == r_count_19_io_out ? io_r_166_b : _GEN_5955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5957 = 9'ha7 == r_count_19_io_out ? io_r_167_b : _GEN_5956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5958 = 9'ha8 == r_count_19_io_out ? io_r_168_b : _GEN_5957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5959 = 9'ha9 == r_count_19_io_out ? io_r_169_b : _GEN_5958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5960 = 9'haa == r_count_19_io_out ? io_r_170_b : _GEN_5959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5961 = 9'hab == r_count_19_io_out ? io_r_171_b : _GEN_5960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5962 = 9'hac == r_count_19_io_out ? io_r_172_b : _GEN_5961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5963 = 9'had == r_count_19_io_out ? io_r_173_b : _GEN_5962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5964 = 9'hae == r_count_19_io_out ? io_r_174_b : _GEN_5963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5965 = 9'haf == r_count_19_io_out ? io_r_175_b : _GEN_5964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5966 = 9'hb0 == r_count_19_io_out ? io_r_176_b : _GEN_5965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5967 = 9'hb1 == r_count_19_io_out ? io_r_177_b : _GEN_5966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5968 = 9'hb2 == r_count_19_io_out ? io_r_178_b : _GEN_5967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5969 = 9'hb3 == r_count_19_io_out ? io_r_179_b : _GEN_5968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5970 = 9'hb4 == r_count_19_io_out ? io_r_180_b : _GEN_5969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5971 = 9'hb5 == r_count_19_io_out ? io_r_181_b : _GEN_5970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5972 = 9'hb6 == r_count_19_io_out ? io_r_182_b : _GEN_5971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5973 = 9'hb7 == r_count_19_io_out ? io_r_183_b : _GEN_5972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5974 = 9'hb8 == r_count_19_io_out ? io_r_184_b : _GEN_5973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5975 = 9'hb9 == r_count_19_io_out ? io_r_185_b : _GEN_5974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5976 = 9'hba == r_count_19_io_out ? io_r_186_b : _GEN_5975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5977 = 9'hbb == r_count_19_io_out ? io_r_187_b : _GEN_5976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5978 = 9'hbc == r_count_19_io_out ? io_r_188_b : _GEN_5977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5979 = 9'hbd == r_count_19_io_out ? io_r_189_b : _GEN_5978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5980 = 9'hbe == r_count_19_io_out ? io_r_190_b : _GEN_5979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5981 = 9'hbf == r_count_19_io_out ? io_r_191_b : _GEN_5980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5982 = 9'hc0 == r_count_19_io_out ? io_r_192_b : _GEN_5981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5983 = 9'hc1 == r_count_19_io_out ? io_r_193_b : _GEN_5982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5984 = 9'hc2 == r_count_19_io_out ? io_r_194_b : _GEN_5983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5985 = 9'hc3 == r_count_19_io_out ? io_r_195_b : _GEN_5984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5986 = 9'hc4 == r_count_19_io_out ? io_r_196_b : _GEN_5985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5987 = 9'hc5 == r_count_19_io_out ? io_r_197_b : _GEN_5986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5988 = 9'hc6 == r_count_19_io_out ? io_r_198_b : _GEN_5987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5989 = 9'hc7 == r_count_19_io_out ? io_r_199_b : _GEN_5988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5990 = 9'hc8 == r_count_19_io_out ? io_r_200_b : _GEN_5989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5991 = 9'hc9 == r_count_19_io_out ? io_r_201_b : _GEN_5990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5992 = 9'hca == r_count_19_io_out ? io_r_202_b : _GEN_5991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5993 = 9'hcb == r_count_19_io_out ? io_r_203_b : _GEN_5992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5994 = 9'hcc == r_count_19_io_out ? io_r_204_b : _GEN_5993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5995 = 9'hcd == r_count_19_io_out ? io_r_205_b : _GEN_5994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5996 = 9'hce == r_count_19_io_out ? io_r_206_b : _GEN_5995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5997 = 9'hcf == r_count_19_io_out ? io_r_207_b : _GEN_5996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5998 = 9'hd0 == r_count_19_io_out ? io_r_208_b : _GEN_5997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5999 = 9'hd1 == r_count_19_io_out ? io_r_209_b : _GEN_5998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6000 = 9'hd2 == r_count_19_io_out ? io_r_210_b : _GEN_5999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6001 = 9'hd3 == r_count_19_io_out ? io_r_211_b : _GEN_6000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6002 = 9'hd4 == r_count_19_io_out ? io_r_212_b : _GEN_6001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6003 = 9'hd5 == r_count_19_io_out ? io_r_213_b : _GEN_6002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6004 = 9'hd6 == r_count_19_io_out ? io_r_214_b : _GEN_6003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6005 = 9'hd7 == r_count_19_io_out ? io_r_215_b : _GEN_6004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6006 = 9'hd8 == r_count_19_io_out ? io_r_216_b : _GEN_6005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6007 = 9'hd9 == r_count_19_io_out ? io_r_217_b : _GEN_6006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6008 = 9'hda == r_count_19_io_out ? io_r_218_b : _GEN_6007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6009 = 9'hdb == r_count_19_io_out ? io_r_219_b : _GEN_6008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6010 = 9'hdc == r_count_19_io_out ? io_r_220_b : _GEN_6009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6011 = 9'hdd == r_count_19_io_out ? io_r_221_b : _GEN_6010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6012 = 9'hde == r_count_19_io_out ? io_r_222_b : _GEN_6011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6013 = 9'hdf == r_count_19_io_out ? io_r_223_b : _GEN_6012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6014 = 9'he0 == r_count_19_io_out ? io_r_224_b : _GEN_6013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6015 = 9'he1 == r_count_19_io_out ? io_r_225_b : _GEN_6014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6016 = 9'he2 == r_count_19_io_out ? io_r_226_b : _GEN_6015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6017 = 9'he3 == r_count_19_io_out ? io_r_227_b : _GEN_6016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6018 = 9'he4 == r_count_19_io_out ? io_r_228_b : _GEN_6017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6019 = 9'he5 == r_count_19_io_out ? io_r_229_b : _GEN_6018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6020 = 9'he6 == r_count_19_io_out ? io_r_230_b : _GEN_6019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6021 = 9'he7 == r_count_19_io_out ? io_r_231_b : _GEN_6020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6022 = 9'he8 == r_count_19_io_out ? io_r_232_b : _GEN_6021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6023 = 9'he9 == r_count_19_io_out ? io_r_233_b : _GEN_6022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6024 = 9'hea == r_count_19_io_out ? io_r_234_b : _GEN_6023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6025 = 9'heb == r_count_19_io_out ? io_r_235_b : _GEN_6024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6026 = 9'hec == r_count_19_io_out ? io_r_236_b : _GEN_6025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6027 = 9'hed == r_count_19_io_out ? io_r_237_b : _GEN_6026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6028 = 9'hee == r_count_19_io_out ? io_r_238_b : _GEN_6027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6029 = 9'hef == r_count_19_io_out ? io_r_239_b : _GEN_6028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6030 = 9'hf0 == r_count_19_io_out ? io_r_240_b : _GEN_6029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6031 = 9'hf1 == r_count_19_io_out ? io_r_241_b : _GEN_6030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6032 = 9'hf2 == r_count_19_io_out ? io_r_242_b : _GEN_6031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6033 = 9'hf3 == r_count_19_io_out ? io_r_243_b : _GEN_6032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6034 = 9'hf4 == r_count_19_io_out ? io_r_244_b : _GEN_6033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6035 = 9'hf5 == r_count_19_io_out ? io_r_245_b : _GEN_6034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6036 = 9'hf6 == r_count_19_io_out ? io_r_246_b : _GEN_6035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6037 = 9'hf7 == r_count_19_io_out ? io_r_247_b : _GEN_6036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6038 = 9'hf8 == r_count_19_io_out ? io_r_248_b : _GEN_6037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6039 = 9'hf9 == r_count_19_io_out ? io_r_249_b : _GEN_6038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6040 = 9'hfa == r_count_19_io_out ? io_r_250_b : _GEN_6039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6041 = 9'hfb == r_count_19_io_out ? io_r_251_b : _GEN_6040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6042 = 9'hfc == r_count_19_io_out ? io_r_252_b : _GEN_6041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6043 = 9'hfd == r_count_19_io_out ? io_r_253_b : _GEN_6042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6044 = 9'hfe == r_count_19_io_out ? io_r_254_b : _GEN_6043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6045 = 9'hff == r_count_19_io_out ? io_r_255_b : _GEN_6044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6046 = 9'h100 == r_count_19_io_out ? io_r_256_b : _GEN_6045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6047 = 9'h101 == r_count_19_io_out ? io_r_257_b : _GEN_6046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6048 = 9'h102 == r_count_19_io_out ? io_r_258_b : _GEN_6047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6049 = 9'h103 == r_count_19_io_out ? io_r_259_b : _GEN_6048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6050 = 9'h104 == r_count_19_io_out ? io_r_260_b : _GEN_6049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6051 = 9'h105 == r_count_19_io_out ? io_r_261_b : _GEN_6050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6052 = 9'h106 == r_count_19_io_out ? io_r_262_b : _GEN_6051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6053 = 9'h107 == r_count_19_io_out ? io_r_263_b : _GEN_6052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6054 = 9'h108 == r_count_19_io_out ? io_r_264_b : _GEN_6053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6055 = 9'h109 == r_count_19_io_out ? io_r_265_b : _GEN_6054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6056 = 9'h10a == r_count_19_io_out ? io_r_266_b : _GEN_6055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6057 = 9'h10b == r_count_19_io_out ? io_r_267_b : _GEN_6056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6058 = 9'h10c == r_count_19_io_out ? io_r_268_b : _GEN_6057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6059 = 9'h10d == r_count_19_io_out ? io_r_269_b : _GEN_6058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6060 = 9'h10e == r_count_19_io_out ? io_r_270_b : _GEN_6059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6061 = 9'h10f == r_count_19_io_out ? io_r_271_b : _GEN_6060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6062 = 9'h110 == r_count_19_io_out ? io_r_272_b : _GEN_6061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6063 = 9'h111 == r_count_19_io_out ? io_r_273_b : _GEN_6062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6064 = 9'h112 == r_count_19_io_out ? io_r_274_b : _GEN_6063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6065 = 9'h113 == r_count_19_io_out ? io_r_275_b : _GEN_6064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6066 = 9'h114 == r_count_19_io_out ? io_r_276_b : _GEN_6065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6067 = 9'h115 == r_count_19_io_out ? io_r_277_b : _GEN_6066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6068 = 9'h116 == r_count_19_io_out ? io_r_278_b : _GEN_6067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6069 = 9'h117 == r_count_19_io_out ? io_r_279_b : _GEN_6068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6070 = 9'h118 == r_count_19_io_out ? io_r_280_b : _GEN_6069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6071 = 9'h119 == r_count_19_io_out ? io_r_281_b : _GEN_6070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6072 = 9'h11a == r_count_19_io_out ? io_r_282_b : _GEN_6071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6073 = 9'h11b == r_count_19_io_out ? io_r_283_b : _GEN_6072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6074 = 9'h11c == r_count_19_io_out ? io_r_284_b : _GEN_6073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6075 = 9'h11d == r_count_19_io_out ? io_r_285_b : _GEN_6074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6076 = 9'h11e == r_count_19_io_out ? io_r_286_b : _GEN_6075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6077 = 9'h11f == r_count_19_io_out ? io_r_287_b : _GEN_6076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6078 = 9'h120 == r_count_19_io_out ? io_r_288_b : _GEN_6077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6079 = 9'h121 == r_count_19_io_out ? io_r_289_b : _GEN_6078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6080 = 9'h122 == r_count_19_io_out ? io_r_290_b : _GEN_6079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6081 = 9'h123 == r_count_19_io_out ? io_r_291_b : _GEN_6080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6082 = 9'h124 == r_count_19_io_out ? io_r_292_b : _GEN_6081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6083 = 9'h125 == r_count_19_io_out ? io_r_293_b : _GEN_6082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6084 = 9'h126 == r_count_19_io_out ? io_r_294_b : _GEN_6083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6085 = 9'h127 == r_count_19_io_out ? io_r_295_b : _GEN_6084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6086 = 9'h128 == r_count_19_io_out ? io_r_296_b : _GEN_6085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6087 = 9'h129 == r_count_19_io_out ? io_r_297_b : _GEN_6086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6088 = 9'h12a == r_count_19_io_out ? io_r_298_b : _GEN_6087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6091 = 9'h1 == r_count_20_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6092 = 9'h2 == r_count_20_io_out ? io_r_2_b : _GEN_6091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6093 = 9'h3 == r_count_20_io_out ? io_r_3_b : _GEN_6092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6094 = 9'h4 == r_count_20_io_out ? io_r_4_b : _GEN_6093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6095 = 9'h5 == r_count_20_io_out ? io_r_5_b : _GEN_6094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6096 = 9'h6 == r_count_20_io_out ? io_r_6_b : _GEN_6095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6097 = 9'h7 == r_count_20_io_out ? io_r_7_b : _GEN_6096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6098 = 9'h8 == r_count_20_io_out ? io_r_8_b : _GEN_6097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6099 = 9'h9 == r_count_20_io_out ? io_r_9_b : _GEN_6098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6100 = 9'ha == r_count_20_io_out ? io_r_10_b : _GEN_6099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6101 = 9'hb == r_count_20_io_out ? io_r_11_b : _GEN_6100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6102 = 9'hc == r_count_20_io_out ? io_r_12_b : _GEN_6101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6103 = 9'hd == r_count_20_io_out ? io_r_13_b : _GEN_6102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6104 = 9'he == r_count_20_io_out ? io_r_14_b : _GEN_6103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6105 = 9'hf == r_count_20_io_out ? io_r_15_b : _GEN_6104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6106 = 9'h10 == r_count_20_io_out ? io_r_16_b : _GEN_6105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6107 = 9'h11 == r_count_20_io_out ? io_r_17_b : _GEN_6106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6108 = 9'h12 == r_count_20_io_out ? io_r_18_b : _GEN_6107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6109 = 9'h13 == r_count_20_io_out ? io_r_19_b : _GEN_6108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6110 = 9'h14 == r_count_20_io_out ? io_r_20_b : _GEN_6109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6111 = 9'h15 == r_count_20_io_out ? io_r_21_b : _GEN_6110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6112 = 9'h16 == r_count_20_io_out ? io_r_22_b : _GEN_6111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6113 = 9'h17 == r_count_20_io_out ? io_r_23_b : _GEN_6112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6114 = 9'h18 == r_count_20_io_out ? io_r_24_b : _GEN_6113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6115 = 9'h19 == r_count_20_io_out ? io_r_25_b : _GEN_6114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6116 = 9'h1a == r_count_20_io_out ? io_r_26_b : _GEN_6115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6117 = 9'h1b == r_count_20_io_out ? io_r_27_b : _GEN_6116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6118 = 9'h1c == r_count_20_io_out ? io_r_28_b : _GEN_6117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6119 = 9'h1d == r_count_20_io_out ? io_r_29_b : _GEN_6118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6120 = 9'h1e == r_count_20_io_out ? io_r_30_b : _GEN_6119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6121 = 9'h1f == r_count_20_io_out ? io_r_31_b : _GEN_6120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6122 = 9'h20 == r_count_20_io_out ? io_r_32_b : _GEN_6121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6123 = 9'h21 == r_count_20_io_out ? io_r_33_b : _GEN_6122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6124 = 9'h22 == r_count_20_io_out ? io_r_34_b : _GEN_6123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6125 = 9'h23 == r_count_20_io_out ? io_r_35_b : _GEN_6124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6126 = 9'h24 == r_count_20_io_out ? io_r_36_b : _GEN_6125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6127 = 9'h25 == r_count_20_io_out ? io_r_37_b : _GEN_6126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6128 = 9'h26 == r_count_20_io_out ? io_r_38_b : _GEN_6127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6129 = 9'h27 == r_count_20_io_out ? io_r_39_b : _GEN_6128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6130 = 9'h28 == r_count_20_io_out ? io_r_40_b : _GEN_6129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6131 = 9'h29 == r_count_20_io_out ? io_r_41_b : _GEN_6130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6132 = 9'h2a == r_count_20_io_out ? io_r_42_b : _GEN_6131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6133 = 9'h2b == r_count_20_io_out ? io_r_43_b : _GEN_6132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6134 = 9'h2c == r_count_20_io_out ? io_r_44_b : _GEN_6133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6135 = 9'h2d == r_count_20_io_out ? io_r_45_b : _GEN_6134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6136 = 9'h2e == r_count_20_io_out ? io_r_46_b : _GEN_6135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6137 = 9'h2f == r_count_20_io_out ? io_r_47_b : _GEN_6136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6138 = 9'h30 == r_count_20_io_out ? io_r_48_b : _GEN_6137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6139 = 9'h31 == r_count_20_io_out ? io_r_49_b : _GEN_6138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6140 = 9'h32 == r_count_20_io_out ? io_r_50_b : _GEN_6139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6141 = 9'h33 == r_count_20_io_out ? io_r_51_b : _GEN_6140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6142 = 9'h34 == r_count_20_io_out ? io_r_52_b : _GEN_6141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6143 = 9'h35 == r_count_20_io_out ? io_r_53_b : _GEN_6142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6144 = 9'h36 == r_count_20_io_out ? io_r_54_b : _GEN_6143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6145 = 9'h37 == r_count_20_io_out ? io_r_55_b : _GEN_6144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6146 = 9'h38 == r_count_20_io_out ? io_r_56_b : _GEN_6145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6147 = 9'h39 == r_count_20_io_out ? io_r_57_b : _GEN_6146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6148 = 9'h3a == r_count_20_io_out ? io_r_58_b : _GEN_6147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6149 = 9'h3b == r_count_20_io_out ? io_r_59_b : _GEN_6148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6150 = 9'h3c == r_count_20_io_out ? io_r_60_b : _GEN_6149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6151 = 9'h3d == r_count_20_io_out ? io_r_61_b : _GEN_6150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6152 = 9'h3e == r_count_20_io_out ? io_r_62_b : _GEN_6151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6153 = 9'h3f == r_count_20_io_out ? io_r_63_b : _GEN_6152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6154 = 9'h40 == r_count_20_io_out ? io_r_64_b : _GEN_6153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6155 = 9'h41 == r_count_20_io_out ? io_r_65_b : _GEN_6154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6156 = 9'h42 == r_count_20_io_out ? io_r_66_b : _GEN_6155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6157 = 9'h43 == r_count_20_io_out ? io_r_67_b : _GEN_6156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6158 = 9'h44 == r_count_20_io_out ? io_r_68_b : _GEN_6157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6159 = 9'h45 == r_count_20_io_out ? io_r_69_b : _GEN_6158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6160 = 9'h46 == r_count_20_io_out ? io_r_70_b : _GEN_6159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6161 = 9'h47 == r_count_20_io_out ? io_r_71_b : _GEN_6160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6162 = 9'h48 == r_count_20_io_out ? io_r_72_b : _GEN_6161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6163 = 9'h49 == r_count_20_io_out ? io_r_73_b : _GEN_6162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6164 = 9'h4a == r_count_20_io_out ? io_r_74_b : _GEN_6163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6165 = 9'h4b == r_count_20_io_out ? io_r_75_b : _GEN_6164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6166 = 9'h4c == r_count_20_io_out ? io_r_76_b : _GEN_6165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6167 = 9'h4d == r_count_20_io_out ? io_r_77_b : _GEN_6166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6168 = 9'h4e == r_count_20_io_out ? io_r_78_b : _GEN_6167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6169 = 9'h4f == r_count_20_io_out ? io_r_79_b : _GEN_6168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6170 = 9'h50 == r_count_20_io_out ? io_r_80_b : _GEN_6169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6171 = 9'h51 == r_count_20_io_out ? io_r_81_b : _GEN_6170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6172 = 9'h52 == r_count_20_io_out ? io_r_82_b : _GEN_6171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6173 = 9'h53 == r_count_20_io_out ? io_r_83_b : _GEN_6172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6174 = 9'h54 == r_count_20_io_out ? io_r_84_b : _GEN_6173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6175 = 9'h55 == r_count_20_io_out ? io_r_85_b : _GEN_6174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6176 = 9'h56 == r_count_20_io_out ? io_r_86_b : _GEN_6175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6177 = 9'h57 == r_count_20_io_out ? io_r_87_b : _GEN_6176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6178 = 9'h58 == r_count_20_io_out ? io_r_88_b : _GEN_6177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6179 = 9'h59 == r_count_20_io_out ? io_r_89_b : _GEN_6178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6180 = 9'h5a == r_count_20_io_out ? io_r_90_b : _GEN_6179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6181 = 9'h5b == r_count_20_io_out ? io_r_91_b : _GEN_6180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6182 = 9'h5c == r_count_20_io_out ? io_r_92_b : _GEN_6181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6183 = 9'h5d == r_count_20_io_out ? io_r_93_b : _GEN_6182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6184 = 9'h5e == r_count_20_io_out ? io_r_94_b : _GEN_6183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6185 = 9'h5f == r_count_20_io_out ? io_r_95_b : _GEN_6184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6186 = 9'h60 == r_count_20_io_out ? io_r_96_b : _GEN_6185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6187 = 9'h61 == r_count_20_io_out ? io_r_97_b : _GEN_6186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6188 = 9'h62 == r_count_20_io_out ? io_r_98_b : _GEN_6187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6189 = 9'h63 == r_count_20_io_out ? io_r_99_b : _GEN_6188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6190 = 9'h64 == r_count_20_io_out ? io_r_100_b : _GEN_6189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6191 = 9'h65 == r_count_20_io_out ? io_r_101_b : _GEN_6190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6192 = 9'h66 == r_count_20_io_out ? io_r_102_b : _GEN_6191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6193 = 9'h67 == r_count_20_io_out ? io_r_103_b : _GEN_6192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6194 = 9'h68 == r_count_20_io_out ? io_r_104_b : _GEN_6193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6195 = 9'h69 == r_count_20_io_out ? io_r_105_b : _GEN_6194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6196 = 9'h6a == r_count_20_io_out ? io_r_106_b : _GEN_6195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6197 = 9'h6b == r_count_20_io_out ? io_r_107_b : _GEN_6196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6198 = 9'h6c == r_count_20_io_out ? io_r_108_b : _GEN_6197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6199 = 9'h6d == r_count_20_io_out ? io_r_109_b : _GEN_6198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6200 = 9'h6e == r_count_20_io_out ? io_r_110_b : _GEN_6199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6201 = 9'h6f == r_count_20_io_out ? io_r_111_b : _GEN_6200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6202 = 9'h70 == r_count_20_io_out ? io_r_112_b : _GEN_6201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6203 = 9'h71 == r_count_20_io_out ? io_r_113_b : _GEN_6202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6204 = 9'h72 == r_count_20_io_out ? io_r_114_b : _GEN_6203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6205 = 9'h73 == r_count_20_io_out ? io_r_115_b : _GEN_6204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6206 = 9'h74 == r_count_20_io_out ? io_r_116_b : _GEN_6205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6207 = 9'h75 == r_count_20_io_out ? io_r_117_b : _GEN_6206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6208 = 9'h76 == r_count_20_io_out ? io_r_118_b : _GEN_6207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6209 = 9'h77 == r_count_20_io_out ? io_r_119_b : _GEN_6208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6210 = 9'h78 == r_count_20_io_out ? io_r_120_b : _GEN_6209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6211 = 9'h79 == r_count_20_io_out ? io_r_121_b : _GEN_6210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6212 = 9'h7a == r_count_20_io_out ? io_r_122_b : _GEN_6211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6213 = 9'h7b == r_count_20_io_out ? io_r_123_b : _GEN_6212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6214 = 9'h7c == r_count_20_io_out ? io_r_124_b : _GEN_6213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6215 = 9'h7d == r_count_20_io_out ? io_r_125_b : _GEN_6214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6216 = 9'h7e == r_count_20_io_out ? io_r_126_b : _GEN_6215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6217 = 9'h7f == r_count_20_io_out ? io_r_127_b : _GEN_6216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6218 = 9'h80 == r_count_20_io_out ? io_r_128_b : _GEN_6217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6219 = 9'h81 == r_count_20_io_out ? io_r_129_b : _GEN_6218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6220 = 9'h82 == r_count_20_io_out ? io_r_130_b : _GEN_6219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6221 = 9'h83 == r_count_20_io_out ? io_r_131_b : _GEN_6220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6222 = 9'h84 == r_count_20_io_out ? io_r_132_b : _GEN_6221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6223 = 9'h85 == r_count_20_io_out ? io_r_133_b : _GEN_6222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6224 = 9'h86 == r_count_20_io_out ? io_r_134_b : _GEN_6223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6225 = 9'h87 == r_count_20_io_out ? io_r_135_b : _GEN_6224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6226 = 9'h88 == r_count_20_io_out ? io_r_136_b : _GEN_6225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6227 = 9'h89 == r_count_20_io_out ? io_r_137_b : _GEN_6226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6228 = 9'h8a == r_count_20_io_out ? io_r_138_b : _GEN_6227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6229 = 9'h8b == r_count_20_io_out ? io_r_139_b : _GEN_6228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6230 = 9'h8c == r_count_20_io_out ? io_r_140_b : _GEN_6229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6231 = 9'h8d == r_count_20_io_out ? io_r_141_b : _GEN_6230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6232 = 9'h8e == r_count_20_io_out ? io_r_142_b : _GEN_6231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6233 = 9'h8f == r_count_20_io_out ? io_r_143_b : _GEN_6232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6234 = 9'h90 == r_count_20_io_out ? io_r_144_b : _GEN_6233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6235 = 9'h91 == r_count_20_io_out ? io_r_145_b : _GEN_6234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6236 = 9'h92 == r_count_20_io_out ? io_r_146_b : _GEN_6235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6237 = 9'h93 == r_count_20_io_out ? io_r_147_b : _GEN_6236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6238 = 9'h94 == r_count_20_io_out ? io_r_148_b : _GEN_6237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6239 = 9'h95 == r_count_20_io_out ? io_r_149_b : _GEN_6238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6240 = 9'h96 == r_count_20_io_out ? io_r_150_b : _GEN_6239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6241 = 9'h97 == r_count_20_io_out ? io_r_151_b : _GEN_6240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6242 = 9'h98 == r_count_20_io_out ? io_r_152_b : _GEN_6241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6243 = 9'h99 == r_count_20_io_out ? io_r_153_b : _GEN_6242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6244 = 9'h9a == r_count_20_io_out ? io_r_154_b : _GEN_6243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6245 = 9'h9b == r_count_20_io_out ? io_r_155_b : _GEN_6244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6246 = 9'h9c == r_count_20_io_out ? io_r_156_b : _GEN_6245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6247 = 9'h9d == r_count_20_io_out ? io_r_157_b : _GEN_6246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6248 = 9'h9e == r_count_20_io_out ? io_r_158_b : _GEN_6247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6249 = 9'h9f == r_count_20_io_out ? io_r_159_b : _GEN_6248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6250 = 9'ha0 == r_count_20_io_out ? io_r_160_b : _GEN_6249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6251 = 9'ha1 == r_count_20_io_out ? io_r_161_b : _GEN_6250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6252 = 9'ha2 == r_count_20_io_out ? io_r_162_b : _GEN_6251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6253 = 9'ha3 == r_count_20_io_out ? io_r_163_b : _GEN_6252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6254 = 9'ha4 == r_count_20_io_out ? io_r_164_b : _GEN_6253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6255 = 9'ha5 == r_count_20_io_out ? io_r_165_b : _GEN_6254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6256 = 9'ha6 == r_count_20_io_out ? io_r_166_b : _GEN_6255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6257 = 9'ha7 == r_count_20_io_out ? io_r_167_b : _GEN_6256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6258 = 9'ha8 == r_count_20_io_out ? io_r_168_b : _GEN_6257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6259 = 9'ha9 == r_count_20_io_out ? io_r_169_b : _GEN_6258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6260 = 9'haa == r_count_20_io_out ? io_r_170_b : _GEN_6259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6261 = 9'hab == r_count_20_io_out ? io_r_171_b : _GEN_6260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6262 = 9'hac == r_count_20_io_out ? io_r_172_b : _GEN_6261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6263 = 9'had == r_count_20_io_out ? io_r_173_b : _GEN_6262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6264 = 9'hae == r_count_20_io_out ? io_r_174_b : _GEN_6263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6265 = 9'haf == r_count_20_io_out ? io_r_175_b : _GEN_6264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6266 = 9'hb0 == r_count_20_io_out ? io_r_176_b : _GEN_6265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6267 = 9'hb1 == r_count_20_io_out ? io_r_177_b : _GEN_6266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6268 = 9'hb2 == r_count_20_io_out ? io_r_178_b : _GEN_6267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6269 = 9'hb3 == r_count_20_io_out ? io_r_179_b : _GEN_6268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6270 = 9'hb4 == r_count_20_io_out ? io_r_180_b : _GEN_6269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6271 = 9'hb5 == r_count_20_io_out ? io_r_181_b : _GEN_6270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6272 = 9'hb6 == r_count_20_io_out ? io_r_182_b : _GEN_6271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6273 = 9'hb7 == r_count_20_io_out ? io_r_183_b : _GEN_6272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6274 = 9'hb8 == r_count_20_io_out ? io_r_184_b : _GEN_6273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6275 = 9'hb9 == r_count_20_io_out ? io_r_185_b : _GEN_6274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6276 = 9'hba == r_count_20_io_out ? io_r_186_b : _GEN_6275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6277 = 9'hbb == r_count_20_io_out ? io_r_187_b : _GEN_6276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6278 = 9'hbc == r_count_20_io_out ? io_r_188_b : _GEN_6277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6279 = 9'hbd == r_count_20_io_out ? io_r_189_b : _GEN_6278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6280 = 9'hbe == r_count_20_io_out ? io_r_190_b : _GEN_6279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6281 = 9'hbf == r_count_20_io_out ? io_r_191_b : _GEN_6280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6282 = 9'hc0 == r_count_20_io_out ? io_r_192_b : _GEN_6281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6283 = 9'hc1 == r_count_20_io_out ? io_r_193_b : _GEN_6282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6284 = 9'hc2 == r_count_20_io_out ? io_r_194_b : _GEN_6283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6285 = 9'hc3 == r_count_20_io_out ? io_r_195_b : _GEN_6284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6286 = 9'hc4 == r_count_20_io_out ? io_r_196_b : _GEN_6285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6287 = 9'hc5 == r_count_20_io_out ? io_r_197_b : _GEN_6286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6288 = 9'hc6 == r_count_20_io_out ? io_r_198_b : _GEN_6287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6289 = 9'hc7 == r_count_20_io_out ? io_r_199_b : _GEN_6288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6290 = 9'hc8 == r_count_20_io_out ? io_r_200_b : _GEN_6289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6291 = 9'hc9 == r_count_20_io_out ? io_r_201_b : _GEN_6290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6292 = 9'hca == r_count_20_io_out ? io_r_202_b : _GEN_6291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6293 = 9'hcb == r_count_20_io_out ? io_r_203_b : _GEN_6292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6294 = 9'hcc == r_count_20_io_out ? io_r_204_b : _GEN_6293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6295 = 9'hcd == r_count_20_io_out ? io_r_205_b : _GEN_6294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6296 = 9'hce == r_count_20_io_out ? io_r_206_b : _GEN_6295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6297 = 9'hcf == r_count_20_io_out ? io_r_207_b : _GEN_6296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6298 = 9'hd0 == r_count_20_io_out ? io_r_208_b : _GEN_6297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6299 = 9'hd1 == r_count_20_io_out ? io_r_209_b : _GEN_6298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6300 = 9'hd2 == r_count_20_io_out ? io_r_210_b : _GEN_6299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6301 = 9'hd3 == r_count_20_io_out ? io_r_211_b : _GEN_6300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6302 = 9'hd4 == r_count_20_io_out ? io_r_212_b : _GEN_6301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6303 = 9'hd5 == r_count_20_io_out ? io_r_213_b : _GEN_6302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6304 = 9'hd6 == r_count_20_io_out ? io_r_214_b : _GEN_6303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6305 = 9'hd7 == r_count_20_io_out ? io_r_215_b : _GEN_6304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6306 = 9'hd8 == r_count_20_io_out ? io_r_216_b : _GEN_6305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6307 = 9'hd9 == r_count_20_io_out ? io_r_217_b : _GEN_6306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6308 = 9'hda == r_count_20_io_out ? io_r_218_b : _GEN_6307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6309 = 9'hdb == r_count_20_io_out ? io_r_219_b : _GEN_6308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6310 = 9'hdc == r_count_20_io_out ? io_r_220_b : _GEN_6309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6311 = 9'hdd == r_count_20_io_out ? io_r_221_b : _GEN_6310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6312 = 9'hde == r_count_20_io_out ? io_r_222_b : _GEN_6311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6313 = 9'hdf == r_count_20_io_out ? io_r_223_b : _GEN_6312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6314 = 9'he0 == r_count_20_io_out ? io_r_224_b : _GEN_6313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6315 = 9'he1 == r_count_20_io_out ? io_r_225_b : _GEN_6314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6316 = 9'he2 == r_count_20_io_out ? io_r_226_b : _GEN_6315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6317 = 9'he3 == r_count_20_io_out ? io_r_227_b : _GEN_6316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6318 = 9'he4 == r_count_20_io_out ? io_r_228_b : _GEN_6317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6319 = 9'he5 == r_count_20_io_out ? io_r_229_b : _GEN_6318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6320 = 9'he6 == r_count_20_io_out ? io_r_230_b : _GEN_6319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6321 = 9'he7 == r_count_20_io_out ? io_r_231_b : _GEN_6320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6322 = 9'he8 == r_count_20_io_out ? io_r_232_b : _GEN_6321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6323 = 9'he9 == r_count_20_io_out ? io_r_233_b : _GEN_6322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6324 = 9'hea == r_count_20_io_out ? io_r_234_b : _GEN_6323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6325 = 9'heb == r_count_20_io_out ? io_r_235_b : _GEN_6324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6326 = 9'hec == r_count_20_io_out ? io_r_236_b : _GEN_6325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6327 = 9'hed == r_count_20_io_out ? io_r_237_b : _GEN_6326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6328 = 9'hee == r_count_20_io_out ? io_r_238_b : _GEN_6327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6329 = 9'hef == r_count_20_io_out ? io_r_239_b : _GEN_6328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6330 = 9'hf0 == r_count_20_io_out ? io_r_240_b : _GEN_6329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6331 = 9'hf1 == r_count_20_io_out ? io_r_241_b : _GEN_6330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6332 = 9'hf2 == r_count_20_io_out ? io_r_242_b : _GEN_6331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6333 = 9'hf3 == r_count_20_io_out ? io_r_243_b : _GEN_6332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6334 = 9'hf4 == r_count_20_io_out ? io_r_244_b : _GEN_6333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6335 = 9'hf5 == r_count_20_io_out ? io_r_245_b : _GEN_6334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6336 = 9'hf6 == r_count_20_io_out ? io_r_246_b : _GEN_6335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6337 = 9'hf7 == r_count_20_io_out ? io_r_247_b : _GEN_6336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6338 = 9'hf8 == r_count_20_io_out ? io_r_248_b : _GEN_6337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6339 = 9'hf9 == r_count_20_io_out ? io_r_249_b : _GEN_6338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6340 = 9'hfa == r_count_20_io_out ? io_r_250_b : _GEN_6339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6341 = 9'hfb == r_count_20_io_out ? io_r_251_b : _GEN_6340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6342 = 9'hfc == r_count_20_io_out ? io_r_252_b : _GEN_6341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6343 = 9'hfd == r_count_20_io_out ? io_r_253_b : _GEN_6342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6344 = 9'hfe == r_count_20_io_out ? io_r_254_b : _GEN_6343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6345 = 9'hff == r_count_20_io_out ? io_r_255_b : _GEN_6344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6346 = 9'h100 == r_count_20_io_out ? io_r_256_b : _GEN_6345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6347 = 9'h101 == r_count_20_io_out ? io_r_257_b : _GEN_6346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6348 = 9'h102 == r_count_20_io_out ? io_r_258_b : _GEN_6347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6349 = 9'h103 == r_count_20_io_out ? io_r_259_b : _GEN_6348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6350 = 9'h104 == r_count_20_io_out ? io_r_260_b : _GEN_6349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6351 = 9'h105 == r_count_20_io_out ? io_r_261_b : _GEN_6350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6352 = 9'h106 == r_count_20_io_out ? io_r_262_b : _GEN_6351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6353 = 9'h107 == r_count_20_io_out ? io_r_263_b : _GEN_6352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6354 = 9'h108 == r_count_20_io_out ? io_r_264_b : _GEN_6353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6355 = 9'h109 == r_count_20_io_out ? io_r_265_b : _GEN_6354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6356 = 9'h10a == r_count_20_io_out ? io_r_266_b : _GEN_6355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6357 = 9'h10b == r_count_20_io_out ? io_r_267_b : _GEN_6356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6358 = 9'h10c == r_count_20_io_out ? io_r_268_b : _GEN_6357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6359 = 9'h10d == r_count_20_io_out ? io_r_269_b : _GEN_6358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6360 = 9'h10e == r_count_20_io_out ? io_r_270_b : _GEN_6359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6361 = 9'h10f == r_count_20_io_out ? io_r_271_b : _GEN_6360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6362 = 9'h110 == r_count_20_io_out ? io_r_272_b : _GEN_6361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6363 = 9'h111 == r_count_20_io_out ? io_r_273_b : _GEN_6362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6364 = 9'h112 == r_count_20_io_out ? io_r_274_b : _GEN_6363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6365 = 9'h113 == r_count_20_io_out ? io_r_275_b : _GEN_6364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6366 = 9'h114 == r_count_20_io_out ? io_r_276_b : _GEN_6365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6367 = 9'h115 == r_count_20_io_out ? io_r_277_b : _GEN_6366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6368 = 9'h116 == r_count_20_io_out ? io_r_278_b : _GEN_6367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6369 = 9'h117 == r_count_20_io_out ? io_r_279_b : _GEN_6368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6370 = 9'h118 == r_count_20_io_out ? io_r_280_b : _GEN_6369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6371 = 9'h119 == r_count_20_io_out ? io_r_281_b : _GEN_6370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6372 = 9'h11a == r_count_20_io_out ? io_r_282_b : _GEN_6371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6373 = 9'h11b == r_count_20_io_out ? io_r_283_b : _GEN_6372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6374 = 9'h11c == r_count_20_io_out ? io_r_284_b : _GEN_6373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6375 = 9'h11d == r_count_20_io_out ? io_r_285_b : _GEN_6374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6376 = 9'h11e == r_count_20_io_out ? io_r_286_b : _GEN_6375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6377 = 9'h11f == r_count_20_io_out ? io_r_287_b : _GEN_6376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6378 = 9'h120 == r_count_20_io_out ? io_r_288_b : _GEN_6377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6379 = 9'h121 == r_count_20_io_out ? io_r_289_b : _GEN_6378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6380 = 9'h122 == r_count_20_io_out ? io_r_290_b : _GEN_6379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6381 = 9'h123 == r_count_20_io_out ? io_r_291_b : _GEN_6380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6382 = 9'h124 == r_count_20_io_out ? io_r_292_b : _GEN_6381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6383 = 9'h125 == r_count_20_io_out ? io_r_293_b : _GEN_6382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6384 = 9'h126 == r_count_20_io_out ? io_r_294_b : _GEN_6383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6385 = 9'h127 == r_count_20_io_out ? io_r_295_b : _GEN_6384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6386 = 9'h128 == r_count_20_io_out ? io_r_296_b : _GEN_6385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6387 = 9'h129 == r_count_20_io_out ? io_r_297_b : _GEN_6386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6388 = 9'h12a == r_count_20_io_out ? io_r_298_b : _GEN_6387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6391 = 9'h1 == r_count_21_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6392 = 9'h2 == r_count_21_io_out ? io_r_2_b : _GEN_6391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6393 = 9'h3 == r_count_21_io_out ? io_r_3_b : _GEN_6392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6394 = 9'h4 == r_count_21_io_out ? io_r_4_b : _GEN_6393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6395 = 9'h5 == r_count_21_io_out ? io_r_5_b : _GEN_6394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6396 = 9'h6 == r_count_21_io_out ? io_r_6_b : _GEN_6395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6397 = 9'h7 == r_count_21_io_out ? io_r_7_b : _GEN_6396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6398 = 9'h8 == r_count_21_io_out ? io_r_8_b : _GEN_6397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6399 = 9'h9 == r_count_21_io_out ? io_r_9_b : _GEN_6398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6400 = 9'ha == r_count_21_io_out ? io_r_10_b : _GEN_6399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6401 = 9'hb == r_count_21_io_out ? io_r_11_b : _GEN_6400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6402 = 9'hc == r_count_21_io_out ? io_r_12_b : _GEN_6401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6403 = 9'hd == r_count_21_io_out ? io_r_13_b : _GEN_6402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6404 = 9'he == r_count_21_io_out ? io_r_14_b : _GEN_6403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6405 = 9'hf == r_count_21_io_out ? io_r_15_b : _GEN_6404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6406 = 9'h10 == r_count_21_io_out ? io_r_16_b : _GEN_6405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6407 = 9'h11 == r_count_21_io_out ? io_r_17_b : _GEN_6406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6408 = 9'h12 == r_count_21_io_out ? io_r_18_b : _GEN_6407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6409 = 9'h13 == r_count_21_io_out ? io_r_19_b : _GEN_6408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6410 = 9'h14 == r_count_21_io_out ? io_r_20_b : _GEN_6409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6411 = 9'h15 == r_count_21_io_out ? io_r_21_b : _GEN_6410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6412 = 9'h16 == r_count_21_io_out ? io_r_22_b : _GEN_6411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6413 = 9'h17 == r_count_21_io_out ? io_r_23_b : _GEN_6412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6414 = 9'h18 == r_count_21_io_out ? io_r_24_b : _GEN_6413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6415 = 9'h19 == r_count_21_io_out ? io_r_25_b : _GEN_6414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6416 = 9'h1a == r_count_21_io_out ? io_r_26_b : _GEN_6415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6417 = 9'h1b == r_count_21_io_out ? io_r_27_b : _GEN_6416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6418 = 9'h1c == r_count_21_io_out ? io_r_28_b : _GEN_6417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6419 = 9'h1d == r_count_21_io_out ? io_r_29_b : _GEN_6418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6420 = 9'h1e == r_count_21_io_out ? io_r_30_b : _GEN_6419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6421 = 9'h1f == r_count_21_io_out ? io_r_31_b : _GEN_6420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6422 = 9'h20 == r_count_21_io_out ? io_r_32_b : _GEN_6421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6423 = 9'h21 == r_count_21_io_out ? io_r_33_b : _GEN_6422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6424 = 9'h22 == r_count_21_io_out ? io_r_34_b : _GEN_6423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6425 = 9'h23 == r_count_21_io_out ? io_r_35_b : _GEN_6424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6426 = 9'h24 == r_count_21_io_out ? io_r_36_b : _GEN_6425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6427 = 9'h25 == r_count_21_io_out ? io_r_37_b : _GEN_6426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6428 = 9'h26 == r_count_21_io_out ? io_r_38_b : _GEN_6427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6429 = 9'h27 == r_count_21_io_out ? io_r_39_b : _GEN_6428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6430 = 9'h28 == r_count_21_io_out ? io_r_40_b : _GEN_6429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6431 = 9'h29 == r_count_21_io_out ? io_r_41_b : _GEN_6430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6432 = 9'h2a == r_count_21_io_out ? io_r_42_b : _GEN_6431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6433 = 9'h2b == r_count_21_io_out ? io_r_43_b : _GEN_6432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6434 = 9'h2c == r_count_21_io_out ? io_r_44_b : _GEN_6433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6435 = 9'h2d == r_count_21_io_out ? io_r_45_b : _GEN_6434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6436 = 9'h2e == r_count_21_io_out ? io_r_46_b : _GEN_6435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6437 = 9'h2f == r_count_21_io_out ? io_r_47_b : _GEN_6436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6438 = 9'h30 == r_count_21_io_out ? io_r_48_b : _GEN_6437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6439 = 9'h31 == r_count_21_io_out ? io_r_49_b : _GEN_6438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6440 = 9'h32 == r_count_21_io_out ? io_r_50_b : _GEN_6439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6441 = 9'h33 == r_count_21_io_out ? io_r_51_b : _GEN_6440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6442 = 9'h34 == r_count_21_io_out ? io_r_52_b : _GEN_6441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6443 = 9'h35 == r_count_21_io_out ? io_r_53_b : _GEN_6442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6444 = 9'h36 == r_count_21_io_out ? io_r_54_b : _GEN_6443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6445 = 9'h37 == r_count_21_io_out ? io_r_55_b : _GEN_6444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6446 = 9'h38 == r_count_21_io_out ? io_r_56_b : _GEN_6445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6447 = 9'h39 == r_count_21_io_out ? io_r_57_b : _GEN_6446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6448 = 9'h3a == r_count_21_io_out ? io_r_58_b : _GEN_6447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6449 = 9'h3b == r_count_21_io_out ? io_r_59_b : _GEN_6448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6450 = 9'h3c == r_count_21_io_out ? io_r_60_b : _GEN_6449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6451 = 9'h3d == r_count_21_io_out ? io_r_61_b : _GEN_6450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6452 = 9'h3e == r_count_21_io_out ? io_r_62_b : _GEN_6451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6453 = 9'h3f == r_count_21_io_out ? io_r_63_b : _GEN_6452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6454 = 9'h40 == r_count_21_io_out ? io_r_64_b : _GEN_6453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6455 = 9'h41 == r_count_21_io_out ? io_r_65_b : _GEN_6454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6456 = 9'h42 == r_count_21_io_out ? io_r_66_b : _GEN_6455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6457 = 9'h43 == r_count_21_io_out ? io_r_67_b : _GEN_6456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6458 = 9'h44 == r_count_21_io_out ? io_r_68_b : _GEN_6457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6459 = 9'h45 == r_count_21_io_out ? io_r_69_b : _GEN_6458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6460 = 9'h46 == r_count_21_io_out ? io_r_70_b : _GEN_6459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6461 = 9'h47 == r_count_21_io_out ? io_r_71_b : _GEN_6460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6462 = 9'h48 == r_count_21_io_out ? io_r_72_b : _GEN_6461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6463 = 9'h49 == r_count_21_io_out ? io_r_73_b : _GEN_6462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6464 = 9'h4a == r_count_21_io_out ? io_r_74_b : _GEN_6463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6465 = 9'h4b == r_count_21_io_out ? io_r_75_b : _GEN_6464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6466 = 9'h4c == r_count_21_io_out ? io_r_76_b : _GEN_6465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6467 = 9'h4d == r_count_21_io_out ? io_r_77_b : _GEN_6466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6468 = 9'h4e == r_count_21_io_out ? io_r_78_b : _GEN_6467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6469 = 9'h4f == r_count_21_io_out ? io_r_79_b : _GEN_6468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6470 = 9'h50 == r_count_21_io_out ? io_r_80_b : _GEN_6469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6471 = 9'h51 == r_count_21_io_out ? io_r_81_b : _GEN_6470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6472 = 9'h52 == r_count_21_io_out ? io_r_82_b : _GEN_6471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6473 = 9'h53 == r_count_21_io_out ? io_r_83_b : _GEN_6472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6474 = 9'h54 == r_count_21_io_out ? io_r_84_b : _GEN_6473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6475 = 9'h55 == r_count_21_io_out ? io_r_85_b : _GEN_6474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6476 = 9'h56 == r_count_21_io_out ? io_r_86_b : _GEN_6475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6477 = 9'h57 == r_count_21_io_out ? io_r_87_b : _GEN_6476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6478 = 9'h58 == r_count_21_io_out ? io_r_88_b : _GEN_6477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6479 = 9'h59 == r_count_21_io_out ? io_r_89_b : _GEN_6478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6480 = 9'h5a == r_count_21_io_out ? io_r_90_b : _GEN_6479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6481 = 9'h5b == r_count_21_io_out ? io_r_91_b : _GEN_6480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6482 = 9'h5c == r_count_21_io_out ? io_r_92_b : _GEN_6481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6483 = 9'h5d == r_count_21_io_out ? io_r_93_b : _GEN_6482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6484 = 9'h5e == r_count_21_io_out ? io_r_94_b : _GEN_6483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6485 = 9'h5f == r_count_21_io_out ? io_r_95_b : _GEN_6484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6486 = 9'h60 == r_count_21_io_out ? io_r_96_b : _GEN_6485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6487 = 9'h61 == r_count_21_io_out ? io_r_97_b : _GEN_6486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6488 = 9'h62 == r_count_21_io_out ? io_r_98_b : _GEN_6487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6489 = 9'h63 == r_count_21_io_out ? io_r_99_b : _GEN_6488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6490 = 9'h64 == r_count_21_io_out ? io_r_100_b : _GEN_6489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6491 = 9'h65 == r_count_21_io_out ? io_r_101_b : _GEN_6490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6492 = 9'h66 == r_count_21_io_out ? io_r_102_b : _GEN_6491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6493 = 9'h67 == r_count_21_io_out ? io_r_103_b : _GEN_6492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6494 = 9'h68 == r_count_21_io_out ? io_r_104_b : _GEN_6493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6495 = 9'h69 == r_count_21_io_out ? io_r_105_b : _GEN_6494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6496 = 9'h6a == r_count_21_io_out ? io_r_106_b : _GEN_6495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6497 = 9'h6b == r_count_21_io_out ? io_r_107_b : _GEN_6496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6498 = 9'h6c == r_count_21_io_out ? io_r_108_b : _GEN_6497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6499 = 9'h6d == r_count_21_io_out ? io_r_109_b : _GEN_6498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6500 = 9'h6e == r_count_21_io_out ? io_r_110_b : _GEN_6499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6501 = 9'h6f == r_count_21_io_out ? io_r_111_b : _GEN_6500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6502 = 9'h70 == r_count_21_io_out ? io_r_112_b : _GEN_6501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6503 = 9'h71 == r_count_21_io_out ? io_r_113_b : _GEN_6502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6504 = 9'h72 == r_count_21_io_out ? io_r_114_b : _GEN_6503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6505 = 9'h73 == r_count_21_io_out ? io_r_115_b : _GEN_6504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6506 = 9'h74 == r_count_21_io_out ? io_r_116_b : _GEN_6505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6507 = 9'h75 == r_count_21_io_out ? io_r_117_b : _GEN_6506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6508 = 9'h76 == r_count_21_io_out ? io_r_118_b : _GEN_6507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6509 = 9'h77 == r_count_21_io_out ? io_r_119_b : _GEN_6508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6510 = 9'h78 == r_count_21_io_out ? io_r_120_b : _GEN_6509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6511 = 9'h79 == r_count_21_io_out ? io_r_121_b : _GEN_6510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6512 = 9'h7a == r_count_21_io_out ? io_r_122_b : _GEN_6511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6513 = 9'h7b == r_count_21_io_out ? io_r_123_b : _GEN_6512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6514 = 9'h7c == r_count_21_io_out ? io_r_124_b : _GEN_6513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6515 = 9'h7d == r_count_21_io_out ? io_r_125_b : _GEN_6514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6516 = 9'h7e == r_count_21_io_out ? io_r_126_b : _GEN_6515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6517 = 9'h7f == r_count_21_io_out ? io_r_127_b : _GEN_6516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6518 = 9'h80 == r_count_21_io_out ? io_r_128_b : _GEN_6517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6519 = 9'h81 == r_count_21_io_out ? io_r_129_b : _GEN_6518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6520 = 9'h82 == r_count_21_io_out ? io_r_130_b : _GEN_6519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6521 = 9'h83 == r_count_21_io_out ? io_r_131_b : _GEN_6520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6522 = 9'h84 == r_count_21_io_out ? io_r_132_b : _GEN_6521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6523 = 9'h85 == r_count_21_io_out ? io_r_133_b : _GEN_6522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6524 = 9'h86 == r_count_21_io_out ? io_r_134_b : _GEN_6523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6525 = 9'h87 == r_count_21_io_out ? io_r_135_b : _GEN_6524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6526 = 9'h88 == r_count_21_io_out ? io_r_136_b : _GEN_6525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6527 = 9'h89 == r_count_21_io_out ? io_r_137_b : _GEN_6526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6528 = 9'h8a == r_count_21_io_out ? io_r_138_b : _GEN_6527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6529 = 9'h8b == r_count_21_io_out ? io_r_139_b : _GEN_6528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6530 = 9'h8c == r_count_21_io_out ? io_r_140_b : _GEN_6529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6531 = 9'h8d == r_count_21_io_out ? io_r_141_b : _GEN_6530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6532 = 9'h8e == r_count_21_io_out ? io_r_142_b : _GEN_6531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6533 = 9'h8f == r_count_21_io_out ? io_r_143_b : _GEN_6532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6534 = 9'h90 == r_count_21_io_out ? io_r_144_b : _GEN_6533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6535 = 9'h91 == r_count_21_io_out ? io_r_145_b : _GEN_6534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6536 = 9'h92 == r_count_21_io_out ? io_r_146_b : _GEN_6535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6537 = 9'h93 == r_count_21_io_out ? io_r_147_b : _GEN_6536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6538 = 9'h94 == r_count_21_io_out ? io_r_148_b : _GEN_6537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6539 = 9'h95 == r_count_21_io_out ? io_r_149_b : _GEN_6538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6540 = 9'h96 == r_count_21_io_out ? io_r_150_b : _GEN_6539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6541 = 9'h97 == r_count_21_io_out ? io_r_151_b : _GEN_6540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6542 = 9'h98 == r_count_21_io_out ? io_r_152_b : _GEN_6541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6543 = 9'h99 == r_count_21_io_out ? io_r_153_b : _GEN_6542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6544 = 9'h9a == r_count_21_io_out ? io_r_154_b : _GEN_6543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6545 = 9'h9b == r_count_21_io_out ? io_r_155_b : _GEN_6544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6546 = 9'h9c == r_count_21_io_out ? io_r_156_b : _GEN_6545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6547 = 9'h9d == r_count_21_io_out ? io_r_157_b : _GEN_6546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6548 = 9'h9e == r_count_21_io_out ? io_r_158_b : _GEN_6547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6549 = 9'h9f == r_count_21_io_out ? io_r_159_b : _GEN_6548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6550 = 9'ha0 == r_count_21_io_out ? io_r_160_b : _GEN_6549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6551 = 9'ha1 == r_count_21_io_out ? io_r_161_b : _GEN_6550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6552 = 9'ha2 == r_count_21_io_out ? io_r_162_b : _GEN_6551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6553 = 9'ha3 == r_count_21_io_out ? io_r_163_b : _GEN_6552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6554 = 9'ha4 == r_count_21_io_out ? io_r_164_b : _GEN_6553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6555 = 9'ha5 == r_count_21_io_out ? io_r_165_b : _GEN_6554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6556 = 9'ha6 == r_count_21_io_out ? io_r_166_b : _GEN_6555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6557 = 9'ha7 == r_count_21_io_out ? io_r_167_b : _GEN_6556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6558 = 9'ha8 == r_count_21_io_out ? io_r_168_b : _GEN_6557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6559 = 9'ha9 == r_count_21_io_out ? io_r_169_b : _GEN_6558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6560 = 9'haa == r_count_21_io_out ? io_r_170_b : _GEN_6559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6561 = 9'hab == r_count_21_io_out ? io_r_171_b : _GEN_6560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6562 = 9'hac == r_count_21_io_out ? io_r_172_b : _GEN_6561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6563 = 9'had == r_count_21_io_out ? io_r_173_b : _GEN_6562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6564 = 9'hae == r_count_21_io_out ? io_r_174_b : _GEN_6563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6565 = 9'haf == r_count_21_io_out ? io_r_175_b : _GEN_6564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6566 = 9'hb0 == r_count_21_io_out ? io_r_176_b : _GEN_6565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6567 = 9'hb1 == r_count_21_io_out ? io_r_177_b : _GEN_6566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6568 = 9'hb2 == r_count_21_io_out ? io_r_178_b : _GEN_6567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6569 = 9'hb3 == r_count_21_io_out ? io_r_179_b : _GEN_6568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6570 = 9'hb4 == r_count_21_io_out ? io_r_180_b : _GEN_6569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6571 = 9'hb5 == r_count_21_io_out ? io_r_181_b : _GEN_6570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6572 = 9'hb6 == r_count_21_io_out ? io_r_182_b : _GEN_6571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6573 = 9'hb7 == r_count_21_io_out ? io_r_183_b : _GEN_6572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6574 = 9'hb8 == r_count_21_io_out ? io_r_184_b : _GEN_6573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6575 = 9'hb9 == r_count_21_io_out ? io_r_185_b : _GEN_6574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6576 = 9'hba == r_count_21_io_out ? io_r_186_b : _GEN_6575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6577 = 9'hbb == r_count_21_io_out ? io_r_187_b : _GEN_6576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6578 = 9'hbc == r_count_21_io_out ? io_r_188_b : _GEN_6577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6579 = 9'hbd == r_count_21_io_out ? io_r_189_b : _GEN_6578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6580 = 9'hbe == r_count_21_io_out ? io_r_190_b : _GEN_6579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6581 = 9'hbf == r_count_21_io_out ? io_r_191_b : _GEN_6580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6582 = 9'hc0 == r_count_21_io_out ? io_r_192_b : _GEN_6581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6583 = 9'hc1 == r_count_21_io_out ? io_r_193_b : _GEN_6582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6584 = 9'hc2 == r_count_21_io_out ? io_r_194_b : _GEN_6583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6585 = 9'hc3 == r_count_21_io_out ? io_r_195_b : _GEN_6584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6586 = 9'hc4 == r_count_21_io_out ? io_r_196_b : _GEN_6585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6587 = 9'hc5 == r_count_21_io_out ? io_r_197_b : _GEN_6586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6588 = 9'hc6 == r_count_21_io_out ? io_r_198_b : _GEN_6587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6589 = 9'hc7 == r_count_21_io_out ? io_r_199_b : _GEN_6588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6590 = 9'hc8 == r_count_21_io_out ? io_r_200_b : _GEN_6589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6591 = 9'hc9 == r_count_21_io_out ? io_r_201_b : _GEN_6590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6592 = 9'hca == r_count_21_io_out ? io_r_202_b : _GEN_6591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6593 = 9'hcb == r_count_21_io_out ? io_r_203_b : _GEN_6592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6594 = 9'hcc == r_count_21_io_out ? io_r_204_b : _GEN_6593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6595 = 9'hcd == r_count_21_io_out ? io_r_205_b : _GEN_6594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6596 = 9'hce == r_count_21_io_out ? io_r_206_b : _GEN_6595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6597 = 9'hcf == r_count_21_io_out ? io_r_207_b : _GEN_6596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6598 = 9'hd0 == r_count_21_io_out ? io_r_208_b : _GEN_6597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6599 = 9'hd1 == r_count_21_io_out ? io_r_209_b : _GEN_6598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6600 = 9'hd2 == r_count_21_io_out ? io_r_210_b : _GEN_6599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6601 = 9'hd3 == r_count_21_io_out ? io_r_211_b : _GEN_6600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6602 = 9'hd4 == r_count_21_io_out ? io_r_212_b : _GEN_6601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6603 = 9'hd5 == r_count_21_io_out ? io_r_213_b : _GEN_6602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6604 = 9'hd6 == r_count_21_io_out ? io_r_214_b : _GEN_6603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6605 = 9'hd7 == r_count_21_io_out ? io_r_215_b : _GEN_6604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6606 = 9'hd8 == r_count_21_io_out ? io_r_216_b : _GEN_6605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6607 = 9'hd9 == r_count_21_io_out ? io_r_217_b : _GEN_6606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6608 = 9'hda == r_count_21_io_out ? io_r_218_b : _GEN_6607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6609 = 9'hdb == r_count_21_io_out ? io_r_219_b : _GEN_6608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6610 = 9'hdc == r_count_21_io_out ? io_r_220_b : _GEN_6609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6611 = 9'hdd == r_count_21_io_out ? io_r_221_b : _GEN_6610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6612 = 9'hde == r_count_21_io_out ? io_r_222_b : _GEN_6611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6613 = 9'hdf == r_count_21_io_out ? io_r_223_b : _GEN_6612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6614 = 9'he0 == r_count_21_io_out ? io_r_224_b : _GEN_6613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6615 = 9'he1 == r_count_21_io_out ? io_r_225_b : _GEN_6614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6616 = 9'he2 == r_count_21_io_out ? io_r_226_b : _GEN_6615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6617 = 9'he3 == r_count_21_io_out ? io_r_227_b : _GEN_6616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6618 = 9'he4 == r_count_21_io_out ? io_r_228_b : _GEN_6617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6619 = 9'he5 == r_count_21_io_out ? io_r_229_b : _GEN_6618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6620 = 9'he6 == r_count_21_io_out ? io_r_230_b : _GEN_6619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6621 = 9'he7 == r_count_21_io_out ? io_r_231_b : _GEN_6620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6622 = 9'he8 == r_count_21_io_out ? io_r_232_b : _GEN_6621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6623 = 9'he9 == r_count_21_io_out ? io_r_233_b : _GEN_6622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6624 = 9'hea == r_count_21_io_out ? io_r_234_b : _GEN_6623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6625 = 9'heb == r_count_21_io_out ? io_r_235_b : _GEN_6624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6626 = 9'hec == r_count_21_io_out ? io_r_236_b : _GEN_6625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6627 = 9'hed == r_count_21_io_out ? io_r_237_b : _GEN_6626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6628 = 9'hee == r_count_21_io_out ? io_r_238_b : _GEN_6627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6629 = 9'hef == r_count_21_io_out ? io_r_239_b : _GEN_6628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6630 = 9'hf0 == r_count_21_io_out ? io_r_240_b : _GEN_6629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6631 = 9'hf1 == r_count_21_io_out ? io_r_241_b : _GEN_6630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6632 = 9'hf2 == r_count_21_io_out ? io_r_242_b : _GEN_6631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6633 = 9'hf3 == r_count_21_io_out ? io_r_243_b : _GEN_6632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6634 = 9'hf4 == r_count_21_io_out ? io_r_244_b : _GEN_6633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6635 = 9'hf5 == r_count_21_io_out ? io_r_245_b : _GEN_6634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6636 = 9'hf6 == r_count_21_io_out ? io_r_246_b : _GEN_6635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6637 = 9'hf7 == r_count_21_io_out ? io_r_247_b : _GEN_6636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6638 = 9'hf8 == r_count_21_io_out ? io_r_248_b : _GEN_6637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6639 = 9'hf9 == r_count_21_io_out ? io_r_249_b : _GEN_6638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6640 = 9'hfa == r_count_21_io_out ? io_r_250_b : _GEN_6639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6641 = 9'hfb == r_count_21_io_out ? io_r_251_b : _GEN_6640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6642 = 9'hfc == r_count_21_io_out ? io_r_252_b : _GEN_6641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6643 = 9'hfd == r_count_21_io_out ? io_r_253_b : _GEN_6642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6644 = 9'hfe == r_count_21_io_out ? io_r_254_b : _GEN_6643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6645 = 9'hff == r_count_21_io_out ? io_r_255_b : _GEN_6644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6646 = 9'h100 == r_count_21_io_out ? io_r_256_b : _GEN_6645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6647 = 9'h101 == r_count_21_io_out ? io_r_257_b : _GEN_6646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6648 = 9'h102 == r_count_21_io_out ? io_r_258_b : _GEN_6647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6649 = 9'h103 == r_count_21_io_out ? io_r_259_b : _GEN_6648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6650 = 9'h104 == r_count_21_io_out ? io_r_260_b : _GEN_6649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6651 = 9'h105 == r_count_21_io_out ? io_r_261_b : _GEN_6650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6652 = 9'h106 == r_count_21_io_out ? io_r_262_b : _GEN_6651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6653 = 9'h107 == r_count_21_io_out ? io_r_263_b : _GEN_6652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6654 = 9'h108 == r_count_21_io_out ? io_r_264_b : _GEN_6653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6655 = 9'h109 == r_count_21_io_out ? io_r_265_b : _GEN_6654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6656 = 9'h10a == r_count_21_io_out ? io_r_266_b : _GEN_6655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6657 = 9'h10b == r_count_21_io_out ? io_r_267_b : _GEN_6656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6658 = 9'h10c == r_count_21_io_out ? io_r_268_b : _GEN_6657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6659 = 9'h10d == r_count_21_io_out ? io_r_269_b : _GEN_6658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6660 = 9'h10e == r_count_21_io_out ? io_r_270_b : _GEN_6659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6661 = 9'h10f == r_count_21_io_out ? io_r_271_b : _GEN_6660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6662 = 9'h110 == r_count_21_io_out ? io_r_272_b : _GEN_6661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6663 = 9'h111 == r_count_21_io_out ? io_r_273_b : _GEN_6662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6664 = 9'h112 == r_count_21_io_out ? io_r_274_b : _GEN_6663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6665 = 9'h113 == r_count_21_io_out ? io_r_275_b : _GEN_6664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6666 = 9'h114 == r_count_21_io_out ? io_r_276_b : _GEN_6665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6667 = 9'h115 == r_count_21_io_out ? io_r_277_b : _GEN_6666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6668 = 9'h116 == r_count_21_io_out ? io_r_278_b : _GEN_6667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6669 = 9'h117 == r_count_21_io_out ? io_r_279_b : _GEN_6668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6670 = 9'h118 == r_count_21_io_out ? io_r_280_b : _GEN_6669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6671 = 9'h119 == r_count_21_io_out ? io_r_281_b : _GEN_6670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6672 = 9'h11a == r_count_21_io_out ? io_r_282_b : _GEN_6671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6673 = 9'h11b == r_count_21_io_out ? io_r_283_b : _GEN_6672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6674 = 9'h11c == r_count_21_io_out ? io_r_284_b : _GEN_6673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6675 = 9'h11d == r_count_21_io_out ? io_r_285_b : _GEN_6674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6676 = 9'h11e == r_count_21_io_out ? io_r_286_b : _GEN_6675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6677 = 9'h11f == r_count_21_io_out ? io_r_287_b : _GEN_6676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6678 = 9'h120 == r_count_21_io_out ? io_r_288_b : _GEN_6677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6679 = 9'h121 == r_count_21_io_out ? io_r_289_b : _GEN_6678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6680 = 9'h122 == r_count_21_io_out ? io_r_290_b : _GEN_6679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6681 = 9'h123 == r_count_21_io_out ? io_r_291_b : _GEN_6680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6682 = 9'h124 == r_count_21_io_out ? io_r_292_b : _GEN_6681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6683 = 9'h125 == r_count_21_io_out ? io_r_293_b : _GEN_6682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6684 = 9'h126 == r_count_21_io_out ? io_r_294_b : _GEN_6683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6685 = 9'h127 == r_count_21_io_out ? io_r_295_b : _GEN_6684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6686 = 9'h128 == r_count_21_io_out ? io_r_296_b : _GEN_6685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6687 = 9'h129 == r_count_21_io_out ? io_r_297_b : _GEN_6686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6688 = 9'h12a == r_count_21_io_out ? io_r_298_b : _GEN_6687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6691 = 9'h1 == r_count_22_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6692 = 9'h2 == r_count_22_io_out ? io_r_2_b : _GEN_6691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6693 = 9'h3 == r_count_22_io_out ? io_r_3_b : _GEN_6692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6694 = 9'h4 == r_count_22_io_out ? io_r_4_b : _GEN_6693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6695 = 9'h5 == r_count_22_io_out ? io_r_5_b : _GEN_6694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6696 = 9'h6 == r_count_22_io_out ? io_r_6_b : _GEN_6695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6697 = 9'h7 == r_count_22_io_out ? io_r_7_b : _GEN_6696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6698 = 9'h8 == r_count_22_io_out ? io_r_8_b : _GEN_6697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6699 = 9'h9 == r_count_22_io_out ? io_r_9_b : _GEN_6698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6700 = 9'ha == r_count_22_io_out ? io_r_10_b : _GEN_6699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6701 = 9'hb == r_count_22_io_out ? io_r_11_b : _GEN_6700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6702 = 9'hc == r_count_22_io_out ? io_r_12_b : _GEN_6701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6703 = 9'hd == r_count_22_io_out ? io_r_13_b : _GEN_6702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6704 = 9'he == r_count_22_io_out ? io_r_14_b : _GEN_6703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6705 = 9'hf == r_count_22_io_out ? io_r_15_b : _GEN_6704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6706 = 9'h10 == r_count_22_io_out ? io_r_16_b : _GEN_6705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6707 = 9'h11 == r_count_22_io_out ? io_r_17_b : _GEN_6706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6708 = 9'h12 == r_count_22_io_out ? io_r_18_b : _GEN_6707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6709 = 9'h13 == r_count_22_io_out ? io_r_19_b : _GEN_6708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6710 = 9'h14 == r_count_22_io_out ? io_r_20_b : _GEN_6709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6711 = 9'h15 == r_count_22_io_out ? io_r_21_b : _GEN_6710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6712 = 9'h16 == r_count_22_io_out ? io_r_22_b : _GEN_6711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6713 = 9'h17 == r_count_22_io_out ? io_r_23_b : _GEN_6712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6714 = 9'h18 == r_count_22_io_out ? io_r_24_b : _GEN_6713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6715 = 9'h19 == r_count_22_io_out ? io_r_25_b : _GEN_6714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6716 = 9'h1a == r_count_22_io_out ? io_r_26_b : _GEN_6715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6717 = 9'h1b == r_count_22_io_out ? io_r_27_b : _GEN_6716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6718 = 9'h1c == r_count_22_io_out ? io_r_28_b : _GEN_6717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6719 = 9'h1d == r_count_22_io_out ? io_r_29_b : _GEN_6718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6720 = 9'h1e == r_count_22_io_out ? io_r_30_b : _GEN_6719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6721 = 9'h1f == r_count_22_io_out ? io_r_31_b : _GEN_6720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6722 = 9'h20 == r_count_22_io_out ? io_r_32_b : _GEN_6721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6723 = 9'h21 == r_count_22_io_out ? io_r_33_b : _GEN_6722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6724 = 9'h22 == r_count_22_io_out ? io_r_34_b : _GEN_6723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6725 = 9'h23 == r_count_22_io_out ? io_r_35_b : _GEN_6724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6726 = 9'h24 == r_count_22_io_out ? io_r_36_b : _GEN_6725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6727 = 9'h25 == r_count_22_io_out ? io_r_37_b : _GEN_6726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6728 = 9'h26 == r_count_22_io_out ? io_r_38_b : _GEN_6727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6729 = 9'h27 == r_count_22_io_out ? io_r_39_b : _GEN_6728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6730 = 9'h28 == r_count_22_io_out ? io_r_40_b : _GEN_6729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6731 = 9'h29 == r_count_22_io_out ? io_r_41_b : _GEN_6730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6732 = 9'h2a == r_count_22_io_out ? io_r_42_b : _GEN_6731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6733 = 9'h2b == r_count_22_io_out ? io_r_43_b : _GEN_6732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6734 = 9'h2c == r_count_22_io_out ? io_r_44_b : _GEN_6733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6735 = 9'h2d == r_count_22_io_out ? io_r_45_b : _GEN_6734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6736 = 9'h2e == r_count_22_io_out ? io_r_46_b : _GEN_6735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6737 = 9'h2f == r_count_22_io_out ? io_r_47_b : _GEN_6736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6738 = 9'h30 == r_count_22_io_out ? io_r_48_b : _GEN_6737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6739 = 9'h31 == r_count_22_io_out ? io_r_49_b : _GEN_6738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6740 = 9'h32 == r_count_22_io_out ? io_r_50_b : _GEN_6739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6741 = 9'h33 == r_count_22_io_out ? io_r_51_b : _GEN_6740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6742 = 9'h34 == r_count_22_io_out ? io_r_52_b : _GEN_6741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6743 = 9'h35 == r_count_22_io_out ? io_r_53_b : _GEN_6742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6744 = 9'h36 == r_count_22_io_out ? io_r_54_b : _GEN_6743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6745 = 9'h37 == r_count_22_io_out ? io_r_55_b : _GEN_6744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6746 = 9'h38 == r_count_22_io_out ? io_r_56_b : _GEN_6745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6747 = 9'h39 == r_count_22_io_out ? io_r_57_b : _GEN_6746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6748 = 9'h3a == r_count_22_io_out ? io_r_58_b : _GEN_6747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6749 = 9'h3b == r_count_22_io_out ? io_r_59_b : _GEN_6748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6750 = 9'h3c == r_count_22_io_out ? io_r_60_b : _GEN_6749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6751 = 9'h3d == r_count_22_io_out ? io_r_61_b : _GEN_6750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6752 = 9'h3e == r_count_22_io_out ? io_r_62_b : _GEN_6751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6753 = 9'h3f == r_count_22_io_out ? io_r_63_b : _GEN_6752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6754 = 9'h40 == r_count_22_io_out ? io_r_64_b : _GEN_6753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6755 = 9'h41 == r_count_22_io_out ? io_r_65_b : _GEN_6754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6756 = 9'h42 == r_count_22_io_out ? io_r_66_b : _GEN_6755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6757 = 9'h43 == r_count_22_io_out ? io_r_67_b : _GEN_6756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6758 = 9'h44 == r_count_22_io_out ? io_r_68_b : _GEN_6757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6759 = 9'h45 == r_count_22_io_out ? io_r_69_b : _GEN_6758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6760 = 9'h46 == r_count_22_io_out ? io_r_70_b : _GEN_6759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6761 = 9'h47 == r_count_22_io_out ? io_r_71_b : _GEN_6760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6762 = 9'h48 == r_count_22_io_out ? io_r_72_b : _GEN_6761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6763 = 9'h49 == r_count_22_io_out ? io_r_73_b : _GEN_6762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6764 = 9'h4a == r_count_22_io_out ? io_r_74_b : _GEN_6763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6765 = 9'h4b == r_count_22_io_out ? io_r_75_b : _GEN_6764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6766 = 9'h4c == r_count_22_io_out ? io_r_76_b : _GEN_6765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6767 = 9'h4d == r_count_22_io_out ? io_r_77_b : _GEN_6766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6768 = 9'h4e == r_count_22_io_out ? io_r_78_b : _GEN_6767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6769 = 9'h4f == r_count_22_io_out ? io_r_79_b : _GEN_6768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6770 = 9'h50 == r_count_22_io_out ? io_r_80_b : _GEN_6769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6771 = 9'h51 == r_count_22_io_out ? io_r_81_b : _GEN_6770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6772 = 9'h52 == r_count_22_io_out ? io_r_82_b : _GEN_6771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6773 = 9'h53 == r_count_22_io_out ? io_r_83_b : _GEN_6772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6774 = 9'h54 == r_count_22_io_out ? io_r_84_b : _GEN_6773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6775 = 9'h55 == r_count_22_io_out ? io_r_85_b : _GEN_6774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6776 = 9'h56 == r_count_22_io_out ? io_r_86_b : _GEN_6775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6777 = 9'h57 == r_count_22_io_out ? io_r_87_b : _GEN_6776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6778 = 9'h58 == r_count_22_io_out ? io_r_88_b : _GEN_6777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6779 = 9'h59 == r_count_22_io_out ? io_r_89_b : _GEN_6778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6780 = 9'h5a == r_count_22_io_out ? io_r_90_b : _GEN_6779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6781 = 9'h5b == r_count_22_io_out ? io_r_91_b : _GEN_6780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6782 = 9'h5c == r_count_22_io_out ? io_r_92_b : _GEN_6781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6783 = 9'h5d == r_count_22_io_out ? io_r_93_b : _GEN_6782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6784 = 9'h5e == r_count_22_io_out ? io_r_94_b : _GEN_6783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6785 = 9'h5f == r_count_22_io_out ? io_r_95_b : _GEN_6784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6786 = 9'h60 == r_count_22_io_out ? io_r_96_b : _GEN_6785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6787 = 9'h61 == r_count_22_io_out ? io_r_97_b : _GEN_6786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6788 = 9'h62 == r_count_22_io_out ? io_r_98_b : _GEN_6787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6789 = 9'h63 == r_count_22_io_out ? io_r_99_b : _GEN_6788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6790 = 9'h64 == r_count_22_io_out ? io_r_100_b : _GEN_6789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6791 = 9'h65 == r_count_22_io_out ? io_r_101_b : _GEN_6790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6792 = 9'h66 == r_count_22_io_out ? io_r_102_b : _GEN_6791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6793 = 9'h67 == r_count_22_io_out ? io_r_103_b : _GEN_6792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6794 = 9'h68 == r_count_22_io_out ? io_r_104_b : _GEN_6793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6795 = 9'h69 == r_count_22_io_out ? io_r_105_b : _GEN_6794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6796 = 9'h6a == r_count_22_io_out ? io_r_106_b : _GEN_6795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6797 = 9'h6b == r_count_22_io_out ? io_r_107_b : _GEN_6796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6798 = 9'h6c == r_count_22_io_out ? io_r_108_b : _GEN_6797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6799 = 9'h6d == r_count_22_io_out ? io_r_109_b : _GEN_6798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6800 = 9'h6e == r_count_22_io_out ? io_r_110_b : _GEN_6799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6801 = 9'h6f == r_count_22_io_out ? io_r_111_b : _GEN_6800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6802 = 9'h70 == r_count_22_io_out ? io_r_112_b : _GEN_6801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6803 = 9'h71 == r_count_22_io_out ? io_r_113_b : _GEN_6802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6804 = 9'h72 == r_count_22_io_out ? io_r_114_b : _GEN_6803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6805 = 9'h73 == r_count_22_io_out ? io_r_115_b : _GEN_6804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6806 = 9'h74 == r_count_22_io_out ? io_r_116_b : _GEN_6805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6807 = 9'h75 == r_count_22_io_out ? io_r_117_b : _GEN_6806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6808 = 9'h76 == r_count_22_io_out ? io_r_118_b : _GEN_6807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6809 = 9'h77 == r_count_22_io_out ? io_r_119_b : _GEN_6808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6810 = 9'h78 == r_count_22_io_out ? io_r_120_b : _GEN_6809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6811 = 9'h79 == r_count_22_io_out ? io_r_121_b : _GEN_6810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6812 = 9'h7a == r_count_22_io_out ? io_r_122_b : _GEN_6811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6813 = 9'h7b == r_count_22_io_out ? io_r_123_b : _GEN_6812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6814 = 9'h7c == r_count_22_io_out ? io_r_124_b : _GEN_6813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6815 = 9'h7d == r_count_22_io_out ? io_r_125_b : _GEN_6814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6816 = 9'h7e == r_count_22_io_out ? io_r_126_b : _GEN_6815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6817 = 9'h7f == r_count_22_io_out ? io_r_127_b : _GEN_6816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6818 = 9'h80 == r_count_22_io_out ? io_r_128_b : _GEN_6817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6819 = 9'h81 == r_count_22_io_out ? io_r_129_b : _GEN_6818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6820 = 9'h82 == r_count_22_io_out ? io_r_130_b : _GEN_6819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6821 = 9'h83 == r_count_22_io_out ? io_r_131_b : _GEN_6820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6822 = 9'h84 == r_count_22_io_out ? io_r_132_b : _GEN_6821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6823 = 9'h85 == r_count_22_io_out ? io_r_133_b : _GEN_6822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6824 = 9'h86 == r_count_22_io_out ? io_r_134_b : _GEN_6823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6825 = 9'h87 == r_count_22_io_out ? io_r_135_b : _GEN_6824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6826 = 9'h88 == r_count_22_io_out ? io_r_136_b : _GEN_6825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6827 = 9'h89 == r_count_22_io_out ? io_r_137_b : _GEN_6826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6828 = 9'h8a == r_count_22_io_out ? io_r_138_b : _GEN_6827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6829 = 9'h8b == r_count_22_io_out ? io_r_139_b : _GEN_6828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6830 = 9'h8c == r_count_22_io_out ? io_r_140_b : _GEN_6829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6831 = 9'h8d == r_count_22_io_out ? io_r_141_b : _GEN_6830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6832 = 9'h8e == r_count_22_io_out ? io_r_142_b : _GEN_6831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6833 = 9'h8f == r_count_22_io_out ? io_r_143_b : _GEN_6832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6834 = 9'h90 == r_count_22_io_out ? io_r_144_b : _GEN_6833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6835 = 9'h91 == r_count_22_io_out ? io_r_145_b : _GEN_6834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6836 = 9'h92 == r_count_22_io_out ? io_r_146_b : _GEN_6835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6837 = 9'h93 == r_count_22_io_out ? io_r_147_b : _GEN_6836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6838 = 9'h94 == r_count_22_io_out ? io_r_148_b : _GEN_6837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6839 = 9'h95 == r_count_22_io_out ? io_r_149_b : _GEN_6838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6840 = 9'h96 == r_count_22_io_out ? io_r_150_b : _GEN_6839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6841 = 9'h97 == r_count_22_io_out ? io_r_151_b : _GEN_6840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6842 = 9'h98 == r_count_22_io_out ? io_r_152_b : _GEN_6841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6843 = 9'h99 == r_count_22_io_out ? io_r_153_b : _GEN_6842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6844 = 9'h9a == r_count_22_io_out ? io_r_154_b : _GEN_6843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6845 = 9'h9b == r_count_22_io_out ? io_r_155_b : _GEN_6844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6846 = 9'h9c == r_count_22_io_out ? io_r_156_b : _GEN_6845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6847 = 9'h9d == r_count_22_io_out ? io_r_157_b : _GEN_6846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6848 = 9'h9e == r_count_22_io_out ? io_r_158_b : _GEN_6847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6849 = 9'h9f == r_count_22_io_out ? io_r_159_b : _GEN_6848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6850 = 9'ha0 == r_count_22_io_out ? io_r_160_b : _GEN_6849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6851 = 9'ha1 == r_count_22_io_out ? io_r_161_b : _GEN_6850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6852 = 9'ha2 == r_count_22_io_out ? io_r_162_b : _GEN_6851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6853 = 9'ha3 == r_count_22_io_out ? io_r_163_b : _GEN_6852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6854 = 9'ha4 == r_count_22_io_out ? io_r_164_b : _GEN_6853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6855 = 9'ha5 == r_count_22_io_out ? io_r_165_b : _GEN_6854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6856 = 9'ha6 == r_count_22_io_out ? io_r_166_b : _GEN_6855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6857 = 9'ha7 == r_count_22_io_out ? io_r_167_b : _GEN_6856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6858 = 9'ha8 == r_count_22_io_out ? io_r_168_b : _GEN_6857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6859 = 9'ha9 == r_count_22_io_out ? io_r_169_b : _GEN_6858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6860 = 9'haa == r_count_22_io_out ? io_r_170_b : _GEN_6859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6861 = 9'hab == r_count_22_io_out ? io_r_171_b : _GEN_6860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6862 = 9'hac == r_count_22_io_out ? io_r_172_b : _GEN_6861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6863 = 9'had == r_count_22_io_out ? io_r_173_b : _GEN_6862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6864 = 9'hae == r_count_22_io_out ? io_r_174_b : _GEN_6863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6865 = 9'haf == r_count_22_io_out ? io_r_175_b : _GEN_6864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6866 = 9'hb0 == r_count_22_io_out ? io_r_176_b : _GEN_6865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6867 = 9'hb1 == r_count_22_io_out ? io_r_177_b : _GEN_6866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6868 = 9'hb2 == r_count_22_io_out ? io_r_178_b : _GEN_6867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6869 = 9'hb3 == r_count_22_io_out ? io_r_179_b : _GEN_6868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6870 = 9'hb4 == r_count_22_io_out ? io_r_180_b : _GEN_6869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6871 = 9'hb5 == r_count_22_io_out ? io_r_181_b : _GEN_6870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6872 = 9'hb6 == r_count_22_io_out ? io_r_182_b : _GEN_6871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6873 = 9'hb7 == r_count_22_io_out ? io_r_183_b : _GEN_6872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6874 = 9'hb8 == r_count_22_io_out ? io_r_184_b : _GEN_6873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6875 = 9'hb9 == r_count_22_io_out ? io_r_185_b : _GEN_6874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6876 = 9'hba == r_count_22_io_out ? io_r_186_b : _GEN_6875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6877 = 9'hbb == r_count_22_io_out ? io_r_187_b : _GEN_6876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6878 = 9'hbc == r_count_22_io_out ? io_r_188_b : _GEN_6877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6879 = 9'hbd == r_count_22_io_out ? io_r_189_b : _GEN_6878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6880 = 9'hbe == r_count_22_io_out ? io_r_190_b : _GEN_6879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6881 = 9'hbf == r_count_22_io_out ? io_r_191_b : _GEN_6880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6882 = 9'hc0 == r_count_22_io_out ? io_r_192_b : _GEN_6881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6883 = 9'hc1 == r_count_22_io_out ? io_r_193_b : _GEN_6882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6884 = 9'hc2 == r_count_22_io_out ? io_r_194_b : _GEN_6883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6885 = 9'hc3 == r_count_22_io_out ? io_r_195_b : _GEN_6884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6886 = 9'hc4 == r_count_22_io_out ? io_r_196_b : _GEN_6885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6887 = 9'hc5 == r_count_22_io_out ? io_r_197_b : _GEN_6886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6888 = 9'hc6 == r_count_22_io_out ? io_r_198_b : _GEN_6887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6889 = 9'hc7 == r_count_22_io_out ? io_r_199_b : _GEN_6888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6890 = 9'hc8 == r_count_22_io_out ? io_r_200_b : _GEN_6889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6891 = 9'hc9 == r_count_22_io_out ? io_r_201_b : _GEN_6890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6892 = 9'hca == r_count_22_io_out ? io_r_202_b : _GEN_6891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6893 = 9'hcb == r_count_22_io_out ? io_r_203_b : _GEN_6892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6894 = 9'hcc == r_count_22_io_out ? io_r_204_b : _GEN_6893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6895 = 9'hcd == r_count_22_io_out ? io_r_205_b : _GEN_6894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6896 = 9'hce == r_count_22_io_out ? io_r_206_b : _GEN_6895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6897 = 9'hcf == r_count_22_io_out ? io_r_207_b : _GEN_6896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6898 = 9'hd0 == r_count_22_io_out ? io_r_208_b : _GEN_6897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6899 = 9'hd1 == r_count_22_io_out ? io_r_209_b : _GEN_6898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6900 = 9'hd2 == r_count_22_io_out ? io_r_210_b : _GEN_6899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6901 = 9'hd3 == r_count_22_io_out ? io_r_211_b : _GEN_6900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6902 = 9'hd4 == r_count_22_io_out ? io_r_212_b : _GEN_6901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6903 = 9'hd5 == r_count_22_io_out ? io_r_213_b : _GEN_6902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6904 = 9'hd6 == r_count_22_io_out ? io_r_214_b : _GEN_6903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6905 = 9'hd7 == r_count_22_io_out ? io_r_215_b : _GEN_6904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6906 = 9'hd8 == r_count_22_io_out ? io_r_216_b : _GEN_6905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6907 = 9'hd9 == r_count_22_io_out ? io_r_217_b : _GEN_6906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6908 = 9'hda == r_count_22_io_out ? io_r_218_b : _GEN_6907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6909 = 9'hdb == r_count_22_io_out ? io_r_219_b : _GEN_6908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6910 = 9'hdc == r_count_22_io_out ? io_r_220_b : _GEN_6909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6911 = 9'hdd == r_count_22_io_out ? io_r_221_b : _GEN_6910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6912 = 9'hde == r_count_22_io_out ? io_r_222_b : _GEN_6911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6913 = 9'hdf == r_count_22_io_out ? io_r_223_b : _GEN_6912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6914 = 9'he0 == r_count_22_io_out ? io_r_224_b : _GEN_6913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6915 = 9'he1 == r_count_22_io_out ? io_r_225_b : _GEN_6914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6916 = 9'he2 == r_count_22_io_out ? io_r_226_b : _GEN_6915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6917 = 9'he3 == r_count_22_io_out ? io_r_227_b : _GEN_6916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6918 = 9'he4 == r_count_22_io_out ? io_r_228_b : _GEN_6917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6919 = 9'he5 == r_count_22_io_out ? io_r_229_b : _GEN_6918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6920 = 9'he6 == r_count_22_io_out ? io_r_230_b : _GEN_6919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6921 = 9'he7 == r_count_22_io_out ? io_r_231_b : _GEN_6920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6922 = 9'he8 == r_count_22_io_out ? io_r_232_b : _GEN_6921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6923 = 9'he9 == r_count_22_io_out ? io_r_233_b : _GEN_6922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6924 = 9'hea == r_count_22_io_out ? io_r_234_b : _GEN_6923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6925 = 9'heb == r_count_22_io_out ? io_r_235_b : _GEN_6924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6926 = 9'hec == r_count_22_io_out ? io_r_236_b : _GEN_6925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6927 = 9'hed == r_count_22_io_out ? io_r_237_b : _GEN_6926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6928 = 9'hee == r_count_22_io_out ? io_r_238_b : _GEN_6927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6929 = 9'hef == r_count_22_io_out ? io_r_239_b : _GEN_6928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6930 = 9'hf0 == r_count_22_io_out ? io_r_240_b : _GEN_6929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6931 = 9'hf1 == r_count_22_io_out ? io_r_241_b : _GEN_6930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6932 = 9'hf2 == r_count_22_io_out ? io_r_242_b : _GEN_6931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6933 = 9'hf3 == r_count_22_io_out ? io_r_243_b : _GEN_6932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6934 = 9'hf4 == r_count_22_io_out ? io_r_244_b : _GEN_6933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6935 = 9'hf5 == r_count_22_io_out ? io_r_245_b : _GEN_6934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6936 = 9'hf6 == r_count_22_io_out ? io_r_246_b : _GEN_6935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6937 = 9'hf7 == r_count_22_io_out ? io_r_247_b : _GEN_6936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6938 = 9'hf8 == r_count_22_io_out ? io_r_248_b : _GEN_6937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6939 = 9'hf9 == r_count_22_io_out ? io_r_249_b : _GEN_6938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6940 = 9'hfa == r_count_22_io_out ? io_r_250_b : _GEN_6939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6941 = 9'hfb == r_count_22_io_out ? io_r_251_b : _GEN_6940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6942 = 9'hfc == r_count_22_io_out ? io_r_252_b : _GEN_6941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6943 = 9'hfd == r_count_22_io_out ? io_r_253_b : _GEN_6942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6944 = 9'hfe == r_count_22_io_out ? io_r_254_b : _GEN_6943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6945 = 9'hff == r_count_22_io_out ? io_r_255_b : _GEN_6944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6946 = 9'h100 == r_count_22_io_out ? io_r_256_b : _GEN_6945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6947 = 9'h101 == r_count_22_io_out ? io_r_257_b : _GEN_6946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6948 = 9'h102 == r_count_22_io_out ? io_r_258_b : _GEN_6947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6949 = 9'h103 == r_count_22_io_out ? io_r_259_b : _GEN_6948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6950 = 9'h104 == r_count_22_io_out ? io_r_260_b : _GEN_6949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6951 = 9'h105 == r_count_22_io_out ? io_r_261_b : _GEN_6950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6952 = 9'h106 == r_count_22_io_out ? io_r_262_b : _GEN_6951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6953 = 9'h107 == r_count_22_io_out ? io_r_263_b : _GEN_6952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6954 = 9'h108 == r_count_22_io_out ? io_r_264_b : _GEN_6953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6955 = 9'h109 == r_count_22_io_out ? io_r_265_b : _GEN_6954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6956 = 9'h10a == r_count_22_io_out ? io_r_266_b : _GEN_6955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6957 = 9'h10b == r_count_22_io_out ? io_r_267_b : _GEN_6956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6958 = 9'h10c == r_count_22_io_out ? io_r_268_b : _GEN_6957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6959 = 9'h10d == r_count_22_io_out ? io_r_269_b : _GEN_6958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6960 = 9'h10e == r_count_22_io_out ? io_r_270_b : _GEN_6959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6961 = 9'h10f == r_count_22_io_out ? io_r_271_b : _GEN_6960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6962 = 9'h110 == r_count_22_io_out ? io_r_272_b : _GEN_6961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6963 = 9'h111 == r_count_22_io_out ? io_r_273_b : _GEN_6962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6964 = 9'h112 == r_count_22_io_out ? io_r_274_b : _GEN_6963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6965 = 9'h113 == r_count_22_io_out ? io_r_275_b : _GEN_6964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6966 = 9'h114 == r_count_22_io_out ? io_r_276_b : _GEN_6965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6967 = 9'h115 == r_count_22_io_out ? io_r_277_b : _GEN_6966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6968 = 9'h116 == r_count_22_io_out ? io_r_278_b : _GEN_6967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6969 = 9'h117 == r_count_22_io_out ? io_r_279_b : _GEN_6968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6970 = 9'h118 == r_count_22_io_out ? io_r_280_b : _GEN_6969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6971 = 9'h119 == r_count_22_io_out ? io_r_281_b : _GEN_6970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6972 = 9'h11a == r_count_22_io_out ? io_r_282_b : _GEN_6971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6973 = 9'h11b == r_count_22_io_out ? io_r_283_b : _GEN_6972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6974 = 9'h11c == r_count_22_io_out ? io_r_284_b : _GEN_6973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6975 = 9'h11d == r_count_22_io_out ? io_r_285_b : _GEN_6974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6976 = 9'h11e == r_count_22_io_out ? io_r_286_b : _GEN_6975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6977 = 9'h11f == r_count_22_io_out ? io_r_287_b : _GEN_6976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6978 = 9'h120 == r_count_22_io_out ? io_r_288_b : _GEN_6977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6979 = 9'h121 == r_count_22_io_out ? io_r_289_b : _GEN_6978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6980 = 9'h122 == r_count_22_io_out ? io_r_290_b : _GEN_6979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6981 = 9'h123 == r_count_22_io_out ? io_r_291_b : _GEN_6980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6982 = 9'h124 == r_count_22_io_out ? io_r_292_b : _GEN_6981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6983 = 9'h125 == r_count_22_io_out ? io_r_293_b : _GEN_6982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6984 = 9'h126 == r_count_22_io_out ? io_r_294_b : _GEN_6983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6985 = 9'h127 == r_count_22_io_out ? io_r_295_b : _GEN_6984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6986 = 9'h128 == r_count_22_io_out ? io_r_296_b : _GEN_6985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6987 = 9'h129 == r_count_22_io_out ? io_r_297_b : _GEN_6986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6988 = 9'h12a == r_count_22_io_out ? io_r_298_b : _GEN_6987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6991 = 9'h1 == r_count_23_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6992 = 9'h2 == r_count_23_io_out ? io_r_2_b : _GEN_6991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6993 = 9'h3 == r_count_23_io_out ? io_r_3_b : _GEN_6992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6994 = 9'h4 == r_count_23_io_out ? io_r_4_b : _GEN_6993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6995 = 9'h5 == r_count_23_io_out ? io_r_5_b : _GEN_6994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6996 = 9'h6 == r_count_23_io_out ? io_r_6_b : _GEN_6995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6997 = 9'h7 == r_count_23_io_out ? io_r_7_b : _GEN_6996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6998 = 9'h8 == r_count_23_io_out ? io_r_8_b : _GEN_6997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6999 = 9'h9 == r_count_23_io_out ? io_r_9_b : _GEN_6998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7000 = 9'ha == r_count_23_io_out ? io_r_10_b : _GEN_6999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7001 = 9'hb == r_count_23_io_out ? io_r_11_b : _GEN_7000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7002 = 9'hc == r_count_23_io_out ? io_r_12_b : _GEN_7001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7003 = 9'hd == r_count_23_io_out ? io_r_13_b : _GEN_7002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7004 = 9'he == r_count_23_io_out ? io_r_14_b : _GEN_7003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7005 = 9'hf == r_count_23_io_out ? io_r_15_b : _GEN_7004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7006 = 9'h10 == r_count_23_io_out ? io_r_16_b : _GEN_7005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7007 = 9'h11 == r_count_23_io_out ? io_r_17_b : _GEN_7006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7008 = 9'h12 == r_count_23_io_out ? io_r_18_b : _GEN_7007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7009 = 9'h13 == r_count_23_io_out ? io_r_19_b : _GEN_7008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7010 = 9'h14 == r_count_23_io_out ? io_r_20_b : _GEN_7009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7011 = 9'h15 == r_count_23_io_out ? io_r_21_b : _GEN_7010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7012 = 9'h16 == r_count_23_io_out ? io_r_22_b : _GEN_7011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7013 = 9'h17 == r_count_23_io_out ? io_r_23_b : _GEN_7012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7014 = 9'h18 == r_count_23_io_out ? io_r_24_b : _GEN_7013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7015 = 9'h19 == r_count_23_io_out ? io_r_25_b : _GEN_7014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7016 = 9'h1a == r_count_23_io_out ? io_r_26_b : _GEN_7015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7017 = 9'h1b == r_count_23_io_out ? io_r_27_b : _GEN_7016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7018 = 9'h1c == r_count_23_io_out ? io_r_28_b : _GEN_7017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7019 = 9'h1d == r_count_23_io_out ? io_r_29_b : _GEN_7018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7020 = 9'h1e == r_count_23_io_out ? io_r_30_b : _GEN_7019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7021 = 9'h1f == r_count_23_io_out ? io_r_31_b : _GEN_7020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7022 = 9'h20 == r_count_23_io_out ? io_r_32_b : _GEN_7021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7023 = 9'h21 == r_count_23_io_out ? io_r_33_b : _GEN_7022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7024 = 9'h22 == r_count_23_io_out ? io_r_34_b : _GEN_7023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7025 = 9'h23 == r_count_23_io_out ? io_r_35_b : _GEN_7024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7026 = 9'h24 == r_count_23_io_out ? io_r_36_b : _GEN_7025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7027 = 9'h25 == r_count_23_io_out ? io_r_37_b : _GEN_7026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7028 = 9'h26 == r_count_23_io_out ? io_r_38_b : _GEN_7027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7029 = 9'h27 == r_count_23_io_out ? io_r_39_b : _GEN_7028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7030 = 9'h28 == r_count_23_io_out ? io_r_40_b : _GEN_7029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7031 = 9'h29 == r_count_23_io_out ? io_r_41_b : _GEN_7030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7032 = 9'h2a == r_count_23_io_out ? io_r_42_b : _GEN_7031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7033 = 9'h2b == r_count_23_io_out ? io_r_43_b : _GEN_7032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7034 = 9'h2c == r_count_23_io_out ? io_r_44_b : _GEN_7033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7035 = 9'h2d == r_count_23_io_out ? io_r_45_b : _GEN_7034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7036 = 9'h2e == r_count_23_io_out ? io_r_46_b : _GEN_7035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7037 = 9'h2f == r_count_23_io_out ? io_r_47_b : _GEN_7036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7038 = 9'h30 == r_count_23_io_out ? io_r_48_b : _GEN_7037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7039 = 9'h31 == r_count_23_io_out ? io_r_49_b : _GEN_7038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7040 = 9'h32 == r_count_23_io_out ? io_r_50_b : _GEN_7039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7041 = 9'h33 == r_count_23_io_out ? io_r_51_b : _GEN_7040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7042 = 9'h34 == r_count_23_io_out ? io_r_52_b : _GEN_7041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7043 = 9'h35 == r_count_23_io_out ? io_r_53_b : _GEN_7042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7044 = 9'h36 == r_count_23_io_out ? io_r_54_b : _GEN_7043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7045 = 9'h37 == r_count_23_io_out ? io_r_55_b : _GEN_7044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7046 = 9'h38 == r_count_23_io_out ? io_r_56_b : _GEN_7045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7047 = 9'h39 == r_count_23_io_out ? io_r_57_b : _GEN_7046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7048 = 9'h3a == r_count_23_io_out ? io_r_58_b : _GEN_7047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7049 = 9'h3b == r_count_23_io_out ? io_r_59_b : _GEN_7048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7050 = 9'h3c == r_count_23_io_out ? io_r_60_b : _GEN_7049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7051 = 9'h3d == r_count_23_io_out ? io_r_61_b : _GEN_7050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7052 = 9'h3e == r_count_23_io_out ? io_r_62_b : _GEN_7051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7053 = 9'h3f == r_count_23_io_out ? io_r_63_b : _GEN_7052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7054 = 9'h40 == r_count_23_io_out ? io_r_64_b : _GEN_7053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7055 = 9'h41 == r_count_23_io_out ? io_r_65_b : _GEN_7054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7056 = 9'h42 == r_count_23_io_out ? io_r_66_b : _GEN_7055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7057 = 9'h43 == r_count_23_io_out ? io_r_67_b : _GEN_7056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7058 = 9'h44 == r_count_23_io_out ? io_r_68_b : _GEN_7057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7059 = 9'h45 == r_count_23_io_out ? io_r_69_b : _GEN_7058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7060 = 9'h46 == r_count_23_io_out ? io_r_70_b : _GEN_7059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7061 = 9'h47 == r_count_23_io_out ? io_r_71_b : _GEN_7060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7062 = 9'h48 == r_count_23_io_out ? io_r_72_b : _GEN_7061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7063 = 9'h49 == r_count_23_io_out ? io_r_73_b : _GEN_7062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7064 = 9'h4a == r_count_23_io_out ? io_r_74_b : _GEN_7063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7065 = 9'h4b == r_count_23_io_out ? io_r_75_b : _GEN_7064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7066 = 9'h4c == r_count_23_io_out ? io_r_76_b : _GEN_7065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7067 = 9'h4d == r_count_23_io_out ? io_r_77_b : _GEN_7066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7068 = 9'h4e == r_count_23_io_out ? io_r_78_b : _GEN_7067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7069 = 9'h4f == r_count_23_io_out ? io_r_79_b : _GEN_7068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7070 = 9'h50 == r_count_23_io_out ? io_r_80_b : _GEN_7069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7071 = 9'h51 == r_count_23_io_out ? io_r_81_b : _GEN_7070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7072 = 9'h52 == r_count_23_io_out ? io_r_82_b : _GEN_7071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7073 = 9'h53 == r_count_23_io_out ? io_r_83_b : _GEN_7072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7074 = 9'h54 == r_count_23_io_out ? io_r_84_b : _GEN_7073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7075 = 9'h55 == r_count_23_io_out ? io_r_85_b : _GEN_7074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7076 = 9'h56 == r_count_23_io_out ? io_r_86_b : _GEN_7075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7077 = 9'h57 == r_count_23_io_out ? io_r_87_b : _GEN_7076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7078 = 9'h58 == r_count_23_io_out ? io_r_88_b : _GEN_7077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7079 = 9'h59 == r_count_23_io_out ? io_r_89_b : _GEN_7078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7080 = 9'h5a == r_count_23_io_out ? io_r_90_b : _GEN_7079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7081 = 9'h5b == r_count_23_io_out ? io_r_91_b : _GEN_7080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7082 = 9'h5c == r_count_23_io_out ? io_r_92_b : _GEN_7081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7083 = 9'h5d == r_count_23_io_out ? io_r_93_b : _GEN_7082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7084 = 9'h5e == r_count_23_io_out ? io_r_94_b : _GEN_7083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7085 = 9'h5f == r_count_23_io_out ? io_r_95_b : _GEN_7084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7086 = 9'h60 == r_count_23_io_out ? io_r_96_b : _GEN_7085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7087 = 9'h61 == r_count_23_io_out ? io_r_97_b : _GEN_7086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7088 = 9'h62 == r_count_23_io_out ? io_r_98_b : _GEN_7087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7089 = 9'h63 == r_count_23_io_out ? io_r_99_b : _GEN_7088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7090 = 9'h64 == r_count_23_io_out ? io_r_100_b : _GEN_7089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7091 = 9'h65 == r_count_23_io_out ? io_r_101_b : _GEN_7090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7092 = 9'h66 == r_count_23_io_out ? io_r_102_b : _GEN_7091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7093 = 9'h67 == r_count_23_io_out ? io_r_103_b : _GEN_7092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7094 = 9'h68 == r_count_23_io_out ? io_r_104_b : _GEN_7093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7095 = 9'h69 == r_count_23_io_out ? io_r_105_b : _GEN_7094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7096 = 9'h6a == r_count_23_io_out ? io_r_106_b : _GEN_7095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7097 = 9'h6b == r_count_23_io_out ? io_r_107_b : _GEN_7096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7098 = 9'h6c == r_count_23_io_out ? io_r_108_b : _GEN_7097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7099 = 9'h6d == r_count_23_io_out ? io_r_109_b : _GEN_7098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7100 = 9'h6e == r_count_23_io_out ? io_r_110_b : _GEN_7099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7101 = 9'h6f == r_count_23_io_out ? io_r_111_b : _GEN_7100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7102 = 9'h70 == r_count_23_io_out ? io_r_112_b : _GEN_7101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7103 = 9'h71 == r_count_23_io_out ? io_r_113_b : _GEN_7102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7104 = 9'h72 == r_count_23_io_out ? io_r_114_b : _GEN_7103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7105 = 9'h73 == r_count_23_io_out ? io_r_115_b : _GEN_7104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7106 = 9'h74 == r_count_23_io_out ? io_r_116_b : _GEN_7105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7107 = 9'h75 == r_count_23_io_out ? io_r_117_b : _GEN_7106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7108 = 9'h76 == r_count_23_io_out ? io_r_118_b : _GEN_7107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7109 = 9'h77 == r_count_23_io_out ? io_r_119_b : _GEN_7108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7110 = 9'h78 == r_count_23_io_out ? io_r_120_b : _GEN_7109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7111 = 9'h79 == r_count_23_io_out ? io_r_121_b : _GEN_7110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7112 = 9'h7a == r_count_23_io_out ? io_r_122_b : _GEN_7111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7113 = 9'h7b == r_count_23_io_out ? io_r_123_b : _GEN_7112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7114 = 9'h7c == r_count_23_io_out ? io_r_124_b : _GEN_7113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7115 = 9'h7d == r_count_23_io_out ? io_r_125_b : _GEN_7114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7116 = 9'h7e == r_count_23_io_out ? io_r_126_b : _GEN_7115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7117 = 9'h7f == r_count_23_io_out ? io_r_127_b : _GEN_7116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7118 = 9'h80 == r_count_23_io_out ? io_r_128_b : _GEN_7117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7119 = 9'h81 == r_count_23_io_out ? io_r_129_b : _GEN_7118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7120 = 9'h82 == r_count_23_io_out ? io_r_130_b : _GEN_7119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7121 = 9'h83 == r_count_23_io_out ? io_r_131_b : _GEN_7120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7122 = 9'h84 == r_count_23_io_out ? io_r_132_b : _GEN_7121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7123 = 9'h85 == r_count_23_io_out ? io_r_133_b : _GEN_7122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7124 = 9'h86 == r_count_23_io_out ? io_r_134_b : _GEN_7123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7125 = 9'h87 == r_count_23_io_out ? io_r_135_b : _GEN_7124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7126 = 9'h88 == r_count_23_io_out ? io_r_136_b : _GEN_7125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7127 = 9'h89 == r_count_23_io_out ? io_r_137_b : _GEN_7126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7128 = 9'h8a == r_count_23_io_out ? io_r_138_b : _GEN_7127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7129 = 9'h8b == r_count_23_io_out ? io_r_139_b : _GEN_7128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7130 = 9'h8c == r_count_23_io_out ? io_r_140_b : _GEN_7129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7131 = 9'h8d == r_count_23_io_out ? io_r_141_b : _GEN_7130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7132 = 9'h8e == r_count_23_io_out ? io_r_142_b : _GEN_7131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7133 = 9'h8f == r_count_23_io_out ? io_r_143_b : _GEN_7132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7134 = 9'h90 == r_count_23_io_out ? io_r_144_b : _GEN_7133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7135 = 9'h91 == r_count_23_io_out ? io_r_145_b : _GEN_7134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7136 = 9'h92 == r_count_23_io_out ? io_r_146_b : _GEN_7135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7137 = 9'h93 == r_count_23_io_out ? io_r_147_b : _GEN_7136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7138 = 9'h94 == r_count_23_io_out ? io_r_148_b : _GEN_7137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7139 = 9'h95 == r_count_23_io_out ? io_r_149_b : _GEN_7138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7140 = 9'h96 == r_count_23_io_out ? io_r_150_b : _GEN_7139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7141 = 9'h97 == r_count_23_io_out ? io_r_151_b : _GEN_7140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7142 = 9'h98 == r_count_23_io_out ? io_r_152_b : _GEN_7141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7143 = 9'h99 == r_count_23_io_out ? io_r_153_b : _GEN_7142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7144 = 9'h9a == r_count_23_io_out ? io_r_154_b : _GEN_7143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7145 = 9'h9b == r_count_23_io_out ? io_r_155_b : _GEN_7144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7146 = 9'h9c == r_count_23_io_out ? io_r_156_b : _GEN_7145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7147 = 9'h9d == r_count_23_io_out ? io_r_157_b : _GEN_7146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7148 = 9'h9e == r_count_23_io_out ? io_r_158_b : _GEN_7147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7149 = 9'h9f == r_count_23_io_out ? io_r_159_b : _GEN_7148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7150 = 9'ha0 == r_count_23_io_out ? io_r_160_b : _GEN_7149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7151 = 9'ha1 == r_count_23_io_out ? io_r_161_b : _GEN_7150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7152 = 9'ha2 == r_count_23_io_out ? io_r_162_b : _GEN_7151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7153 = 9'ha3 == r_count_23_io_out ? io_r_163_b : _GEN_7152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7154 = 9'ha4 == r_count_23_io_out ? io_r_164_b : _GEN_7153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7155 = 9'ha5 == r_count_23_io_out ? io_r_165_b : _GEN_7154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7156 = 9'ha6 == r_count_23_io_out ? io_r_166_b : _GEN_7155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7157 = 9'ha7 == r_count_23_io_out ? io_r_167_b : _GEN_7156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7158 = 9'ha8 == r_count_23_io_out ? io_r_168_b : _GEN_7157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7159 = 9'ha9 == r_count_23_io_out ? io_r_169_b : _GEN_7158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7160 = 9'haa == r_count_23_io_out ? io_r_170_b : _GEN_7159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7161 = 9'hab == r_count_23_io_out ? io_r_171_b : _GEN_7160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7162 = 9'hac == r_count_23_io_out ? io_r_172_b : _GEN_7161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7163 = 9'had == r_count_23_io_out ? io_r_173_b : _GEN_7162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7164 = 9'hae == r_count_23_io_out ? io_r_174_b : _GEN_7163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7165 = 9'haf == r_count_23_io_out ? io_r_175_b : _GEN_7164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7166 = 9'hb0 == r_count_23_io_out ? io_r_176_b : _GEN_7165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7167 = 9'hb1 == r_count_23_io_out ? io_r_177_b : _GEN_7166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7168 = 9'hb2 == r_count_23_io_out ? io_r_178_b : _GEN_7167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7169 = 9'hb3 == r_count_23_io_out ? io_r_179_b : _GEN_7168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7170 = 9'hb4 == r_count_23_io_out ? io_r_180_b : _GEN_7169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7171 = 9'hb5 == r_count_23_io_out ? io_r_181_b : _GEN_7170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7172 = 9'hb6 == r_count_23_io_out ? io_r_182_b : _GEN_7171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7173 = 9'hb7 == r_count_23_io_out ? io_r_183_b : _GEN_7172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7174 = 9'hb8 == r_count_23_io_out ? io_r_184_b : _GEN_7173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7175 = 9'hb9 == r_count_23_io_out ? io_r_185_b : _GEN_7174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7176 = 9'hba == r_count_23_io_out ? io_r_186_b : _GEN_7175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7177 = 9'hbb == r_count_23_io_out ? io_r_187_b : _GEN_7176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7178 = 9'hbc == r_count_23_io_out ? io_r_188_b : _GEN_7177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7179 = 9'hbd == r_count_23_io_out ? io_r_189_b : _GEN_7178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7180 = 9'hbe == r_count_23_io_out ? io_r_190_b : _GEN_7179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7181 = 9'hbf == r_count_23_io_out ? io_r_191_b : _GEN_7180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7182 = 9'hc0 == r_count_23_io_out ? io_r_192_b : _GEN_7181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7183 = 9'hc1 == r_count_23_io_out ? io_r_193_b : _GEN_7182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7184 = 9'hc2 == r_count_23_io_out ? io_r_194_b : _GEN_7183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7185 = 9'hc3 == r_count_23_io_out ? io_r_195_b : _GEN_7184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7186 = 9'hc4 == r_count_23_io_out ? io_r_196_b : _GEN_7185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7187 = 9'hc5 == r_count_23_io_out ? io_r_197_b : _GEN_7186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7188 = 9'hc6 == r_count_23_io_out ? io_r_198_b : _GEN_7187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7189 = 9'hc7 == r_count_23_io_out ? io_r_199_b : _GEN_7188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7190 = 9'hc8 == r_count_23_io_out ? io_r_200_b : _GEN_7189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7191 = 9'hc9 == r_count_23_io_out ? io_r_201_b : _GEN_7190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7192 = 9'hca == r_count_23_io_out ? io_r_202_b : _GEN_7191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7193 = 9'hcb == r_count_23_io_out ? io_r_203_b : _GEN_7192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7194 = 9'hcc == r_count_23_io_out ? io_r_204_b : _GEN_7193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7195 = 9'hcd == r_count_23_io_out ? io_r_205_b : _GEN_7194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7196 = 9'hce == r_count_23_io_out ? io_r_206_b : _GEN_7195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7197 = 9'hcf == r_count_23_io_out ? io_r_207_b : _GEN_7196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7198 = 9'hd0 == r_count_23_io_out ? io_r_208_b : _GEN_7197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7199 = 9'hd1 == r_count_23_io_out ? io_r_209_b : _GEN_7198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7200 = 9'hd2 == r_count_23_io_out ? io_r_210_b : _GEN_7199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7201 = 9'hd3 == r_count_23_io_out ? io_r_211_b : _GEN_7200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7202 = 9'hd4 == r_count_23_io_out ? io_r_212_b : _GEN_7201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7203 = 9'hd5 == r_count_23_io_out ? io_r_213_b : _GEN_7202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7204 = 9'hd6 == r_count_23_io_out ? io_r_214_b : _GEN_7203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7205 = 9'hd7 == r_count_23_io_out ? io_r_215_b : _GEN_7204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7206 = 9'hd8 == r_count_23_io_out ? io_r_216_b : _GEN_7205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7207 = 9'hd9 == r_count_23_io_out ? io_r_217_b : _GEN_7206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7208 = 9'hda == r_count_23_io_out ? io_r_218_b : _GEN_7207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7209 = 9'hdb == r_count_23_io_out ? io_r_219_b : _GEN_7208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7210 = 9'hdc == r_count_23_io_out ? io_r_220_b : _GEN_7209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7211 = 9'hdd == r_count_23_io_out ? io_r_221_b : _GEN_7210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7212 = 9'hde == r_count_23_io_out ? io_r_222_b : _GEN_7211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7213 = 9'hdf == r_count_23_io_out ? io_r_223_b : _GEN_7212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7214 = 9'he0 == r_count_23_io_out ? io_r_224_b : _GEN_7213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7215 = 9'he1 == r_count_23_io_out ? io_r_225_b : _GEN_7214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7216 = 9'he2 == r_count_23_io_out ? io_r_226_b : _GEN_7215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7217 = 9'he3 == r_count_23_io_out ? io_r_227_b : _GEN_7216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7218 = 9'he4 == r_count_23_io_out ? io_r_228_b : _GEN_7217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7219 = 9'he5 == r_count_23_io_out ? io_r_229_b : _GEN_7218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7220 = 9'he6 == r_count_23_io_out ? io_r_230_b : _GEN_7219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7221 = 9'he7 == r_count_23_io_out ? io_r_231_b : _GEN_7220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7222 = 9'he8 == r_count_23_io_out ? io_r_232_b : _GEN_7221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7223 = 9'he9 == r_count_23_io_out ? io_r_233_b : _GEN_7222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7224 = 9'hea == r_count_23_io_out ? io_r_234_b : _GEN_7223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7225 = 9'heb == r_count_23_io_out ? io_r_235_b : _GEN_7224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7226 = 9'hec == r_count_23_io_out ? io_r_236_b : _GEN_7225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7227 = 9'hed == r_count_23_io_out ? io_r_237_b : _GEN_7226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7228 = 9'hee == r_count_23_io_out ? io_r_238_b : _GEN_7227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7229 = 9'hef == r_count_23_io_out ? io_r_239_b : _GEN_7228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7230 = 9'hf0 == r_count_23_io_out ? io_r_240_b : _GEN_7229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7231 = 9'hf1 == r_count_23_io_out ? io_r_241_b : _GEN_7230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7232 = 9'hf2 == r_count_23_io_out ? io_r_242_b : _GEN_7231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7233 = 9'hf3 == r_count_23_io_out ? io_r_243_b : _GEN_7232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7234 = 9'hf4 == r_count_23_io_out ? io_r_244_b : _GEN_7233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7235 = 9'hf5 == r_count_23_io_out ? io_r_245_b : _GEN_7234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7236 = 9'hf6 == r_count_23_io_out ? io_r_246_b : _GEN_7235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7237 = 9'hf7 == r_count_23_io_out ? io_r_247_b : _GEN_7236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7238 = 9'hf8 == r_count_23_io_out ? io_r_248_b : _GEN_7237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7239 = 9'hf9 == r_count_23_io_out ? io_r_249_b : _GEN_7238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7240 = 9'hfa == r_count_23_io_out ? io_r_250_b : _GEN_7239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7241 = 9'hfb == r_count_23_io_out ? io_r_251_b : _GEN_7240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7242 = 9'hfc == r_count_23_io_out ? io_r_252_b : _GEN_7241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7243 = 9'hfd == r_count_23_io_out ? io_r_253_b : _GEN_7242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7244 = 9'hfe == r_count_23_io_out ? io_r_254_b : _GEN_7243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7245 = 9'hff == r_count_23_io_out ? io_r_255_b : _GEN_7244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7246 = 9'h100 == r_count_23_io_out ? io_r_256_b : _GEN_7245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7247 = 9'h101 == r_count_23_io_out ? io_r_257_b : _GEN_7246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7248 = 9'h102 == r_count_23_io_out ? io_r_258_b : _GEN_7247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7249 = 9'h103 == r_count_23_io_out ? io_r_259_b : _GEN_7248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7250 = 9'h104 == r_count_23_io_out ? io_r_260_b : _GEN_7249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7251 = 9'h105 == r_count_23_io_out ? io_r_261_b : _GEN_7250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7252 = 9'h106 == r_count_23_io_out ? io_r_262_b : _GEN_7251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7253 = 9'h107 == r_count_23_io_out ? io_r_263_b : _GEN_7252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7254 = 9'h108 == r_count_23_io_out ? io_r_264_b : _GEN_7253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7255 = 9'h109 == r_count_23_io_out ? io_r_265_b : _GEN_7254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7256 = 9'h10a == r_count_23_io_out ? io_r_266_b : _GEN_7255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7257 = 9'h10b == r_count_23_io_out ? io_r_267_b : _GEN_7256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7258 = 9'h10c == r_count_23_io_out ? io_r_268_b : _GEN_7257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7259 = 9'h10d == r_count_23_io_out ? io_r_269_b : _GEN_7258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7260 = 9'h10e == r_count_23_io_out ? io_r_270_b : _GEN_7259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7261 = 9'h10f == r_count_23_io_out ? io_r_271_b : _GEN_7260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7262 = 9'h110 == r_count_23_io_out ? io_r_272_b : _GEN_7261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7263 = 9'h111 == r_count_23_io_out ? io_r_273_b : _GEN_7262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7264 = 9'h112 == r_count_23_io_out ? io_r_274_b : _GEN_7263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7265 = 9'h113 == r_count_23_io_out ? io_r_275_b : _GEN_7264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7266 = 9'h114 == r_count_23_io_out ? io_r_276_b : _GEN_7265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7267 = 9'h115 == r_count_23_io_out ? io_r_277_b : _GEN_7266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7268 = 9'h116 == r_count_23_io_out ? io_r_278_b : _GEN_7267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7269 = 9'h117 == r_count_23_io_out ? io_r_279_b : _GEN_7268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7270 = 9'h118 == r_count_23_io_out ? io_r_280_b : _GEN_7269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7271 = 9'h119 == r_count_23_io_out ? io_r_281_b : _GEN_7270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7272 = 9'h11a == r_count_23_io_out ? io_r_282_b : _GEN_7271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7273 = 9'h11b == r_count_23_io_out ? io_r_283_b : _GEN_7272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7274 = 9'h11c == r_count_23_io_out ? io_r_284_b : _GEN_7273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7275 = 9'h11d == r_count_23_io_out ? io_r_285_b : _GEN_7274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7276 = 9'h11e == r_count_23_io_out ? io_r_286_b : _GEN_7275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7277 = 9'h11f == r_count_23_io_out ? io_r_287_b : _GEN_7276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7278 = 9'h120 == r_count_23_io_out ? io_r_288_b : _GEN_7277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7279 = 9'h121 == r_count_23_io_out ? io_r_289_b : _GEN_7278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7280 = 9'h122 == r_count_23_io_out ? io_r_290_b : _GEN_7279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7281 = 9'h123 == r_count_23_io_out ? io_r_291_b : _GEN_7280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7282 = 9'h124 == r_count_23_io_out ? io_r_292_b : _GEN_7281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7283 = 9'h125 == r_count_23_io_out ? io_r_293_b : _GEN_7282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7284 = 9'h126 == r_count_23_io_out ? io_r_294_b : _GEN_7283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7285 = 9'h127 == r_count_23_io_out ? io_r_295_b : _GEN_7284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7286 = 9'h128 == r_count_23_io_out ? io_r_296_b : _GEN_7285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7287 = 9'h129 == r_count_23_io_out ? io_r_297_b : _GEN_7286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7288 = 9'h12a == r_count_23_io_out ? io_r_298_b : _GEN_7287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7291 = 9'h1 == r_count_24_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7292 = 9'h2 == r_count_24_io_out ? io_r_2_b : _GEN_7291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7293 = 9'h3 == r_count_24_io_out ? io_r_3_b : _GEN_7292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7294 = 9'h4 == r_count_24_io_out ? io_r_4_b : _GEN_7293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7295 = 9'h5 == r_count_24_io_out ? io_r_5_b : _GEN_7294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7296 = 9'h6 == r_count_24_io_out ? io_r_6_b : _GEN_7295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7297 = 9'h7 == r_count_24_io_out ? io_r_7_b : _GEN_7296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7298 = 9'h8 == r_count_24_io_out ? io_r_8_b : _GEN_7297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7299 = 9'h9 == r_count_24_io_out ? io_r_9_b : _GEN_7298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7300 = 9'ha == r_count_24_io_out ? io_r_10_b : _GEN_7299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7301 = 9'hb == r_count_24_io_out ? io_r_11_b : _GEN_7300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7302 = 9'hc == r_count_24_io_out ? io_r_12_b : _GEN_7301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7303 = 9'hd == r_count_24_io_out ? io_r_13_b : _GEN_7302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7304 = 9'he == r_count_24_io_out ? io_r_14_b : _GEN_7303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7305 = 9'hf == r_count_24_io_out ? io_r_15_b : _GEN_7304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7306 = 9'h10 == r_count_24_io_out ? io_r_16_b : _GEN_7305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7307 = 9'h11 == r_count_24_io_out ? io_r_17_b : _GEN_7306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7308 = 9'h12 == r_count_24_io_out ? io_r_18_b : _GEN_7307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7309 = 9'h13 == r_count_24_io_out ? io_r_19_b : _GEN_7308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7310 = 9'h14 == r_count_24_io_out ? io_r_20_b : _GEN_7309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7311 = 9'h15 == r_count_24_io_out ? io_r_21_b : _GEN_7310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7312 = 9'h16 == r_count_24_io_out ? io_r_22_b : _GEN_7311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7313 = 9'h17 == r_count_24_io_out ? io_r_23_b : _GEN_7312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7314 = 9'h18 == r_count_24_io_out ? io_r_24_b : _GEN_7313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7315 = 9'h19 == r_count_24_io_out ? io_r_25_b : _GEN_7314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7316 = 9'h1a == r_count_24_io_out ? io_r_26_b : _GEN_7315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7317 = 9'h1b == r_count_24_io_out ? io_r_27_b : _GEN_7316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7318 = 9'h1c == r_count_24_io_out ? io_r_28_b : _GEN_7317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7319 = 9'h1d == r_count_24_io_out ? io_r_29_b : _GEN_7318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7320 = 9'h1e == r_count_24_io_out ? io_r_30_b : _GEN_7319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7321 = 9'h1f == r_count_24_io_out ? io_r_31_b : _GEN_7320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7322 = 9'h20 == r_count_24_io_out ? io_r_32_b : _GEN_7321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7323 = 9'h21 == r_count_24_io_out ? io_r_33_b : _GEN_7322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7324 = 9'h22 == r_count_24_io_out ? io_r_34_b : _GEN_7323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7325 = 9'h23 == r_count_24_io_out ? io_r_35_b : _GEN_7324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7326 = 9'h24 == r_count_24_io_out ? io_r_36_b : _GEN_7325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7327 = 9'h25 == r_count_24_io_out ? io_r_37_b : _GEN_7326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7328 = 9'h26 == r_count_24_io_out ? io_r_38_b : _GEN_7327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7329 = 9'h27 == r_count_24_io_out ? io_r_39_b : _GEN_7328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7330 = 9'h28 == r_count_24_io_out ? io_r_40_b : _GEN_7329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7331 = 9'h29 == r_count_24_io_out ? io_r_41_b : _GEN_7330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7332 = 9'h2a == r_count_24_io_out ? io_r_42_b : _GEN_7331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7333 = 9'h2b == r_count_24_io_out ? io_r_43_b : _GEN_7332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7334 = 9'h2c == r_count_24_io_out ? io_r_44_b : _GEN_7333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7335 = 9'h2d == r_count_24_io_out ? io_r_45_b : _GEN_7334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7336 = 9'h2e == r_count_24_io_out ? io_r_46_b : _GEN_7335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7337 = 9'h2f == r_count_24_io_out ? io_r_47_b : _GEN_7336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7338 = 9'h30 == r_count_24_io_out ? io_r_48_b : _GEN_7337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7339 = 9'h31 == r_count_24_io_out ? io_r_49_b : _GEN_7338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7340 = 9'h32 == r_count_24_io_out ? io_r_50_b : _GEN_7339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7341 = 9'h33 == r_count_24_io_out ? io_r_51_b : _GEN_7340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7342 = 9'h34 == r_count_24_io_out ? io_r_52_b : _GEN_7341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7343 = 9'h35 == r_count_24_io_out ? io_r_53_b : _GEN_7342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7344 = 9'h36 == r_count_24_io_out ? io_r_54_b : _GEN_7343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7345 = 9'h37 == r_count_24_io_out ? io_r_55_b : _GEN_7344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7346 = 9'h38 == r_count_24_io_out ? io_r_56_b : _GEN_7345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7347 = 9'h39 == r_count_24_io_out ? io_r_57_b : _GEN_7346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7348 = 9'h3a == r_count_24_io_out ? io_r_58_b : _GEN_7347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7349 = 9'h3b == r_count_24_io_out ? io_r_59_b : _GEN_7348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7350 = 9'h3c == r_count_24_io_out ? io_r_60_b : _GEN_7349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7351 = 9'h3d == r_count_24_io_out ? io_r_61_b : _GEN_7350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7352 = 9'h3e == r_count_24_io_out ? io_r_62_b : _GEN_7351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7353 = 9'h3f == r_count_24_io_out ? io_r_63_b : _GEN_7352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7354 = 9'h40 == r_count_24_io_out ? io_r_64_b : _GEN_7353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7355 = 9'h41 == r_count_24_io_out ? io_r_65_b : _GEN_7354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7356 = 9'h42 == r_count_24_io_out ? io_r_66_b : _GEN_7355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7357 = 9'h43 == r_count_24_io_out ? io_r_67_b : _GEN_7356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7358 = 9'h44 == r_count_24_io_out ? io_r_68_b : _GEN_7357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7359 = 9'h45 == r_count_24_io_out ? io_r_69_b : _GEN_7358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7360 = 9'h46 == r_count_24_io_out ? io_r_70_b : _GEN_7359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7361 = 9'h47 == r_count_24_io_out ? io_r_71_b : _GEN_7360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7362 = 9'h48 == r_count_24_io_out ? io_r_72_b : _GEN_7361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7363 = 9'h49 == r_count_24_io_out ? io_r_73_b : _GEN_7362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7364 = 9'h4a == r_count_24_io_out ? io_r_74_b : _GEN_7363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7365 = 9'h4b == r_count_24_io_out ? io_r_75_b : _GEN_7364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7366 = 9'h4c == r_count_24_io_out ? io_r_76_b : _GEN_7365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7367 = 9'h4d == r_count_24_io_out ? io_r_77_b : _GEN_7366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7368 = 9'h4e == r_count_24_io_out ? io_r_78_b : _GEN_7367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7369 = 9'h4f == r_count_24_io_out ? io_r_79_b : _GEN_7368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7370 = 9'h50 == r_count_24_io_out ? io_r_80_b : _GEN_7369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7371 = 9'h51 == r_count_24_io_out ? io_r_81_b : _GEN_7370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7372 = 9'h52 == r_count_24_io_out ? io_r_82_b : _GEN_7371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7373 = 9'h53 == r_count_24_io_out ? io_r_83_b : _GEN_7372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7374 = 9'h54 == r_count_24_io_out ? io_r_84_b : _GEN_7373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7375 = 9'h55 == r_count_24_io_out ? io_r_85_b : _GEN_7374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7376 = 9'h56 == r_count_24_io_out ? io_r_86_b : _GEN_7375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7377 = 9'h57 == r_count_24_io_out ? io_r_87_b : _GEN_7376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7378 = 9'h58 == r_count_24_io_out ? io_r_88_b : _GEN_7377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7379 = 9'h59 == r_count_24_io_out ? io_r_89_b : _GEN_7378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7380 = 9'h5a == r_count_24_io_out ? io_r_90_b : _GEN_7379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7381 = 9'h5b == r_count_24_io_out ? io_r_91_b : _GEN_7380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7382 = 9'h5c == r_count_24_io_out ? io_r_92_b : _GEN_7381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7383 = 9'h5d == r_count_24_io_out ? io_r_93_b : _GEN_7382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7384 = 9'h5e == r_count_24_io_out ? io_r_94_b : _GEN_7383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7385 = 9'h5f == r_count_24_io_out ? io_r_95_b : _GEN_7384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7386 = 9'h60 == r_count_24_io_out ? io_r_96_b : _GEN_7385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7387 = 9'h61 == r_count_24_io_out ? io_r_97_b : _GEN_7386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7388 = 9'h62 == r_count_24_io_out ? io_r_98_b : _GEN_7387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7389 = 9'h63 == r_count_24_io_out ? io_r_99_b : _GEN_7388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7390 = 9'h64 == r_count_24_io_out ? io_r_100_b : _GEN_7389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7391 = 9'h65 == r_count_24_io_out ? io_r_101_b : _GEN_7390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7392 = 9'h66 == r_count_24_io_out ? io_r_102_b : _GEN_7391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7393 = 9'h67 == r_count_24_io_out ? io_r_103_b : _GEN_7392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7394 = 9'h68 == r_count_24_io_out ? io_r_104_b : _GEN_7393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7395 = 9'h69 == r_count_24_io_out ? io_r_105_b : _GEN_7394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7396 = 9'h6a == r_count_24_io_out ? io_r_106_b : _GEN_7395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7397 = 9'h6b == r_count_24_io_out ? io_r_107_b : _GEN_7396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7398 = 9'h6c == r_count_24_io_out ? io_r_108_b : _GEN_7397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7399 = 9'h6d == r_count_24_io_out ? io_r_109_b : _GEN_7398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7400 = 9'h6e == r_count_24_io_out ? io_r_110_b : _GEN_7399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7401 = 9'h6f == r_count_24_io_out ? io_r_111_b : _GEN_7400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7402 = 9'h70 == r_count_24_io_out ? io_r_112_b : _GEN_7401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7403 = 9'h71 == r_count_24_io_out ? io_r_113_b : _GEN_7402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7404 = 9'h72 == r_count_24_io_out ? io_r_114_b : _GEN_7403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7405 = 9'h73 == r_count_24_io_out ? io_r_115_b : _GEN_7404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7406 = 9'h74 == r_count_24_io_out ? io_r_116_b : _GEN_7405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7407 = 9'h75 == r_count_24_io_out ? io_r_117_b : _GEN_7406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7408 = 9'h76 == r_count_24_io_out ? io_r_118_b : _GEN_7407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7409 = 9'h77 == r_count_24_io_out ? io_r_119_b : _GEN_7408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7410 = 9'h78 == r_count_24_io_out ? io_r_120_b : _GEN_7409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7411 = 9'h79 == r_count_24_io_out ? io_r_121_b : _GEN_7410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7412 = 9'h7a == r_count_24_io_out ? io_r_122_b : _GEN_7411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7413 = 9'h7b == r_count_24_io_out ? io_r_123_b : _GEN_7412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7414 = 9'h7c == r_count_24_io_out ? io_r_124_b : _GEN_7413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7415 = 9'h7d == r_count_24_io_out ? io_r_125_b : _GEN_7414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7416 = 9'h7e == r_count_24_io_out ? io_r_126_b : _GEN_7415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7417 = 9'h7f == r_count_24_io_out ? io_r_127_b : _GEN_7416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7418 = 9'h80 == r_count_24_io_out ? io_r_128_b : _GEN_7417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7419 = 9'h81 == r_count_24_io_out ? io_r_129_b : _GEN_7418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7420 = 9'h82 == r_count_24_io_out ? io_r_130_b : _GEN_7419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7421 = 9'h83 == r_count_24_io_out ? io_r_131_b : _GEN_7420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7422 = 9'h84 == r_count_24_io_out ? io_r_132_b : _GEN_7421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7423 = 9'h85 == r_count_24_io_out ? io_r_133_b : _GEN_7422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7424 = 9'h86 == r_count_24_io_out ? io_r_134_b : _GEN_7423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7425 = 9'h87 == r_count_24_io_out ? io_r_135_b : _GEN_7424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7426 = 9'h88 == r_count_24_io_out ? io_r_136_b : _GEN_7425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7427 = 9'h89 == r_count_24_io_out ? io_r_137_b : _GEN_7426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7428 = 9'h8a == r_count_24_io_out ? io_r_138_b : _GEN_7427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7429 = 9'h8b == r_count_24_io_out ? io_r_139_b : _GEN_7428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7430 = 9'h8c == r_count_24_io_out ? io_r_140_b : _GEN_7429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7431 = 9'h8d == r_count_24_io_out ? io_r_141_b : _GEN_7430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7432 = 9'h8e == r_count_24_io_out ? io_r_142_b : _GEN_7431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7433 = 9'h8f == r_count_24_io_out ? io_r_143_b : _GEN_7432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7434 = 9'h90 == r_count_24_io_out ? io_r_144_b : _GEN_7433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7435 = 9'h91 == r_count_24_io_out ? io_r_145_b : _GEN_7434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7436 = 9'h92 == r_count_24_io_out ? io_r_146_b : _GEN_7435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7437 = 9'h93 == r_count_24_io_out ? io_r_147_b : _GEN_7436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7438 = 9'h94 == r_count_24_io_out ? io_r_148_b : _GEN_7437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7439 = 9'h95 == r_count_24_io_out ? io_r_149_b : _GEN_7438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7440 = 9'h96 == r_count_24_io_out ? io_r_150_b : _GEN_7439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7441 = 9'h97 == r_count_24_io_out ? io_r_151_b : _GEN_7440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7442 = 9'h98 == r_count_24_io_out ? io_r_152_b : _GEN_7441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7443 = 9'h99 == r_count_24_io_out ? io_r_153_b : _GEN_7442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7444 = 9'h9a == r_count_24_io_out ? io_r_154_b : _GEN_7443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7445 = 9'h9b == r_count_24_io_out ? io_r_155_b : _GEN_7444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7446 = 9'h9c == r_count_24_io_out ? io_r_156_b : _GEN_7445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7447 = 9'h9d == r_count_24_io_out ? io_r_157_b : _GEN_7446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7448 = 9'h9e == r_count_24_io_out ? io_r_158_b : _GEN_7447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7449 = 9'h9f == r_count_24_io_out ? io_r_159_b : _GEN_7448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7450 = 9'ha0 == r_count_24_io_out ? io_r_160_b : _GEN_7449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7451 = 9'ha1 == r_count_24_io_out ? io_r_161_b : _GEN_7450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7452 = 9'ha2 == r_count_24_io_out ? io_r_162_b : _GEN_7451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7453 = 9'ha3 == r_count_24_io_out ? io_r_163_b : _GEN_7452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7454 = 9'ha4 == r_count_24_io_out ? io_r_164_b : _GEN_7453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7455 = 9'ha5 == r_count_24_io_out ? io_r_165_b : _GEN_7454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7456 = 9'ha6 == r_count_24_io_out ? io_r_166_b : _GEN_7455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7457 = 9'ha7 == r_count_24_io_out ? io_r_167_b : _GEN_7456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7458 = 9'ha8 == r_count_24_io_out ? io_r_168_b : _GEN_7457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7459 = 9'ha9 == r_count_24_io_out ? io_r_169_b : _GEN_7458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7460 = 9'haa == r_count_24_io_out ? io_r_170_b : _GEN_7459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7461 = 9'hab == r_count_24_io_out ? io_r_171_b : _GEN_7460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7462 = 9'hac == r_count_24_io_out ? io_r_172_b : _GEN_7461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7463 = 9'had == r_count_24_io_out ? io_r_173_b : _GEN_7462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7464 = 9'hae == r_count_24_io_out ? io_r_174_b : _GEN_7463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7465 = 9'haf == r_count_24_io_out ? io_r_175_b : _GEN_7464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7466 = 9'hb0 == r_count_24_io_out ? io_r_176_b : _GEN_7465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7467 = 9'hb1 == r_count_24_io_out ? io_r_177_b : _GEN_7466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7468 = 9'hb2 == r_count_24_io_out ? io_r_178_b : _GEN_7467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7469 = 9'hb3 == r_count_24_io_out ? io_r_179_b : _GEN_7468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7470 = 9'hb4 == r_count_24_io_out ? io_r_180_b : _GEN_7469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7471 = 9'hb5 == r_count_24_io_out ? io_r_181_b : _GEN_7470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7472 = 9'hb6 == r_count_24_io_out ? io_r_182_b : _GEN_7471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7473 = 9'hb7 == r_count_24_io_out ? io_r_183_b : _GEN_7472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7474 = 9'hb8 == r_count_24_io_out ? io_r_184_b : _GEN_7473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7475 = 9'hb9 == r_count_24_io_out ? io_r_185_b : _GEN_7474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7476 = 9'hba == r_count_24_io_out ? io_r_186_b : _GEN_7475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7477 = 9'hbb == r_count_24_io_out ? io_r_187_b : _GEN_7476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7478 = 9'hbc == r_count_24_io_out ? io_r_188_b : _GEN_7477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7479 = 9'hbd == r_count_24_io_out ? io_r_189_b : _GEN_7478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7480 = 9'hbe == r_count_24_io_out ? io_r_190_b : _GEN_7479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7481 = 9'hbf == r_count_24_io_out ? io_r_191_b : _GEN_7480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7482 = 9'hc0 == r_count_24_io_out ? io_r_192_b : _GEN_7481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7483 = 9'hc1 == r_count_24_io_out ? io_r_193_b : _GEN_7482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7484 = 9'hc2 == r_count_24_io_out ? io_r_194_b : _GEN_7483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7485 = 9'hc3 == r_count_24_io_out ? io_r_195_b : _GEN_7484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7486 = 9'hc4 == r_count_24_io_out ? io_r_196_b : _GEN_7485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7487 = 9'hc5 == r_count_24_io_out ? io_r_197_b : _GEN_7486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7488 = 9'hc6 == r_count_24_io_out ? io_r_198_b : _GEN_7487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7489 = 9'hc7 == r_count_24_io_out ? io_r_199_b : _GEN_7488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7490 = 9'hc8 == r_count_24_io_out ? io_r_200_b : _GEN_7489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7491 = 9'hc9 == r_count_24_io_out ? io_r_201_b : _GEN_7490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7492 = 9'hca == r_count_24_io_out ? io_r_202_b : _GEN_7491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7493 = 9'hcb == r_count_24_io_out ? io_r_203_b : _GEN_7492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7494 = 9'hcc == r_count_24_io_out ? io_r_204_b : _GEN_7493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7495 = 9'hcd == r_count_24_io_out ? io_r_205_b : _GEN_7494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7496 = 9'hce == r_count_24_io_out ? io_r_206_b : _GEN_7495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7497 = 9'hcf == r_count_24_io_out ? io_r_207_b : _GEN_7496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7498 = 9'hd0 == r_count_24_io_out ? io_r_208_b : _GEN_7497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7499 = 9'hd1 == r_count_24_io_out ? io_r_209_b : _GEN_7498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7500 = 9'hd2 == r_count_24_io_out ? io_r_210_b : _GEN_7499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7501 = 9'hd3 == r_count_24_io_out ? io_r_211_b : _GEN_7500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7502 = 9'hd4 == r_count_24_io_out ? io_r_212_b : _GEN_7501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7503 = 9'hd5 == r_count_24_io_out ? io_r_213_b : _GEN_7502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7504 = 9'hd6 == r_count_24_io_out ? io_r_214_b : _GEN_7503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7505 = 9'hd7 == r_count_24_io_out ? io_r_215_b : _GEN_7504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7506 = 9'hd8 == r_count_24_io_out ? io_r_216_b : _GEN_7505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7507 = 9'hd9 == r_count_24_io_out ? io_r_217_b : _GEN_7506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7508 = 9'hda == r_count_24_io_out ? io_r_218_b : _GEN_7507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7509 = 9'hdb == r_count_24_io_out ? io_r_219_b : _GEN_7508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7510 = 9'hdc == r_count_24_io_out ? io_r_220_b : _GEN_7509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7511 = 9'hdd == r_count_24_io_out ? io_r_221_b : _GEN_7510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7512 = 9'hde == r_count_24_io_out ? io_r_222_b : _GEN_7511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7513 = 9'hdf == r_count_24_io_out ? io_r_223_b : _GEN_7512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7514 = 9'he0 == r_count_24_io_out ? io_r_224_b : _GEN_7513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7515 = 9'he1 == r_count_24_io_out ? io_r_225_b : _GEN_7514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7516 = 9'he2 == r_count_24_io_out ? io_r_226_b : _GEN_7515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7517 = 9'he3 == r_count_24_io_out ? io_r_227_b : _GEN_7516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7518 = 9'he4 == r_count_24_io_out ? io_r_228_b : _GEN_7517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7519 = 9'he5 == r_count_24_io_out ? io_r_229_b : _GEN_7518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7520 = 9'he6 == r_count_24_io_out ? io_r_230_b : _GEN_7519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7521 = 9'he7 == r_count_24_io_out ? io_r_231_b : _GEN_7520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7522 = 9'he8 == r_count_24_io_out ? io_r_232_b : _GEN_7521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7523 = 9'he9 == r_count_24_io_out ? io_r_233_b : _GEN_7522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7524 = 9'hea == r_count_24_io_out ? io_r_234_b : _GEN_7523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7525 = 9'heb == r_count_24_io_out ? io_r_235_b : _GEN_7524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7526 = 9'hec == r_count_24_io_out ? io_r_236_b : _GEN_7525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7527 = 9'hed == r_count_24_io_out ? io_r_237_b : _GEN_7526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7528 = 9'hee == r_count_24_io_out ? io_r_238_b : _GEN_7527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7529 = 9'hef == r_count_24_io_out ? io_r_239_b : _GEN_7528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7530 = 9'hf0 == r_count_24_io_out ? io_r_240_b : _GEN_7529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7531 = 9'hf1 == r_count_24_io_out ? io_r_241_b : _GEN_7530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7532 = 9'hf2 == r_count_24_io_out ? io_r_242_b : _GEN_7531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7533 = 9'hf3 == r_count_24_io_out ? io_r_243_b : _GEN_7532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7534 = 9'hf4 == r_count_24_io_out ? io_r_244_b : _GEN_7533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7535 = 9'hf5 == r_count_24_io_out ? io_r_245_b : _GEN_7534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7536 = 9'hf6 == r_count_24_io_out ? io_r_246_b : _GEN_7535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7537 = 9'hf7 == r_count_24_io_out ? io_r_247_b : _GEN_7536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7538 = 9'hf8 == r_count_24_io_out ? io_r_248_b : _GEN_7537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7539 = 9'hf9 == r_count_24_io_out ? io_r_249_b : _GEN_7538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7540 = 9'hfa == r_count_24_io_out ? io_r_250_b : _GEN_7539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7541 = 9'hfb == r_count_24_io_out ? io_r_251_b : _GEN_7540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7542 = 9'hfc == r_count_24_io_out ? io_r_252_b : _GEN_7541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7543 = 9'hfd == r_count_24_io_out ? io_r_253_b : _GEN_7542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7544 = 9'hfe == r_count_24_io_out ? io_r_254_b : _GEN_7543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7545 = 9'hff == r_count_24_io_out ? io_r_255_b : _GEN_7544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7546 = 9'h100 == r_count_24_io_out ? io_r_256_b : _GEN_7545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7547 = 9'h101 == r_count_24_io_out ? io_r_257_b : _GEN_7546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7548 = 9'h102 == r_count_24_io_out ? io_r_258_b : _GEN_7547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7549 = 9'h103 == r_count_24_io_out ? io_r_259_b : _GEN_7548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7550 = 9'h104 == r_count_24_io_out ? io_r_260_b : _GEN_7549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7551 = 9'h105 == r_count_24_io_out ? io_r_261_b : _GEN_7550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7552 = 9'h106 == r_count_24_io_out ? io_r_262_b : _GEN_7551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7553 = 9'h107 == r_count_24_io_out ? io_r_263_b : _GEN_7552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7554 = 9'h108 == r_count_24_io_out ? io_r_264_b : _GEN_7553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7555 = 9'h109 == r_count_24_io_out ? io_r_265_b : _GEN_7554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7556 = 9'h10a == r_count_24_io_out ? io_r_266_b : _GEN_7555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7557 = 9'h10b == r_count_24_io_out ? io_r_267_b : _GEN_7556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7558 = 9'h10c == r_count_24_io_out ? io_r_268_b : _GEN_7557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7559 = 9'h10d == r_count_24_io_out ? io_r_269_b : _GEN_7558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7560 = 9'h10e == r_count_24_io_out ? io_r_270_b : _GEN_7559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7561 = 9'h10f == r_count_24_io_out ? io_r_271_b : _GEN_7560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7562 = 9'h110 == r_count_24_io_out ? io_r_272_b : _GEN_7561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7563 = 9'h111 == r_count_24_io_out ? io_r_273_b : _GEN_7562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7564 = 9'h112 == r_count_24_io_out ? io_r_274_b : _GEN_7563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7565 = 9'h113 == r_count_24_io_out ? io_r_275_b : _GEN_7564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7566 = 9'h114 == r_count_24_io_out ? io_r_276_b : _GEN_7565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7567 = 9'h115 == r_count_24_io_out ? io_r_277_b : _GEN_7566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7568 = 9'h116 == r_count_24_io_out ? io_r_278_b : _GEN_7567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7569 = 9'h117 == r_count_24_io_out ? io_r_279_b : _GEN_7568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7570 = 9'h118 == r_count_24_io_out ? io_r_280_b : _GEN_7569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7571 = 9'h119 == r_count_24_io_out ? io_r_281_b : _GEN_7570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7572 = 9'h11a == r_count_24_io_out ? io_r_282_b : _GEN_7571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7573 = 9'h11b == r_count_24_io_out ? io_r_283_b : _GEN_7572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7574 = 9'h11c == r_count_24_io_out ? io_r_284_b : _GEN_7573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7575 = 9'h11d == r_count_24_io_out ? io_r_285_b : _GEN_7574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7576 = 9'h11e == r_count_24_io_out ? io_r_286_b : _GEN_7575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7577 = 9'h11f == r_count_24_io_out ? io_r_287_b : _GEN_7576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7578 = 9'h120 == r_count_24_io_out ? io_r_288_b : _GEN_7577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7579 = 9'h121 == r_count_24_io_out ? io_r_289_b : _GEN_7578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7580 = 9'h122 == r_count_24_io_out ? io_r_290_b : _GEN_7579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7581 = 9'h123 == r_count_24_io_out ? io_r_291_b : _GEN_7580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7582 = 9'h124 == r_count_24_io_out ? io_r_292_b : _GEN_7581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7583 = 9'h125 == r_count_24_io_out ? io_r_293_b : _GEN_7582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7584 = 9'h126 == r_count_24_io_out ? io_r_294_b : _GEN_7583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7585 = 9'h127 == r_count_24_io_out ? io_r_295_b : _GEN_7584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7586 = 9'h128 == r_count_24_io_out ? io_r_296_b : _GEN_7585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7587 = 9'h129 == r_count_24_io_out ? io_r_297_b : _GEN_7586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7588 = 9'h12a == r_count_24_io_out ? io_r_298_b : _GEN_7587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7591 = 9'h1 == r_count_25_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7592 = 9'h2 == r_count_25_io_out ? io_r_2_b : _GEN_7591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7593 = 9'h3 == r_count_25_io_out ? io_r_3_b : _GEN_7592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7594 = 9'h4 == r_count_25_io_out ? io_r_4_b : _GEN_7593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7595 = 9'h5 == r_count_25_io_out ? io_r_5_b : _GEN_7594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7596 = 9'h6 == r_count_25_io_out ? io_r_6_b : _GEN_7595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7597 = 9'h7 == r_count_25_io_out ? io_r_7_b : _GEN_7596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7598 = 9'h8 == r_count_25_io_out ? io_r_8_b : _GEN_7597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7599 = 9'h9 == r_count_25_io_out ? io_r_9_b : _GEN_7598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7600 = 9'ha == r_count_25_io_out ? io_r_10_b : _GEN_7599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7601 = 9'hb == r_count_25_io_out ? io_r_11_b : _GEN_7600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7602 = 9'hc == r_count_25_io_out ? io_r_12_b : _GEN_7601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7603 = 9'hd == r_count_25_io_out ? io_r_13_b : _GEN_7602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7604 = 9'he == r_count_25_io_out ? io_r_14_b : _GEN_7603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7605 = 9'hf == r_count_25_io_out ? io_r_15_b : _GEN_7604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7606 = 9'h10 == r_count_25_io_out ? io_r_16_b : _GEN_7605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7607 = 9'h11 == r_count_25_io_out ? io_r_17_b : _GEN_7606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7608 = 9'h12 == r_count_25_io_out ? io_r_18_b : _GEN_7607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7609 = 9'h13 == r_count_25_io_out ? io_r_19_b : _GEN_7608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7610 = 9'h14 == r_count_25_io_out ? io_r_20_b : _GEN_7609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7611 = 9'h15 == r_count_25_io_out ? io_r_21_b : _GEN_7610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7612 = 9'h16 == r_count_25_io_out ? io_r_22_b : _GEN_7611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7613 = 9'h17 == r_count_25_io_out ? io_r_23_b : _GEN_7612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7614 = 9'h18 == r_count_25_io_out ? io_r_24_b : _GEN_7613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7615 = 9'h19 == r_count_25_io_out ? io_r_25_b : _GEN_7614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7616 = 9'h1a == r_count_25_io_out ? io_r_26_b : _GEN_7615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7617 = 9'h1b == r_count_25_io_out ? io_r_27_b : _GEN_7616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7618 = 9'h1c == r_count_25_io_out ? io_r_28_b : _GEN_7617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7619 = 9'h1d == r_count_25_io_out ? io_r_29_b : _GEN_7618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7620 = 9'h1e == r_count_25_io_out ? io_r_30_b : _GEN_7619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7621 = 9'h1f == r_count_25_io_out ? io_r_31_b : _GEN_7620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7622 = 9'h20 == r_count_25_io_out ? io_r_32_b : _GEN_7621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7623 = 9'h21 == r_count_25_io_out ? io_r_33_b : _GEN_7622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7624 = 9'h22 == r_count_25_io_out ? io_r_34_b : _GEN_7623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7625 = 9'h23 == r_count_25_io_out ? io_r_35_b : _GEN_7624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7626 = 9'h24 == r_count_25_io_out ? io_r_36_b : _GEN_7625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7627 = 9'h25 == r_count_25_io_out ? io_r_37_b : _GEN_7626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7628 = 9'h26 == r_count_25_io_out ? io_r_38_b : _GEN_7627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7629 = 9'h27 == r_count_25_io_out ? io_r_39_b : _GEN_7628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7630 = 9'h28 == r_count_25_io_out ? io_r_40_b : _GEN_7629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7631 = 9'h29 == r_count_25_io_out ? io_r_41_b : _GEN_7630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7632 = 9'h2a == r_count_25_io_out ? io_r_42_b : _GEN_7631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7633 = 9'h2b == r_count_25_io_out ? io_r_43_b : _GEN_7632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7634 = 9'h2c == r_count_25_io_out ? io_r_44_b : _GEN_7633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7635 = 9'h2d == r_count_25_io_out ? io_r_45_b : _GEN_7634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7636 = 9'h2e == r_count_25_io_out ? io_r_46_b : _GEN_7635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7637 = 9'h2f == r_count_25_io_out ? io_r_47_b : _GEN_7636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7638 = 9'h30 == r_count_25_io_out ? io_r_48_b : _GEN_7637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7639 = 9'h31 == r_count_25_io_out ? io_r_49_b : _GEN_7638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7640 = 9'h32 == r_count_25_io_out ? io_r_50_b : _GEN_7639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7641 = 9'h33 == r_count_25_io_out ? io_r_51_b : _GEN_7640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7642 = 9'h34 == r_count_25_io_out ? io_r_52_b : _GEN_7641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7643 = 9'h35 == r_count_25_io_out ? io_r_53_b : _GEN_7642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7644 = 9'h36 == r_count_25_io_out ? io_r_54_b : _GEN_7643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7645 = 9'h37 == r_count_25_io_out ? io_r_55_b : _GEN_7644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7646 = 9'h38 == r_count_25_io_out ? io_r_56_b : _GEN_7645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7647 = 9'h39 == r_count_25_io_out ? io_r_57_b : _GEN_7646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7648 = 9'h3a == r_count_25_io_out ? io_r_58_b : _GEN_7647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7649 = 9'h3b == r_count_25_io_out ? io_r_59_b : _GEN_7648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7650 = 9'h3c == r_count_25_io_out ? io_r_60_b : _GEN_7649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7651 = 9'h3d == r_count_25_io_out ? io_r_61_b : _GEN_7650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7652 = 9'h3e == r_count_25_io_out ? io_r_62_b : _GEN_7651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7653 = 9'h3f == r_count_25_io_out ? io_r_63_b : _GEN_7652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7654 = 9'h40 == r_count_25_io_out ? io_r_64_b : _GEN_7653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7655 = 9'h41 == r_count_25_io_out ? io_r_65_b : _GEN_7654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7656 = 9'h42 == r_count_25_io_out ? io_r_66_b : _GEN_7655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7657 = 9'h43 == r_count_25_io_out ? io_r_67_b : _GEN_7656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7658 = 9'h44 == r_count_25_io_out ? io_r_68_b : _GEN_7657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7659 = 9'h45 == r_count_25_io_out ? io_r_69_b : _GEN_7658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7660 = 9'h46 == r_count_25_io_out ? io_r_70_b : _GEN_7659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7661 = 9'h47 == r_count_25_io_out ? io_r_71_b : _GEN_7660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7662 = 9'h48 == r_count_25_io_out ? io_r_72_b : _GEN_7661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7663 = 9'h49 == r_count_25_io_out ? io_r_73_b : _GEN_7662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7664 = 9'h4a == r_count_25_io_out ? io_r_74_b : _GEN_7663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7665 = 9'h4b == r_count_25_io_out ? io_r_75_b : _GEN_7664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7666 = 9'h4c == r_count_25_io_out ? io_r_76_b : _GEN_7665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7667 = 9'h4d == r_count_25_io_out ? io_r_77_b : _GEN_7666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7668 = 9'h4e == r_count_25_io_out ? io_r_78_b : _GEN_7667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7669 = 9'h4f == r_count_25_io_out ? io_r_79_b : _GEN_7668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7670 = 9'h50 == r_count_25_io_out ? io_r_80_b : _GEN_7669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7671 = 9'h51 == r_count_25_io_out ? io_r_81_b : _GEN_7670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7672 = 9'h52 == r_count_25_io_out ? io_r_82_b : _GEN_7671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7673 = 9'h53 == r_count_25_io_out ? io_r_83_b : _GEN_7672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7674 = 9'h54 == r_count_25_io_out ? io_r_84_b : _GEN_7673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7675 = 9'h55 == r_count_25_io_out ? io_r_85_b : _GEN_7674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7676 = 9'h56 == r_count_25_io_out ? io_r_86_b : _GEN_7675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7677 = 9'h57 == r_count_25_io_out ? io_r_87_b : _GEN_7676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7678 = 9'h58 == r_count_25_io_out ? io_r_88_b : _GEN_7677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7679 = 9'h59 == r_count_25_io_out ? io_r_89_b : _GEN_7678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7680 = 9'h5a == r_count_25_io_out ? io_r_90_b : _GEN_7679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7681 = 9'h5b == r_count_25_io_out ? io_r_91_b : _GEN_7680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7682 = 9'h5c == r_count_25_io_out ? io_r_92_b : _GEN_7681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7683 = 9'h5d == r_count_25_io_out ? io_r_93_b : _GEN_7682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7684 = 9'h5e == r_count_25_io_out ? io_r_94_b : _GEN_7683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7685 = 9'h5f == r_count_25_io_out ? io_r_95_b : _GEN_7684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7686 = 9'h60 == r_count_25_io_out ? io_r_96_b : _GEN_7685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7687 = 9'h61 == r_count_25_io_out ? io_r_97_b : _GEN_7686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7688 = 9'h62 == r_count_25_io_out ? io_r_98_b : _GEN_7687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7689 = 9'h63 == r_count_25_io_out ? io_r_99_b : _GEN_7688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7690 = 9'h64 == r_count_25_io_out ? io_r_100_b : _GEN_7689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7691 = 9'h65 == r_count_25_io_out ? io_r_101_b : _GEN_7690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7692 = 9'h66 == r_count_25_io_out ? io_r_102_b : _GEN_7691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7693 = 9'h67 == r_count_25_io_out ? io_r_103_b : _GEN_7692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7694 = 9'h68 == r_count_25_io_out ? io_r_104_b : _GEN_7693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7695 = 9'h69 == r_count_25_io_out ? io_r_105_b : _GEN_7694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7696 = 9'h6a == r_count_25_io_out ? io_r_106_b : _GEN_7695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7697 = 9'h6b == r_count_25_io_out ? io_r_107_b : _GEN_7696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7698 = 9'h6c == r_count_25_io_out ? io_r_108_b : _GEN_7697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7699 = 9'h6d == r_count_25_io_out ? io_r_109_b : _GEN_7698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7700 = 9'h6e == r_count_25_io_out ? io_r_110_b : _GEN_7699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7701 = 9'h6f == r_count_25_io_out ? io_r_111_b : _GEN_7700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7702 = 9'h70 == r_count_25_io_out ? io_r_112_b : _GEN_7701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7703 = 9'h71 == r_count_25_io_out ? io_r_113_b : _GEN_7702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7704 = 9'h72 == r_count_25_io_out ? io_r_114_b : _GEN_7703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7705 = 9'h73 == r_count_25_io_out ? io_r_115_b : _GEN_7704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7706 = 9'h74 == r_count_25_io_out ? io_r_116_b : _GEN_7705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7707 = 9'h75 == r_count_25_io_out ? io_r_117_b : _GEN_7706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7708 = 9'h76 == r_count_25_io_out ? io_r_118_b : _GEN_7707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7709 = 9'h77 == r_count_25_io_out ? io_r_119_b : _GEN_7708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7710 = 9'h78 == r_count_25_io_out ? io_r_120_b : _GEN_7709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7711 = 9'h79 == r_count_25_io_out ? io_r_121_b : _GEN_7710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7712 = 9'h7a == r_count_25_io_out ? io_r_122_b : _GEN_7711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7713 = 9'h7b == r_count_25_io_out ? io_r_123_b : _GEN_7712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7714 = 9'h7c == r_count_25_io_out ? io_r_124_b : _GEN_7713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7715 = 9'h7d == r_count_25_io_out ? io_r_125_b : _GEN_7714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7716 = 9'h7e == r_count_25_io_out ? io_r_126_b : _GEN_7715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7717 = 9'h7f == r_count_25_io_out ? io_r_127_b : _GEN_7716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7718 = 9'h80 == r_count_25_io_out ? io_r_128_b : _GEN_7717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7719 = 9'h81 == r_count_25_io_out ? io_r_129_b : _GEN_7718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7720 = 9'h82 == r_count_25_io_out ? io_r_130_b : _GEN_7719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7721 = 9'h83 == r_count_25_io_out ? io_r_131_b : _GEN_7720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7722 = 9'h84 == r_count_25_io_out ? io_r_132_b : _GEN_7721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7723 = 9'h85 == r_count_25_io_out ? io_r_133_b : _GEN_7722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7724 = 9'h86 == r_count_25_io_out ? io_r_134_b : _GEN_7723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7725 = 9'h87 == r_count_25_io_out ? io_r_135_b : _GEN_7724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7726 = 9'h88 == r_count_25_io_out ? io_r_136_b : _GEN_7725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7727 = 9'h89 == r_count_25_io_out ? io_r_137_b : _GEN_7726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7728 = 9'h8a == r_count_25_io_out ? io_r_138_b : _GEN_7727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7729 = 9'h8b == r_count_25_io_out ? io_r_139_b : _GEN_7728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7730 = 9'h8c == r_count_25_io_out ? io_r_140_b : _GEN_7729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7731 = 9'h8d == r_count_25_io_out ? io_r_141_b : _GEN_7730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7732 = 9'h8e == r_count_25_io_out ? io_r_142_b : _GEN_7731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7733 = 9'h8f == r_count_25_io_out ? io_r_143_b : _GEN_7732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7734 = 9'h90 == r_count_25_io_out ? io_r_144_b : _GEN_7733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7735 = 9'h91 == r_count_25_io_out ? io_r_145_b : _GEN_7734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7736 = 9'h92 == r_count_25_io_out ? io_r_146_b : _GEN_7735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7737 = 9'h93 == r_count_25_io_out ? io_r_147_b : _GEN_7736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7738 = 9'h94 == r_count_25_io_out ? io_r_148_b : _GEN_7737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7739 = 9'h95 == r_count_25_io_out ? io_r_149_b : _GEN_7738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7740 = 9'h96 == r_count_25_io_out ? io_r_150_b : _GEN_7739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7741 = 9'h97 == r_count_25_io_out ? io_r_151_b : _GEN_7740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7742 = 9'h98 == r_count_25_io_out ? io_r_152_b : _GEN_7741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7743 = 9'h99 == r_count_25_io_out ? io_r_153_b : _GEN_7742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7744 = 9'h9a == r_count_25_io_out ? io_r_154_b : _GEN_7743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7745 = 9'h9b == r_count_25_io_out ? io_r_155_b : _GEN_7744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7746 = 9'h9c == r_count_25_io_out ? io_r_156_b : _GEN_7745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7747 = 9'h9d == r_count_25_io_out ? io_r_157_b : _GEN_7746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7748 = 9'h9e == r_count_25_io_out ? io_r_158_b : _GEN_7747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7749 = 9'h9f == r_count_25_io_out ? io_r_159_b : _GEN_7748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7750 = 9'ha0 == r_count_25_io_out ? io_r_160_b : _GEN_7749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7751 = 9'ha1 == r_count_25_io_out ? io_r_161_b : _GEN_7750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7752 = 9'ha2 == r_count_25_io_out ? io_r_162_b : _GEN_7751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7753 = 9'ha3 == r_count_25_io_out ? io_r_163_b : _GEN_7752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7754 = 9'ha4 == r_count_25_io_out ? io_r_164_b : _GEN_7753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7755 = 9'ha5 == r_count_25_io_out ? io_r_165_b : _GEN_7754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7756 = 9'ha6 == r_count_25_io_out ? io_r_166_b : _GEN_7755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7757 = 9'ha7 == r_count_25_io_out ? io_r_167_b : _GEN_7756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7758 = 9'ha8 == r_count_25_io_out ? io_r_168_b : _GEN_7757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7759 = 9'ha9 == r_count_25_io_out ? io_r_169_b : _GEN_7758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7760 = 9'haa == r_count_25_io_out ? io_r_170_b : _GEN_7759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7761 = 9'hab == r_count_25_io_out ? io_r_171_b : _GEN_7760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7762 = 9'hac == r_count_25_io_out ? io_r_172_b : _GEN_7761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7763 = 9'had == r_count_25_io_out ? io_r_173_b : _GEN_7762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7764 = 9'hae == r_count_25_io_out ? io_r_174_b : _GEN_7763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7765 = 9'haf == r_count_25_io_out ? io_r_175_b : _GEN_7764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7766 = 9'hb0 == r_count_25_io_out ? io_r_176_b : _GEN_7765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7767 = 9'hb1 == r_count_25_io_out ? io_r_177_b : _GEN_7766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7768 = 9'hb2 == r_count_25_io_out ? io_r_178_b : _GEN_7767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7769 = 9'hb3 == r_count_25_io_out ? io_r_179_b : _GEN_7768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7770 = 9'hb4 == r_count_25_io_out ? io_r_180_b : _GEN_7769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7771 = 9'hb5 == r_count_25_io_out ? io_r_181_b : _GEN_7770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7772 = 9'hb6 == r_count_25_io_out ? io_r_182_b : _GEN_7771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7773 = 9'hb7 == r_count_25_io_out ? io_r_183_b : _GEN_7772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7774 = 9'hb8 == r_count_25_io_out ? io_r_184_b : _GEN_7773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7775 = 9'hb9 == r_count_25_io_out ? io_r_185_b : _GEN_7774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7776 = 9'hba == r_count_25_io_out ? io_r_186_b : _GEN_7775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7777 = 9'hbb == r_count_25_io_out ? io_r_187_b : _GEN_7776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7778 = 9'hbc == r_count_25_io_out ? io_r_188_b : _GEN_7777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7779 = 9'hbd == r_count_25_io_out ? io_r_189_b : _GEN_7778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7780 = 9'hbe == r_count_25_io_out ? io_r_190_b : _GEN_7779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7781 = 9'hbf == r_count_25_io_out ? io_r_191_b : _GEN_7780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7782 = 9'hc0 == r_count_25_io_out ? io_r_192_b : _GEN_7781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7783 = 9'hc1 == r_count_25_io_out ? io_r_193_b : _GEN_7782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7784 = 9'hc2 == r_count_25_io_out ? io_r_194_b : _GEN_7783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7785 = 9'hc3 == r_count_25_io_out ? io_r_195_b : _GEN_7784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7786 = 9'hc4 == r_count_25_io_out ? io_r_196_b : _GEN_7785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7787 = 9'hc5 == r_count_25_io_out ? io_r_197_b : _GEN_7786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7788 = 9'hc6 == r_count_25_io_out ? io_r_198_b : _GEN_7787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7789 = 9'hc7 == r_count_25_io_out ? io_r_199_b : _GEN_7788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7790 = 9'hc8 == r_count_25_io_out ? io_r_200_b : _GEN_7789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7791 = 9'hc9 == r_count_25_io_out ? io_r_201_b : _GEN_7790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7792 = 9'hca == r_count_25_io_out ? io_r_202_b : _GEN_7791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7793 = 9'hcb == r_count_25_io_out ? io_r_203_b : _GEN_7792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7794 = 9'hcc == r_count_25_io_out ? io_r_204_b : _GEN_7793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7795 = 9'hcd == r_count_25_io_out ? io_r_205_b : _GEN_7794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7796 = 9'hce == r_count_25_io_out ? io_r_206_b : _GEN_7795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7797 = 9'hcf == r_count_25_io_out ? io_r_207_b : _GEN_7796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7798 = 9'hd0 == r_count_25_io_out ? io_r_208_b : _GEN_7797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7799 = 9'hd1 == r_count_25_io_out ? io_r_209_b : _GEN_7798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7800 = 9'hd2 == r_count_25_io_out ? io_r_210_b : _GEN_7799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7801 = 9'hd3 == r_count_25_io_out ? io_r_211_b : _GEN_7800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7802 = 9'hd4 == r_count_25_io_out ? io_r_212_b : _GEN_7801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7803 = 9'hd5 == r_count_25_io_out ? io_r_213_b : _GEN_7802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7804 = 9'hd6 == r_count_25_io_out ? io_r_214_b : _GEN_7803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7805 = 9'hd7 == r_count_25_io_out ? io_r_215_b : _GEN_7804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7806 = 9'hd8 == r_count_25_io_out ? io_r_216_b : _GEN_7805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7807 = 9'hd9 == r_count_25_io_out ? io_r_217_b : _GEN_7806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7808 = 9'hda == r_count_25_io_out ? io_r_218_b : _GEN_7807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7809 = 9'hdb == r_count_25_io_out ? io_r_219_b : _GEN_7808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7810 = 9'hdc == r_count_25_io_out ? io_r_220_b : _GEN_7809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7811 = 9'hdd == r_count_25_io_out ? io_r_221_b : _GEN_7810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7812 = 9'hde == r_count_25_io_out ? io_r_222_b : _GEN_7811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7813 = 9'hdf == r_count_25_io_out ? io_r_223_b : _GEN_7812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7814 = 9'he0 == r_count_25_io_out ? io_r_224_b : _GEN_7813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7815 = 9'he1 == r_count_25_io_out ? io_r_225_b : _GEN_7814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7816 = 9'he2 == r_count_25_io_out ? io_r_226_b : _GEN_7815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7817 = 9'he3 == r_count_25_io_out ? io_r_227_b : _GEN_7816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7818 = 9'he4 == r_count_25_io_out ? io_r_228_b : _GEN_7817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7819 = 9'he5 == r_count_25_io_out ? io_r_229_b : _GEN_7818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7820 = 9'he6 == r_count_25_io_out ? io_r_230_b : _GEN_7819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7821 = 9'he7 == r_count_25_io_out ? io_r_231_b : _GEN_7820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7822 = 9'he8 == r_count_25_io_out ? io_r_232_b : _GEN_7821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7823 = 9'he9 == r_count_25_io_out ? io_r_233_b : _GEN_7822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7824 = 9'hea == r_count_25_io_out ? io_r_234_b : _GEN_7823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7825 = 9'heb == r_count_25_io_out ? io_r_235_b : _GEN_7824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7826 = 9'hec == r_count_25_io_out ? io_r_236_b : _GEN_7825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7827 = 9'hed == r_count_25_io_out ? io_r_237_b : _GEN_7826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7828 = 9'hee == r_count_25_io_out ? io_r_238_b : _GEN_7827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7829 = 9'hef == r_count_25_io_out ? io_r_239_b : _GEN_7828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7830 = 9'hf0 == r_count_25_io_out ? io_r_240_b : _GEN_7829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7831 = 9'hf1 == r_count_25_io_out ? io_r_241_b : _GEN_7830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7832 = 9'hf2 == r_count_25_io_out ? io_r_242_b : _GEN_7831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7833 = 9'hf3 == r_count_25_io_out ? io_r_243_b : _GEN_7832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7834 = 9'hf4 == r_count_25_io_out ? io_r_244_b : _GEN_7833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7835 = 9'hf5 == r_count_25_io_out ? io_r_245_b : _GEN_7834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7836 = 9'hf6 == r_count_25_io_out ? io_r_246_b : _GEN_7835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7837 = 9'hf7 == r_count_25_io_out ? io_r_247_b : _GEN_7836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7838 = 9'hf8 == r_count_25_io_out ? io_r_248_b : _GEN_7837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7839 = 9'hf9 == r_count_25_io_out ? io_r_249_b : _GEN_7838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7840 = 9'hfa == r_count_25_io_out ? io_r_250_b : _GEN_7839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7841 = 9'hfb == r_count_25_io_out ? io_r_251_b : _GEN_7840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7842 = 9'hfc == r_count_25_io_out ? io_r_252_b : _GEN_7841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7843 = 9'hfd == r_count_25_io_out ? io_r_253_b : _GEN_7842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7844 = 9'hfe == r_count_25_io_out ? io_r_254_b : _GEN_7843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7845 = 9'hff == r_count_25_io_out ? io_r_255_b : _GEN_7844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7846 = 9'h100 == r_count_25_io_out ? io_r_256_b : _GEN_7845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7847 = 9'h101 == r_count_25_io_out ? io_r_257_b : _GEN_7846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7848 = 9'h102 == r_count_25_io_out ? io_r_258_b : _GEN_7847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7849 = 9'h103 == r_count_25_io_out ? io_r_259_b : _GEN_7848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7850 = 9'h104 == r_count_25_io_out ? io_r_260_b : _GEN_7849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7851 = 9'h105 == r_count_25_io_out ? io_r_261_b : _GEN_7850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7852 = 9'h106 == r_count_25_io_out ? io_r_262_b : _GEN_7851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7853 = 9'h107 == r_count_25_io_out ? io_r_263_b : _GEN_7852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7854 = 9'h108 == r_count_25_io_out ? io_r_264_b : _GEN_7853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7855 = 9'h109 == r_count_25_io_out ? io_r_265_b : _GEN_7854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7856 = 9'h10a == r_count_25_io_out ? io_r_266_b : _GEN_7855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7857 = 9'h10b == r_count_25_io_out ? io_r_267_b : _GEN_7856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7858 = 9'h10c == r_count_25_io_out ? io_r_268_b : _GEN_7857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7859 = 9'h10d == r_count_25_io_out ? io_r_269_b : _GEN_7858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7860 = 9'h10e == r_count_25_io_out ? io_r_270_b : _GEN_7859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7861 = 9'h10f == r_count_25_io_out ? io_r_271_b : _GEN_7860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7862 = 9'h110 == r_count_25_io_out ? io_r_272_b : _GEN_7861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7863 = 9'h111 == r_count_25_io_out ? io_r_273_b : _GEN_7862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7864 = 9'h112 == r_count_25_io_out ? io_r_274_b : _GEN_7863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7865 = 9'h113 == r_count_25_io_out ? io_r_275_b : _GEN_7864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7866 = 9'h114 == r_count_25_io_out ? io_r_276_b : _GEN_7865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7867 = 9'h115 == r_count_25_io_out ? io_r_277_b : _GEN_7866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7868 = 9'h116 == r_count_25_io_out ? io_r_278_b : _GEN_7867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7869 = 9'h117 == r_count_25_io_out ? io_r_279_b : _GEN_7868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7870 = 9'h118 == r_count_25_io_out ? io_r_280_b : _GEN_7869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7871 = 9'h119 == r_count_25_io_out ? io_r_281_b : _GEN_7870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7872 = 9'h11a == r_count_25_io_out ? io_r_282_b : _GEN_7871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7873 = 9'h11b == r_count_25_io_out ? io_r_283_b : _GEN_7872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7874 = 9'h11c == r_count_25_io_out ? io_r_284_b : _GEN_7873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7875 = 9'h11d == r_count_25_io_out ? io_r_285_b : _GEN_7874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7876 = 9'h11e == r_count_25_io_out ? io_r_286_b : _GEN_7875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7877 = 9'h11f == r_count_25_io_out ? io_r_287_b : _GEN_7876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7878 = 9'h120 == r_count_25_io_out ? io_r_288_b : _GEN_7877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7879 = 9'h121 == r_count_25_io_out ? io_r_289_b : _GEN_7878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7880 = 9'h122 == r_count_25_io_out ? io_r_290_b : _GEN_7879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7881 = 9'h123 == r_count_25_io_out ? io_r_291_b : _GEN_7880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7882 = 9'h124 == r_count_25_io_out ? io_r_292_b : _GEN_7881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7883 = 9'h125 == r_count_25_io_out ? io_r_293_b : _GEN_7882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7884 = 9'h126 == r_count_25_io_out ? io_r_294_b : _GEN_7883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7885 = 9'h127 == r_count_25_io_out ? io_r_295_b : _GEN_7884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7886 = 9'h128 == r_count_25_io_out ? io_r_296_b : _GEN_7885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7887 = 9'h129 == r_count_25_io_out ? io_r_297_b : _GEN_7886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7888 = 9'h12a == r_count_25_io_out ? io_r_298_b : _GEN_7887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7891 = 9'h1 == r_count_26_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7892 = 9'h2 == r_count_26_io_out ? io_r_2_b : _GEN_7891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7893 = 9'h3 == r_count_26_io_out ? io_r_3_b : _GEN_7892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7894 = 9'h4 == r_count_26_io_out ? io_r_4_b : _GEN_7893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7895 = 9'h5 == r_count_26_io_out ? io_r_5_b : _GEN_7894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7896 = 9'h6 == r_count_26_io_out ? io_r_6_b : _GEN_7895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7897 = 9'h7 == r_count_26_io_out ? io_r_7_b : _GEN_7896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7898 = 9'h8 == r_count_26_io_out ? io_r_8_b : _GEN_7897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7899 = 9'h9 == r_count_26_io_out ? io_r_9_b : _GEN_7898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7900 = 9'ha == r_count_26_io_out ? io_r_10_b : _GEN_7899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7901 = 9'hb == r_count_26_io_out ? io_r_11_b : _GEN_7900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7902 = 9'hc == r_count_26_io_out ? io_r_12_b : _GEN_7901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7903 = 9'hd == r_count_26_io_out ? io_r_13_b : _GEN_7902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7904 = 9'he == r_count_26_io_out ? io_r_14_b : _GEN_7903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7905 = 9'hf == r_count_26_io_out ? io_r_15_b : _GEN_7904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7906 = 9'h10 == r_count_26_io_out ? io_r_16_b : _GEN_7905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7907 = 9'h11 == r_count_26_io_out ? io_r_17_b : _GEN_7906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7908 = 9'h12 == r_count_26_io_out ? io_r_18_b : _GEN_7907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7909 = 9'h13 == r_count_26_io_out ? io_r_19_b : _GEN_7908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7910 = 9'h14 == r_count_26_io_out ? io_r_20_b : _GEN_7909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7911 = 9'h15 == r_count_26_io_out ? io_r_21_b : _GEN_7910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7912 = 9'h16 == r_count_26_io_out ? io_r_22_b : _GEN_7911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7913 = 9'h17 == r_count_26_io_out ? io_r_23_b : _GEN_7912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7914 = 9'h18 == r_count_26_io_out ? io_r_24_b : _GEN_7913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7915 = 9'h19 == r_count_26_io_out ? io_r_25_b : _GEN_7914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7916 = 9'h1a == r_count_26_io_out ? io_r_26_b : _GEN_7915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7917 = 9'h1b == r_count_26_io_out ? io_r_27_b : _GEN_7916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7918 = 9'h1c == r_count_26_io_out ? io_r_28_b : _GEN_7917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7919 = 9'h1d == r_count_26_io_out ? io_r_29_b : _GEN_7918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7920 = 9'h1e == r_count_26_io_out ? io_r_30_b : _GEN_7919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7921 = 9'h1f == r_count_26_io_out ? io_r_31_b : _GEN_7920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7922 = 9'h20 == r_count_26_io_out ? io_r_32_b : _GEN_7921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7923 = 9'h21 == r_count_26_io_out ? io_r_33_b : _GEN_7922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7924 = 9'h22 == r_count_26_io_out ? io_r_34_b : _GEN_7923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7925 = 9'h23 == r_count_26_io_out ? io_r_35_b : _GEN_7924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7926 = 9'h24 == r_count_26_io_out ? io_r_36_b : _GEN_7925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7927 = 9'h25 == r_count_26_io_out ? io_r_37_b : _GEN_7926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7928 = 9'h26 == r_count_26_io_out ? io_r_38_b : _GEN_7927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7929 = 9'h27 == r_count_26_io_out ? io_r_39_b : _GEN_7928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7930 = 9'h28 == r_count_26_io_out ? io_r_40_b : _GEN_7929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7931 = 9'h29 == r_count_26_io_out ? io_r_41_b : _GEN_7930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7932 = 9'h2a == r_count_26_io_out ? io_r_42_b : _GEN_7931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7933 = 9'h2b == r_count_26_io_out ? io_r_43_b : _GEN_7932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7934 = 9'h2c == r_count_26_io_out ? io_r_44_b : _GEN_7933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7935 = 9'h2d == r_count_26_io_out ? io_r_45_b : _GEN_7934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7936 = 9'h2e == r_count_26_io_out ? io_r_46_b : _GEN_7935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7937 = 9'h2f == r_count_26_io_out ? io_r_47_b : _GEN_7936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7938 = 9'h30 == r_count_26_io_out ? io_r_48_b : _GEN_7937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7939 = 9'h31 == r_count_26_io_out ? io_r_49_b : _GEN_7938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7940 = 9'h32 == r_count_26_io_out ? io_r_50_b : _GEN_7939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7941 = 9'h33 == r_count_26_io_out ? io_r_51_b : _GEN_7940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7942 = 9'h34 == r_count_26_io_out ? io_r_52_b : _GEN_7941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7943 = 9'h35 == r_count_26_io_out ? io_r_53_b : _GEN_7942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7944 = 9'h36 == r_count_26_io_out ? io_r_54_b : _GEN_7943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7945 = 9'h37 == r_count_26_io_out ? io_r_55_b : _GEN_7944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7946 = 9'h38 == r_count_26_io_out ? io_r_56_b : _GEN_7945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7947 = 9'h39 == r_count_26_io_out ? io_r_57_b : _GEN_7946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7948 = 9'h3a == r_count_26_io_out ? io_r_58_b : _GEN_7947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7949 = 9'h3b == r_count_26_io_out ? io_r_59_b : _GEN_7948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7950 = 9'h3c == r_count_26_io_out ? io_r_60_b : _GEN_7949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7951 = 9'h3d == r_count_26_io_out ? io_r_61_b : _GEN_7950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7952 = 9'h3e == r_count_26_io_out ? io_r_62_b : _GEN_7951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7953 = 9'h3f == r_count_26_io_out ? io_r_63_b : _GEN_7952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7954 = 9'h40 == r_count_26_io_out ? io_r_64_b : _GEN_7953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7955 = 9'h41 == r_count_26_io_out ? io_r_65_b : _GEN_7954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7956 = 9'h42 == r_count_26_io_out ? io_r_66_b : _GEN_7955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7957 = 9'h43 == r_count_26_io_out ? io_r_67_b : _GEN_7956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7958 = 9'h44 == r_count_26_io_out ? io_r_68_b : _GEN_7957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7959 = 9'h45 == r_count_26_io_out ? io_r_69_b : _GEN_7958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7960 = 9'h46 == r_count_26_io_out ? io_r_70_b : _GEN_7959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7961 = 9'h47 == r_count_26_io_out ? io_r_71_b : _GEN_7960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7962 = 9'h48 == r_count_26_io_out ? io_r_72_b : _GEN_7961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7963 = 9'h49 == r_count_26_io_out ? io_r_73_b : _GEN_7962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7964 = 9'h4a == r_count_26_io_out ? io_r_74_b : _GEN_7963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7965 = 9'h4b == r_count_26_io_out ? io_r_75_b : _GEN_7964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7966 = 9'h4c == r_count_26_io_out ? io_r_76_b : _GEN_7965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7967 = 9'h4d == r_count_26_io_out ? io_r_77_b : _GEN_7966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7968 = 9'h4e == r_count_26_io_out ? io_r_78_b : _GEN_7967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7969 = 9'h4f == r_count_26_io_out ? io_r_79_b : _GEN_7968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7970 = 9'h50 == r_count_26_io_out ? io_r_80_b : _GEN_7969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7971 = 9'h51 == r_count_26_io_out ? io_r_81_b : _GEN_7970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7972 = 9'h52 == r_count_26_io_out ? io_r_82_b : _GEN_7971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7973 = 9'h53 == r_count_26_io_out ? io_r_83_b : _GEN_7972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7974 = 9'h54 == r_count_26_io_out ? io_r_84_b : _GEN_7973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7975 = 9'h55 == r_count_26_io_out ? io_r_85_b : _GEN_7974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7976 = 9'h56 == r_count_26_io_out ? io_r_86_b : _GEN_7975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7977 = 9'h57 == r_count_26_io_out ? io_r_87_b : _GEN_7976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7978 = 9'h58 == r_count_26_io_out ? io_r_88_b : _GEN_7977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7979 = 9'h59 == r_count_26_io_out ? io_r_89_b : _GEN_7978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7980 = 9'h5a == r_count_26_io_out ? io_r_90_b : _GEN_7979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7981 = 9'h5b == r_count_26_io_out ? io_r_91_b : _GEN_7980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7982 = 9'h5c == r_count_26_io_out ? io_r_92_b : _GEN_7981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7983 = 9'h5d == r_count_26_io_out ? io_r_93_b : _GEN_7982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7984 = 9'h5e == r_count_26_io_out ? io_r_94_b : _GEN_7983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7985 = 9'h5f == r_count_26_io_out ? io_r_95_b : _GEN_7984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7986 = 9'h60 == r_count_26_io_out ? io_r_96_b : _GEN_7985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7987 = 9'h61 == r_count_26_io_out ? io_r_97_b : _GEN_7986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7988 = 9'h62 == r_count_26_io_out ? io_r_98_b : _GEN_7987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7989 = 9'h63 == r_count_26_io_out ? io_r_99_b : _GEN_7988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7990 = 9'h64 == r_count_26_io_out ? io_r_100_b : _GEN_7989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7991 = 9'h65 == r_count_26_io_out ? io_r_101_b : _GEN_7990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7992 = 9'h66 == r_count_26_io_out ? io_r_102_b : _GEN_7991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7993 = 9'h67 == r_count_26_io_out ? io_r_103_b : _GEN_7992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7994 = 9'h68 == r_count_26_io_out ? io_r_104_b : _GEN_7993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7995 = 9'h69 == r_count_26_io_out ? io_r_105_b : _GEN_7994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7996 = 9'h6a == r_count_26_io_out ? io_r_106_b : _GEN_7995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7997 = 9'h6b == r_count_26_io_out ? io_r_107_b : _GEN_7996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7998 = 9'h6c == r_count_26_io_out ? io_r_108_b : _GEN_7997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7999 = 9'h6d == r_count_26_io_out ? io_r_109_b : _GEN_7998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8000 = 9'h6e == r_count_26_io_out ? io_r_110_b : _GEN_7999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8001 = 9'h6f == r_count_26_io_out ? io_r_111_b : _GEN_8000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8002 = 9'h70 == r_count_26_io_out ? io_r_112_b : _GEN_8001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8003 = 9'h71 == r_count_26_io_out ? io_r_113_b : _GEN_8002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8004 = 9'h72 == r_count_26_io_out ? io_r_114_b : _GEN_8003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8005 = 9'h73 == r_count_26_io_out ? io_r_115_b : _GEN_8004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8006 = 9'h74 == r_count_26_io_out ? io_r_116_b : _GEN_8005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8007 = 9'h75 == r_count_26_io_out ? io_r_117_b : _GEN_8006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8008 = 9'h76 == r_count_26_io_out ? io_r_118_b : _GEN_8007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8009 = 9'h77 == r_count_26_io_out ? io_r_119_b : _GEN_8008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8010 = 9'h78 == r_count_26_io_out ? io_r_120_b : _GEN_8009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8011 = 9'h79 == r_count_26_io_out ? io_r_121_b : _GEN_8010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8012 = 9'h7a == r_count_26_io_out ? io_r_122_b : _GEN_8011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8013 = 9'h7b == r_count_26_io_out ? io_r_123_b : _GEN_8012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8014 = 9'h7c == r_count_26_io_out ? io_r_124_b : _GEN_8013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8015 = 9'h7d == r_count_26_io_out ? io_r_125_b : _GEN_8014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8016 = 9'h7e == r_count_26_io_out ? io_r_126_b : _GEN_8015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8017 = 9'h7f == r_count_26_io_out ? io_r_127_b : _GEN_8016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8018 = 9'h80 == r_count_26_io_out ? io_r_128_b : _GEN_8017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8019 = 9'h81 == r_count_26_io_out ? io_r_129_b : _GEN_8018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8020 = 9'h82 == r_count_26_io_out ? io_r_130_b : _GEN_8019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8021 = 9'h83 == r_count_26_io_out ? io_r_131_b : _GEN_8020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8022 = 9'h84 == r_count_26_io_out ? io_r_132_b : _GEN_8021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8023 = 9'h85 == r_count_26_io_out ? io_r_133_b : _GEN_8022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8024 = 9'h86 == r_count_26_io_out ? io_r_134_b : _GEN_8023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8025 = 9'h87 == r_count_26_io_out ? io_r_135_b : _GEN_8024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8026 = 9'h88 == r_count_26_io_out ? io_r_136_b : _GEN_8025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8027 = 9'h89 == r_count_26_io_out ? io_r_137_b : _GEN_8026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8028 = 9'h8a == r_count_26_io_out ? io_r_138_b : _GEN_8027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8029 = 9'h8b == r_count_26_io_out ? io_r_139_b : _GEN_8028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8030 = 9'h8c == r_count_26_io_out ? io_r_140_b : _GEN_8029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8031 = 9'h8d == r_count_26_io_out ? io_r_141_b : _GEN_8030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8032 = 9'h8e == r_count_26_io_out ? io_r_142_b : _GEN_8031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8033 = 9'h8f == r_count_26_io_out ? io_r_143_b : _GEN_8032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8034 = 9'h90 == r_count_26_io_out ? io_r_144_b : _GEN_8033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8035 = 9'h91 == r_count_26_io_out ? io_r_145_b : _GEN_8034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8036 = 9'h92 == r_count_26_io_out ? io_r_146_b : _GEN_8035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8037 = 9'h93 == r_count_26_io_out ? io_r_147_b : _GEN_8036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8038 = 9'h94 == r_count_26_io_out ? io_r_148_b : _GEN_8037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8039 = 9'h95 == r_count_26_io_out ? io_r_149_b : _GEN_8038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8040 = 9'h96 == r_count_26_io_out ? io_r_150_b : _GEN_8039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8041 = 9'h97 == r_count_26_io_out ? io_r_151_b : _GEN_8040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8042 = 9'h98 == r_count_26_io_out ? io_r_152_b : _GEN_8041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8043 = 9'h99 == r_count_26_io_out ? io_r_153_b : _GEN_8042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8044 = 9'h9a == r_count_26_io_out ? io_r_154_b : _GEN_8043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8045 = 9'h9b == r_count_26_io_out ? io_r_155_b : _GEN_8044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8046 = 9'h9c == r_count_26_io_out ? io_r_156_b : _GEN_8045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8047 = 9'h9d == r_count_26_io_out ? io_r_157_b : _GEN_8046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8048 = 9'h9e == r_count_26_io_out ? io_r_158_b : _GEN_8047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8049 = 9'h9f == r_count_26_io_out ? io_r_159_b : _GEN_8048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8050 = 9'ha0 == r_count_26_io_out ? io_r_160_b : _GEN_8049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8051 = 9'ha1 == r_count_26_io_out ? io_r_161_b : _GEN_8050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8052 = 9'ha2 == r_count_26_io_out ? io_r_162_b : _GEN_8051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8053 = 9'ha3 == r_count_26_io_out ? io_r_163_b : _GEN_8052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8054 = 9'ha4 == r_count_26_io_out ? io_r_164_b : _GEN_8053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8055 = 9'ha5 == r_count_26_io_out ? io_r_165_b : _GEN_8054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8056 = 9'ha6 == r_count_26_io_out ? io_r_166_b : _GEN_8055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8057 = 9'ha7 == r_count_26_io_out ? io_r_167_b : _GEN_8056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8058 = 9'ha8 == r_count_26_io_out ? io_r_168_b : _GEN_8057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8059 = 9'ha9 == r_count_26_io_out ? io_r_169_b : _GEN_8058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8060 = 9'haa == r_count_26_io_out ? io_r_170_b : _GEN_8059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8061 = 9'hab == r_count_26_io_out ? io_r_171_b : _GEN_8060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8062 = 9'hac == r_count_26_io_out ? io_r_172_b : _GEN_8061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8063 = 9'had == r_count_26_io_out ? io_r_173_b : _GEN_8062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8064 = 9'hae == r_count_26_io_out ? io_r_174_b : _GEN_8063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8065 = 9'haf == r_count_26_io_out ? io_r_175_b : _GEN_8064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8066 = 9'hb0 == r_count_26_io_out ? io_r_176_b : _GEN_8065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8067 = 9'hb1 == r_count_26_io_out ? io_r_177_b : _GEN_8066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8068 = 9'hb2 == r_count_26_io_out ? io_r_178_b : _GEN_8067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8069 = 9'hb3 == r_count_26_io_out ? io_r_179_b : _GEN_8068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8070 = 9'hb4 == r_count_26_io_out ? io_r_180_b : _GEN_8069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8071 = 9'hb5 == r_count_26_io_out ? io_r_181_b : _GEN_8070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8072 = 9'hb6 == r_count_26_io_out ? io_r_182_b : _GEN_8071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8073 = 9'hb7 == r_count_26_io_out ? io_r_183_b : _GEN_8072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8074 = 9'hb8 == r_count_26_io_out ? io_r_184_b : _GEN_8073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8075 = 9'hb9 == r_count_26_io_out ? io_r_185_b : _GEN_8074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8076 = 9'hba == r_count_26_io_out ? io_r_186_b : _GEN_8075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8077 = 9'hbb == r_count_26_io_out ? io_r_187_b : _GEN_8076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8078 = 9'hbc == r_count_26_io_out ? io_r_188_b : _GEN_8077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8079 = 9'hbd == r_count_26_io_out ? io_r_189_b : _GEN_8078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8080 = 9'hbe == r_count_26_io_out ? io_r_190_b : _GEN_8079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8081 = 9'hbf == r_count_26_io_out ? io_r_191_b : _GEN_8080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8082 = 9'hc0 == r_count_26_io_out ? io_r_192_b : _GEN_8081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8083 = 9'hc1 == r_count_26_io_out ? io_r_193_b : _GEN_8082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8084 = 9'hc2 == r_count_26_io_out ? io_r_194_b : _GEN_8083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8085 = 9'hc3 == r_count_26_io_out ? io_r_195_b : _GEN_8084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8086 = 9'hc4 == r_count_26_io_out ? io_r_196_b : _GEN_8085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8087 = 9'hc5 == r_count_26_io_out ? io_r_197_b : _GEN_8086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8088 = 9'hc6 == r_count_26_io_out ? io_r_198_b : _GEN_8087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8089 = 9'hc7 == r_count_26_io_out ? io_r_199_b : _GEN_8088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8090 = 9'hc8 == r_count_26_io_out ? io_r_200_b : _GEN_8089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8091 = 9'hc9 == r_count_26_io_out ? io_r_201_b : _GEN_8090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8092 = 9'hca == r_count_26_io_out ? io_r_202_b : _GEN_8091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8093 = 9'hcb == r_count_26_io_out ? io_r_203_b : _GEN_8092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8094 = 9'hcc == r_count_26_io_out ? io_r_204_b : _GEN_8093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8095 = 9'hcd == r_count_26_io_out ? io_r_205_b : _GEN_8094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8096 = 9'hce == r_count_26_io_out ? io_r_206_b : _GEN_8095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8097 = 9'hcf == r_count_26_io_out ? io_r_207_b : _GEN_8096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8098 = 9'hd0 == r_count_26_io_out ? io_r_208_b : _GEN_8097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8099 = 9'hd1 == r_count_26_io_out ? io_r_209_b : _GEN_8098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8100 = 9'hd2 == r_count_26_io_out ? io_r_210_b : _GEN_8099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8101 = 9'hd3 == r_count_26_io_out ? io_r_211_b : _GEN_8100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8102 = 9'hd4 == r_count_26_io_out ? io_r_212_b : _GEN_8101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8103 = 9'hd5 == r_count_26_io_out ? io_r_213_b : _GEN_8102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8104 = 9'hd6 == r_count_26_io_out ? io_r_214_b : _GEN_8103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8105 = 9'hd7 == r_count_26_io_out ? io_r_215_b : _GEN_8104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8106 = 9'hd8 == r_count_26_io_out ? io_r_216_b : _GEN_8105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8107 = 9'hd9 == r_count_26_io_out ? io_r_217_b : _GEN_8106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8108 = 9'hda == r_count_26_io_out ? io_r_218_b : _GEN_8107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8109 = 9'hdb == r_count_26_io_out ? io_r_219_b : _GEN_8108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8110 = 9'hdc == r_count_26_io_out ? io_r_220_b : _GEN_8109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8111 = 9'hdd == r_count_26_io_out ? io_r_221_b : _GEN_8110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8112 = 9'hde == r_count_26_io_out ? io_r_222_b : _GEN_8111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8113 = 9'hdf == r_count_26_io_out ? io_r_223_b : _GEN_8112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8114 = 9'he0 == r_count_26_io_out ? io_r_224_b : _GEN_8113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8115 = 9'he1 == r_count_26_io_out ? io_r_225_b : _GEN_8114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8116 = 9'he2 == r_count_26_io_out ? io_r_226_b : _GEN_8115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8117 = 9'he3 == r_count_26_io_out ? io_r_227_b : _GEN_8116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8118 = 9'he4 == r_count_26_io_out ? io_r_228_b : _GEN_8117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8119 = 9'he5 == r_count_26_io_out ? io_r_229_b : _GEN_8118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8120 = 9'he6 == r_count_26_io_out ? io_r_230_b : _GEN_8119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8121 = 9'he7 == r_count_26_io_out ? io_r_231_b : _GEN_8120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8122 = 9'he8 == r_count_26_io_out ? io_r_232_b : _GEN_8121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8123 = 9'he9 == r_count_26_io_out ? io_r_233_b : _GEN_8122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8124 = 9'hea == r_count_26_io_out ? io_r_234_b : _GEN_8123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8125 = 9'heb == r_count_26_io_out ? io_r_235_b : _GEN_8124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8126 = 9'hec == r_count_26_io_out ? io_r_236_b : _GEN_8125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8127 = 9'hed == r_count_26_io_out ? io_r_237_b : _GEN_8126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8128 = 9'hee == r_count_26_io_out ? io_r_238_b : _GEN_8127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8129 = 9'hef == r_count_26_io_out ? io_r_239_b : _GEN_8128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8130 = 9'hf0 == r_count_26_io_out ? io_r_240_b : _GEN_8129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8131 = 9'hf1 == r_count_26_io_out ? io_r_241_b : _GEN_8130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8132 = 9'hf2 == r_count_26_io_out ? io_r_242_b : _GEN_8131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8133 = 9'hf3 == r_count_26_io_out ? io_r_243_b : _GEN_8132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8134 = 9'hf4 == r_count_26_io_out ? io_r_244_b : _GEN_8133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8135 = 9'hf5 == r_count_26_io_out ? io_r_245_b : _GEN_8134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8136 = 9'hf6 == r_count_26_io_out ? io_r_246_b : _GEN_8135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8137 = 9'hf7 == r_count_26_io_out ? io_r_247_b : _GEN_8136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8138 = 9'hf8 == r_count_26_io_out ? io_r_248_b : _GEN_8137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8139 = 9'hf9 == r_count_26_io_out ? io_r_249_b : _GEN_8138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8140 = 9'hfa == r_count_26_io_out ? io_r_250_b : _GEN_8139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8141 = 9'hfb == r_count_26_io_out ? io_r_251_b : _GEN_8140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8142 = 9'hfc == r_count_26_io_out ? io_r_252_b : _GEN_8141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8143 = 9'hfd == r_count_26_io_out ? io_r_253_b : _GEN_8142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8144 = 9'hfe == r_count_26_io_out ? io_r_254_b : _GEN_8143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8145 = 9'hff == r_count_26_io_out ? io_r_255_b : _GEN_8144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8146 = 9'h100 == r_count_26_io_out ? io_r_256_b : _GEN_8145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8147 = 9'h101 == r_count_26_io_out ? io_r_257_b : _GEN_8146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8148 = 9'h102 == r_count_26_io_out ? io_r_258_b : _GEN_8147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8149 = 9'h103 == r_count_26_io_out ? io_r_259_b : _GEN_8148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8150 = 9'h104 == r_count_26_io_out ? io_r_260_b : _GEN_8149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8151 = 9'h105 == r_count_26_io_out ? io_r_261_b : _GEN_8150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8152 = 9'h106 == r_count_26_io_out ? io_r_262_b : _GEN_8151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8153 = 9'h107 == r_count_26_io_out ? io_r_263_b : _GEN_8152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8154 = 9'h108 == r_count_26_io_out ? io_r_264_b : _GEN_8153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8155 = 9'h109 == r_count_26_io_out ? io_r_265_b : _GEN_8154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8156 = 9'h10a == r_count_26_io_out ? io_r_266_b : _GEN_8155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8157 = 9'h10b == r_count_26_io_out ? io_r_267_b : _GEN_8156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8158 = 9'h10c == r_count_26_io_out ? io_r_268_b : _GEN_8157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8159 = 9'h10d == r_count_26_io_out ? io_r_269_b : _GEN_8158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8160 = 9'h10e == r_count_26_io_out ? io_r_270_b : _GEN_8159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8161 = 9'h10f == r_count_26_io_out ? io_r_271_b : _GEN_8160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8162 = 9'h110 == r_count_26_io_out ? io_r_272_b : _GEN_8161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8163 = 9'h111 == r_count_26_io_out ? io_r_273_b : _GEN_8162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8164 = 9'h112 == r_count_26_io_out ? io_r_274_b : _GEN_8163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8165 = 9'h113 == r_count_26_io_out ? io_r_275_b : _GEN_8164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8166 = 9'h114 == r_count_26_io_out ? io_r_276_b : _GEN_8165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8167 = 9'h115 == r_count_26_io_out ? io_r_277_b : _GEN_8166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8168 = 9'h116 == r_count_26_io_out ? io_r_278_b : _GEN_8167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8169 = 9'h117 == r_count_26_io_out ? io_r_279_b : _GEN_8168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8170 = 9'h118 == r_count_26_io_out ? io_r_280_b : _GEN_8169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8171 = 9'h119 == r_count_26_io_out ? io_r_281_b : _GEN_8170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8172 = 9'h11a == r_count_26_io_out ? io_r_282_b : _GEN_8171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8173 = 9'h11b == r_count_26_io_out ? io_r_283_b : _GEN_8172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8174 = 9'h11c == r_count_26_io_out ? io_r_284_b : _GEN_8173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8175 = 9'h11d == r_count_26_io_out ? io_r_285_b : _GEN_8174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8176 = 9'h11e == r_count_26_io_out ? io_r_286_b : _GEN_8175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8177 = 9'h11f == r_count_26_io_out ? io_r_287_b : _GEN_8176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8178 = 9'h120 == r_count_26_io_out ? io_r_288_b : _GEN_8177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8179 = 9'h121 == r_count_26_io_out ? io_r_289_b : _GEN_8178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8180 = 9'h122 == r_count_26_io_out ? io_r_290_b : _GEN_8179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8181 = 9'h123 == r_count_26_io_out ? io_r_291_b : _GEN_8180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8182 = 9'h124 == r_count_26_io_out ? io_r_292_b : _GEN_8181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8183 = 9'h125 == r_count_26_io_out ? io_r_293_b : _GEN_8182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8184 = 9'h126 == r_count_26_io_out ? io_r_294_b : _GEN_8183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8185 = 9'h127 == r_count_26_io_out ? io_r_295_b : _GEN_8184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8186 = 9'h128 == r_count_26_io_out ? io_r_296_b : _GEN_8185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8187 = 9'h129 == r_count_26_io_out ? io_r_297_b : _GEN_8186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8188 = 9'h12a == r_count_26_io_out ? io_r_298_b : _GEN_8187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8191 = 9'h1 == r_count_27_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8192 = 9'h2 == r_count_27_io_out ? io_r_2_b : _GEN_8191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8193 = 9'h3 == r_count_27_io_out ? io_r_3_b : _GEN_8192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8194 = 9'h4 == r_count_27_io_out ? io_r_4_b : _GEN_8193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8195 = 9'h5 == r_count_27_io_out ? io_r_5_b : _GEN_8194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8196 = 9'h6 == r_count_27_io_out ? io_r_6_b : _GEN_8195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8197 = 9'h7 == r_count_27_io_out ? io_r_7_b : _GEN_8196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8198 = 9'h8 == r_count_27_io_out ? io_r_8_b : _GEN_8197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8199 = 9'h9 == r_count_27_io_out ? io_r_9_b : _GEN_8198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8200 = 9'ha == r_count_27_io_out ? io_r_10_b : _GEN_8199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8201 = 9'hb == r_count_27_io_out ? io_r_11_b : _GEN_8200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8202 = 9'hc == r_count_27_io_out ? io_r_12_b : _GEN_8201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8203 = 9'hd == r_count_27_io_out ? io_r_13_b : _GEN_8202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8204 = 9'he == r_count_27_io_out ? io_r_14_b : _GEN_8203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8205 = 9'hf == r_count_27_io_out ? io_r_15_b : _GEN_8204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8206 = 9'h10 == r_count_27_io_out ? io_r_16_b : _GEN_8205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8207 = 9'h11 == r_count_27_io_out ? io_r_17_b : _GEN_8206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8208 = 9'h12 == r_count_27_io_out ? io_r_18_b : _GEN_8207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8209 = 9'h13 == r_count_27_io_out ? io_r_19_b : _GEN_8208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8210 = 9'h14 == r_count_27_io_out ? io_r_20_b : _GEN_8209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8211 = 9'h15 == r_count_27_io_out ? io_r_21_b : _GEN_8210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8212 = 9'h16 == r_count_27_io_out ? io_r_22_b : _GEN_8211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8213 = 9'h17 == r_count_27_io_out ? io_r_23_b : _GEN_8212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8214 = 9'h18 == r_count_27_io_out ? io_r_24_b : _GEN_8213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8215 = 9'h19 == r_count_27_io_out ? io_r_25_b : _GEN_8214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8216 = 9'h1a == r_count_27_io_out ? io_r_26_b : _GEN_8215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8217 = 9'h1b == r_count_27_io_out ? io_r_27_b : _GEN_8216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8218 = 9'h1c == r_count_27_io_out ? io_r_28_b : _GEN_8217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8219 = 9'h1d == r_count_27_io_out ? io_r_29_b : _GEN_8218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8220 = 9'h1e == r_count_27_io_out ? io_r_30_b : _GEN_8219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8221 = 9'h1f == r_count_27_io_out ? io_r_31_b : _GEN_8220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8222 = 9'h20 == r_count_27_io_out ? io_r_32_b : _GEN_8221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8223 = 9'h21 == r_count_27_io_out ? io_r_33_b : _GEN_8222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8224 = 9'h22 == r_count_27_io_out ? io_r_34_b : _GEN_8223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8225 = 9'h23 == r_count_27_io_out ? io_r_35_b : _GEN_8224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8226 = 9'h24 == r_count_27_io_out ? io_r_36_b : _GEN_8225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8227 = 9'h25 == r_count_27_io_out ? io_r_37_b : _GEN_8226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8228 = 9'h26 == r_count_27_io_out ? io_r_38_b : _GEN_8227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8229 = 9'h27 == r_count_27_io_out ? io_r_39_b : _GEN_8228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8230 = 9'h28 == r_count_27_io_out ? io_r_40_b : _GEN_8229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8231 = 9'h29 == r_count_27_io_out ? io_r_41_b : _GEN_8230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8232 = 9'h2a == r_count_27_io_out ? io_r_42_b : _GEN_8231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8233 = 9'h2b == r_count_27_io_out ? io_r_43_b : _GEN_8232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8234 = 9'h2c == r_count_27_io_out ? io_r_44_b : _GEN_8233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8235 = 9'h2d == r_count_27_io_out ? io_r_45_b : _GEN_8234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8236 = 9'h2e == r_count_27_io_out ? io_r_46_b : _GEN_8235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8237 = 9'h2f == r_count_27_io_out ? io_r_47_b : _GEN_8236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8238 = 9'h30 == r_count_27_io_out ? io_r_48_b : _GEN_8237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8239 = 9'h31 == r_count_27_io_out ? io_r_49_b : _GEN_8238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8240 = 9'h32 == r_count_27_io_out ? io_r_50_b : _GEN_8239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8241 = 9'h33 == r_count_27_io_out ? io_r_51_b : _GEN_8240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8242 = 9'h34 == r_count_27_io_out ? io_r_52_b : _GEN_8241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8243 = 9'h35 == r_count_27_io_out ? io_r_53_b : _GEN_8242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8244 = 9'h36 == r_count_27_io_out ? io_r_54_b : _GEN_8243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8245 = 9'h37 == r_count_27_io_out ? io_r_55_b : _GEN_8244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8246 = 9'h38 == r_count_27_io_out ? io_r_56_b : _GEN_8245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8247 = 9'h39 == r_count_27_io_out ? io_r_57_b : _GEN_8246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8248 = 9'h3a == r_count_27_io_out ? io_r_58_b : _GEN_8247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8249 = 9'h3b == r_count_27_io_out ? io_r_59_b : _GEN_8248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8250 = 9'h3c == r_count_27_io_out ? io_r_60_b : _GEN_8249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8251 = 9'h3d == r_count_27_io_out ? io_r_61_b : _GEN_8250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8252 = 9'h3e == r_count_27_io_out ? io_r_62_b : _GEN_8251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8253 = 9'h3f == r_count_27_io_out ? io_r_63_b : _GEN_8252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8254 = 9'h40 == r_count_27_io_out ? io_r_64_b : _GEN_8253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8255 = 9'h41 == r_count_27_io_out ? io_r_65_b : _GEN_8254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8256 = 9'h42 == r_count_27_io_out ? io_r_66_b : _GEN_8255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8257 = 9'h43 == r_count_27_io_out ? io_r_67_b : _GEN_8256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8258 = 9'h44 == r_count_27_io_out ? io_r_68_b : _GEN_8257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8259 = 9'h45 == r_count_27_io_out ? io_r_69_b : _GEN_8258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8260 = 9'h46 == r_count_27_io_out ? io_r_70_b : _GEN_8259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8261 = 9'h47 == r_count_27_io_out ? io_r_71_b : _GEN_8260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8262 = 9'h48 == r_count_27_io_out ? io_r_72_b : _GEN_8261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8263 = 9'h49 == r_count_27_io_out ? io_r_73_b : _GEN_8262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8264 = 9'h4a == r_count_27_io_out ? io_r_74_b : _GEN_8263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8265 = 9'h4b == r_count_27_io_out ? io_r_75_b : _GEN_8264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8266 = 9'h4c == r_count_27_io_out ? io_r_76_b : _GEN_8265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8267 = 9'h4d == r_count_27_io_out ? io_r_77_b : _GEN_8266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8268 = 9'h4e == r_count_27_io_out ? io_r_78_b : _GEN_8267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8269 = 9'h4f == r_count_27_io_out ? io_r_79_b : _GEN_8268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8270 = 9'h50 == r_count_27_io_out ? io_r_80_b : _GEN_8269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8271 = 9'h51 == r_count_27_io_out ? io_r_81_b : _GEN_8270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8272 = 9'h52 == r_count_27_io_out ? io_r_82_b : _GEN_8271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8273 = 9'h53 == r_count_27_io_out ? io_r_83_b : _GEN_8272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8274 = 9'h54 == r_count_27_io_out ? io_r_84_b : _GEN_8273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8275 = 9'h55 == r_count_27_io_out ? io_r_85_b : _GEN_8274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8276 = 9'h56 == r_count_27_io_out ? io_r_86_b : _GEN_8275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8277 = 9'h57 == r_count_27_io_out ? io_r_87_b : _GEN_8276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8278 = 9'h58 == r_count_27_io_out ? io_r_88_b : _GEN_8277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8279 = 9'h59 == r_count_27_io_out ? io_r_89_b : _GEN_8278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8280 = 9'h5a == r_count_27_io_out ? io_r_90_b : _GEN_8279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8281 = 9'h5b == r_count_27_io_out ? io_r_91_b : _GEN_8280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8282 = 9'h5c == r_count_27_io_out ? io_r_92_b : _GEN_8281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8283 = 9'h5d == r_count_27_io_out ? io_r_93_b : _GEN_8282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8284 = 9'h5e == r_count_27_io_out ? io_r_94_b : _GEN_8283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8285 = 9'h5f == r_count_27_io_out ? io_r_95_b : _GEN_8284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8286 = 9'h60 == r_count_27_io_out ? io_r_96_b : _GEN_8285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8287 = 9'h61 == r_count_27_io_out ? io_r_97_b : _GEN_8286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8288 = 9'h62 == r_count_27_io_out ? io_r_98_b : _GEN_8287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8289 = 9'h63 == r_count_27_io_out ? io_r_99_b : _GEN_8288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8290 = 9'h64 == r_count_27_io_out ? io_r_100_b : _GEN_8289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8291 = 9'h65 == r_count_27_io_out ? io_r_101_b : _GEN_8290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8292 = 9'h66 == r_count_27_io_out ? io_r_102_b : _GEN_8291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8293 = 9'h67 == r_count_27_io_out ? io_r_103_b : _GEN_8292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8294 = 9'h68 == r_count_27_io_out ? io_r_104_b : _GEN_8293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8295 = 9'h69 == r_count_27_io_out ? io_r_105_b : _GEN_8294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8296 = 9'h6a == r_count_27_io_out ? io_r_106_b : _GEN_8295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8297 = 9'h6b == r_count_27_io_out ? io_r_107_b : _GEN_8296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8298 = 9'h6c == r_count_27_io_out ? io_r_108_b : _GEN_8297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8299 = 9'h6d == r_count_27_io_out ? io_r_109_b : _GEN_8298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8300 = 9'h6e == r_count_27_io_out ? io_r_110_b : _GEN_8299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8301 = 9'h6f == r_count_27_io_out ? io_r_111_b : _GEN_8300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8302 = 9'h70 == r_count_27_io_out ? io_r_112_b : _GEN_8301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8303 = 9'h71 == r_count_27_io_out ? io_r_113_b : _GEN_8302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8304 = 9'h72 == r_count_27_io_out ? io_r_114_b : _GEN_8303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8305 = 9'h73 == r_count_27_io_out ? io_r_115_b : _GEN_8304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8306 = 9'h74 == r_count_27_io_out ? io_r_116_b : _GEN_8305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8307 = 9'h75 == r_count_27_io_out ? io_r_117_b : _GEN_8306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8308 = 9'h76 == r_count_27_io_out ? io_r_118_b : _GEN_8307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8309 = 9'h77 == r_count_27_io_out ? io_r_119_b : _GEN_8308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8310 = 9'h78 == r_count_27_io_out ? io_r_120_b : _GEN_8309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8311 = 9'h79 == r_count_27_io_out ? io_r_121_b : _GEN_8310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8312 = 9'h7a == r_count_27_io_out ? io_r_122_b : _GEN_8311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8313 = 9'h7b == r_count_27_io_out ? io_r_123_b : _GEN_8312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8314 = 9'h7c == r_count_27_io_out ? io_r_124_b : _GEN_8313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8315 = 9'h7d == r_count_27_io_out ? io_r_125_b : _GEN_8314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8316 = 9'h7e == r_count_27_io_out ? io_r_126_b : _GEN_8315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8317 = 9'h7f == r_count_27_io_out ? io_r_127_b : _GEN_8316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8318 = 9'h80 == r_count_27_io_out ? io_r_128_b : _GEN_8317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8319 = 9'h81 == r_count_27_io_out ? io_r_129_b : _GEN_8318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8320 = 9'h82 == r_count_27_io_out ? io_r_130_b : _GEN_8319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8321 = 9'h83 == r_count_27_io_out ? io_r_131_b : _GEN_8320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8322 = 9'h84 == r_count_27_io_out ? io_r_132_b : _GEN_8321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8323 = 9'h85 == r_count_27_io_out ? io_r_133_b : _GEN_8322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8324 = 9'h86 == r_count_27_io_out ? io_r_134_b : _GEN_8323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8325 = 9'h87 == r_count_27_io_out ? io_r_135_b : _GEN_8324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8326 = 9'h88 == r_count_27_io_out ? io_r_136_b : _GEN_8325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8327 = 9'h89 == r_count_27_io_out ? io_r_137_b : _GEN_8326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8328 = 9'h8a == r_count_27_io_out ? io_r_138_b : _GEN_8327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8329 = 9'h8b == r_count_27_io_out ? io_r_139_b : _GEN_8328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8330 = 9'h8c == r_count_27_io_out ? io_r_140_b : _GEN_8329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8331 = 9'h8d == r_count_27_io_out ? io_r_141_b : _GEN_8330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8332 = 9'h8e == r_count_27_io_out ? io_r_142_b : _GEN_8331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8333 = 9'h8f == r_count_27_io_out ? io_r_143_b : _GEN_8332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8334 = 9'h90 == r_count_27_io_out ? io_r_144_b : _GEN_8333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8335 = 9'h91 == r_count_27_io_out ? io_r_145_b : _GEN_8334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8336 = 9'h92 == r_count_27_io_out ? io_r_146_b : _GEN_8335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8337 = 9'h93 == r_count_27_io_out ? io_r_147_b : _GEN_8336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8338 = 9'h94 == r_count_27_io_out ? io_r_148_b : _GEN_8337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8339 = 9'h95 == r_count_27_io_out ? io_r_149_b : _GEN_8338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8340 = 9'h96 == r_count_27_io_out ? io_r_150_b : _GEN_8339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8341 = 9'h97 == r_count_27_io_out ? io_r_151_b : _GEN_8340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8342 = 9'h98 == r_count_27_io_out ? io_r_152_b : _GEN_8341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8343 = 9'h99 == r_count_27_io_out ? io_r_153_b : _GEN_8342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8344 = 9'h9a == r_count_27_io_out ? io_r_154_b : _GEN_8343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8345 = 9'h9b == r_count_27_io_out ? io_r_155_b : _GEN_8344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8346 = 9'h9c == r_count_27_io_out ? io_r_156_b : _GEN_8345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8347 = 9'h9d == r_count_27_io_out ? io_r_157_b : _GEN_8346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8348 = 9'h9e == r_count_27_io_out ? io_r_158_b : _GEN_8347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8349 = 9'h9f == r_count_27_io_out ? io_r_159_b : _GEN_8348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8350 = 9'ha0 == r_count_27_io_out ? io_r_160_b : _GEN_8349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8351 = 9'ha1 == r_count_27_io_out ? io_r_161_b : _GEN_8350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8352 = 9'ha2 == r_count_27_io_out ? io_r_162_b : _GEN_8351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8353 = 9'ha3 == r_count_27_io_out ? io_r_163_b : _GEN_8352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8354 = 9'ha4 == r_count_27_io_out ? io_r_164_b : _GEN_8353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8355 = 9'ha5 == r_count_27_io_out ? io_r_165_b : _GEN_8354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8356 = 9'ha6 == r_count_27_io_out ? io_r_166_b : _GEN_8355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8357 = 9'ha7 == r_count_27_io_out ? io_r_167_b : _GEN_8356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8358 = 9'ha8 == r_count_27_io_out ? io_r_168_b : _GEN_8357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8359 = 9'ha9 == r_count_27_io_out ? io_r_169_b : _GEN_8358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8360 = 9'haa == r_count_27_io_out ? io_r_170_b : _GEN_8359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8361 = 9'hab == r_count_27_io_out ? io_r_171_b : _GEN_8360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8362 = 9'hac == r_count_27_io_out ? io_r_172_b : _GEN_8361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8363 = 9'had == r_count_27_io_out ? io_r_173_b : _GEN_8362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8364 = 9'hae == r_count_27_io_out ? io_r_174_b : _GEN_8363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8365 = 9'haf == r_count_27_io_out ? io_r_175_b : _GEN_8364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8366 = 9'hb0 == r_count_27_io_out ? io_r_176_b : _GEN_8365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8367 = 9'hb1 == r_count_27_io_out ? io_r_177_b : _GEN_8366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8368 = 9'hb2 == r_count_27_io_out ? io_r_178_b : _GEN_8367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8369 = 9'hb3 == r_count_27_io_out ? io_r_179_b : _GEN_8368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8370 = 9'hb4 == r_count_27_io_out ? io_r_180_b : _GEN_8369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8371 = 9'hb5 == r_count_27_io_out ? io_r_181_b : _GEN_8370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8372 = 9'hb6 == r_count_27_io_out ? io_r_182_b : _GEN_8371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8373 = 9'hb7 == r_count_27_io_out ? io_r_183_b : _GEN_8372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8374 = 9'hb8 == r_count_27_io_out ? io_r_184_b : _GEN_8373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8375 = 9'hb9 == r_count_27_io_out ? io_r_185_b : _GEN_8374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8376 = 9'hba == r_count_27_io_out ? io_r_186_b : _GEN_8375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8377 = 9'hbb == r_count_27_io_out ? io_r_187_b : _GEN_8376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8378 = 9'hbc == r_count_27_io_out ? io_r_188_b : _GEN_8377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8379 = 9'hbd == r_count_27_io_out ? io_r_189_b : _GEN_8378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8380 = 9'hbe == r_count_27_io_out ? io_r_190_b : _GEN_8379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8381 = 9'hbf == r_count_27_io_out ? io_r_191_b : _GEN_8380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8382 = 9'hc0 == r_count_27_io_out ? io_r_192_b : _GEN_8381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8383 = 9'hc1 == r_count_27_io_out ? io_r_193_b : _GEN_8382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8384 = 9'hc2 == r_count_27_io_out ? io_r_194_b : _GEN_8383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8385 = 9'hc3 == r_count_27_io_out ? io_r_195_b : _GEN_8384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8386 = 9'hc4 == r_count_27_io_out ? io_r_196_b : _GEN_8385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8387 = 9'hc5 == r_count_27_io_out ? io_r_197_b : _GEN_8386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8388 = 9'hc6 == r_count_27_io_out ? io_r_198_b : _GEN_8387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8389 = 9'hc7 == r_count_27_io_out ? io_r_199_b : _GEN_8388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8390 = 9'hc8 == r_count_27_io_out ? io_r_200_b : _GEN_8389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8391 = 9'hc9 == r_count_27_io_out ? io_r_201_b : _GEN_8390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8392 = 9'hca == r_count_27_io_out ? io_r_202_b : _GEN_8391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8393 = 9'hcb == r_count_27_io_out ? io_r_203_b : _GEN_8392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8394 = 9'hcc == r_count_27_io_out ? io_r_204_b : _GEN_8393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8395 = 9'hcd == r_count_27_io_out ? io_r_205_b : _GEN_8394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8396 = 9'hce == r_count_27_io_out ? io_r_206_b : _GEN_8395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8397 = 9'hcf == r_count_27_io_out ? io_r_207_b : _GEN_8396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8398 = 9'hd0 == r_count_27_io_out ? io_r_208_b : _GEN_8397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8399 = 9'hd1 == r_count_27_io_out ? io_r_209_b : _GEN_8398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8400 = 9'hd2 == r_count_27_io_out ? io_r_210_b : _GEN_8399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8401 = 9'hd3 == r_count_27_io_out ? io_r_211_b : _GEN_8400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8402 = 9'hd4 == r_count_27_io_out ? io_r_212_b : _GEN_8401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8403 = 9'hd5 == r_count_27_io_out ? io_r_213_b : _GEN_8402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8404 = 9'hd6 == r_count_27_io_out ? io_r_214_b : _GEN_8403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8405 = 9'hd7 == r_count_27_io_out ? io_r_215_b : _GEN_8404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8406 = 9'hd8 == r_count_27_io_out ? io_r_216_b : _GEN_8405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8407 = 9'hd9 == r_count_27_io_out ? io_r_217_b : _GEN_8406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8408 = 9'hda == r_count_27_io_out ? io_r_218_b : _GEN_8407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8409 = 9'hdb == r_count_27_io_out ? io_r_219_b : _GEN_8408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8410 = 9'hdc == r_count_27_io_out ? io_r_220_b : _GEN_8409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8411 = 9'hdd == r_count_27_io_out ? io_r_221_b : _GEN_8410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8412 = 9'hde == r_count_27_io_out ? io_r_222_b : _GEN_8411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8413 = 9'hdf == r_count_27_io_out ? io_r_223_b : _GEN_8412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8414 = 9'he0 == r_count_27_io_out ? io_r_224_b : _GEN_8413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8415 = 9'he1 == r_count_27_io_out ? io_r_225_b : _GEN_8414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8416 = 9'he2 == r_count_27_io_out ? io_r_226_b : _GEN_8415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8417 = 9'he3 == r_count_27_io_out ? io_r_227_b : _GEN_8416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8418 = 9'he4 == r_count_27_io_out ? io_r_228_b : _GEN_8417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8419 = 9'he5 == r_count_27_io_out ? io_r_229_b : _GEN_8418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8420 = 9'he6 == r_count_27_io_out ? io_r_230_b : _GEN_8419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8421 = 9'he7 == r_count_27_io_out ? io_r_231_b : _GEN_8420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8422 = 9'he8 == r_count_27_io_out ? io_r_232_b : _GEN_8421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8423 = 9'he9 == r_count_27_io_out ? io_r_233_b : _GEN_8422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8424 = 9'hea == r_count_27_io_out ? io_r_234_b : _GEN_8423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8425 = 9'heb == r_count_27_io_out ? io_r_235_b : _GEN_8424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8426 = 9'hec == r_count_27_io_out ? io_r_236_b : _GEN_8425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8427 = 9'hed == r_count_27_io_out ? io_r_237_b : _GEN_8426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8428 = 9'hee == r_count_27_io_out ? io_r_238_b : _GEN_8427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8429 = 9'hef == r_count_27_io_out ? io_r_239_b : _GEN_8428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8430 = 9'hf0 == r_count_27_io_out ? io_r_240_b : _GEN_8429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8431 = 9'hf1 == r_count_27_io_out ? io_r_241_b : _GEN_8430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8432 = 9'hf2 == r_count_27_io_out ? io_r_242_b : _GEN_8431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8433 = 9'hf3 == r_count_27_io_out ? io_r_243_b : _GEN_8432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8434 = 9'hf4 == r_count_27_io_out ? io_r_244_b : _GEN_8433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8435 = 9'hf5 == r_count_27_io_out ? io_r_245_b : _GEN_8434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8436 = 9'hf6 == r_count_27_io_out ? io_r_246_b : _GEN_8435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8437 = 9'hf7 == r_count_27_io_out ? io_r_247_b : _GEN_8436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8438 = 9'hf8 == r_count_27_io_out ? io_r_248_b : _GEN_8437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8439 = 9'hf9 == r_count_27_io_out ? io_r_249_b : _GEN_8438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8440 = 9'hfa == r_count_27_io_out ? io_r_250_b : _GEN_8439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8441 = 9'hfb == r_count_27_io_out ? io_r_251_b : _GEN_8440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8442 = 9'hfc == r_count_27_io_out ? io_r_252_b : _GEN_8441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8443 = 9'hfd == r_count_27_io_out ? io_r_253_b : _GEN_8442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8444 = 9'hfe == r_count_27_io_out ? io_r_254_b : _GEN_8443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8445 = 9'hff == r_count_27_io_out ? io_r_255_b : _GEN_8444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8446 = 9'h100 == r_count_27_io_out ? io_r_256_b : _GEN_8445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8447 = 9'h101 == r_count_27_io_out ? io_r_257_b : _GEN_8446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8448 = 9'h102 == r_count_27_io_out ? io_r_258_b : _GEN_8447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8449 = 9'h103 == r_count_27_io_out ? io_r_259_b : _GEN_8448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8450 = 9'h104 == r_count_27_io_out ? io_r_260_b : _GEN_8449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8451 = 9'h105 == r_count_27_io_out ? io_r_261_b : _GEN_8450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8452 = 9'h106 == r_count_27_io_out ? io_r_262_b : _GEN_8451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8453 = 9'h107 == r_count_27_io_out ? io_r_263_b : _GEN_8452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8454 = 9'h108 == r_count_27_io_out ? io_r_264_b : _GEN_8453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8455 = 9'h109 == r_count_27_io_out ? io_r_265_b : _GEN_8454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8456 = 9'h10a == r_count_27_io_out ? io_r_266_b : _GEN_8455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8457 = 9'h10b == r_count_27_io_out ? io_r_267_b : _GEN_8456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8458 = 9'h10c == r_count_27_io_out ? io_r_268_b : _GEN_8457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8459 = 9'h10d == r_count_27_io_out ? io_r_269_b : _GEN_8458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8460 = 9'h10e == r_count_27_io_out ? io_r_270_b : _GEN_8459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8461 = 9'h10f == r_count_27_io_out ? io_r_271_b : _GEN_8460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8462 = 9'h110 == r_count_27_io_out ? io_r_272_b : _GEN_8461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8463 = 9'h111 == r_count_27_io_out ? io_r_273_b : _GEN_8462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8464 = 9'h112 == r_count_27_io_out ? io_r_274_b : _GEN_8463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8465 = 9'h113 == r_count_27_io_out ? io_r_275_b : _GEN_8464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8466 = 9'h114 == r_count_27_io_out ? io_r_276_b : _GEN_8465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8467 = 9'h115 == r_count_27_io_out ? io_r_277_b : _GEN_8466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8468 = 9'h116 == r_count_27_io_out ? io_r_278_b : _GEN_8467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8469 = 9'h117 == r_count_27_io_out ? io_r_279_b : _GEN_8468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8470 = 9'h118 == r_count_27_io_out ? io_r_280_b : _GEN_8469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8471 = 9'h119 == r_count_27_io_out ? io_r_281_b : _GEN_8470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8472 = 9'h11a == r_count_27_io_out ? io_r_282_b : _GEN_8471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8473 = 9'h11b == r_count_27_io_out ? io_r_283_b : _GEN_8472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8474 = 9'h11c == r_count_27_io_out ? io_r_284_b : _GEN_8473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8475 = 9'h11d == r_count_27_io_out ? io_r_285_b : _GEN_8474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8476 = 9'h11e == r_count_27_io_out ? io_r_286_b : _GEN_8475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8477 = 9'h11f == r_count_27_io_out ? io_r_287_b : _GEN_8476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8478 = 9'h120 == r_count_27_io_out ? io_r_288_b : _GEN_8477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8479 = 9'h121 == r_count_27_io_out ? io_r_289_b : _GEN_8478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8480 = 9'h122 == r_count_27_io_out ? io_r_290_b : _GEN_8479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8481 = 9'h123 == r_count_27_io_out ? io_r_291_b : _GEN_8480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8482 = 9'h124 == r_count_27_io_out ? io_r_292_b : _GEN_8481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8483 = 9'h125 == r_count_27_io_out ? io_r_293_b : _GEN_8482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8484 = 9'h126 == r_count_27_io_out ? io_r_294_b : _GEN_8483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8485 = 9'h127 == r_count_27_io_out ? io_r_295_b : _GEN_8484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8486 = 9'h128 == r_count_27_io_out ? io_r_296_b : _GEN_8485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8487 = 9'h129 == r_count_27_io_out ? io_r_297_b : _GEN_8486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8488 = 9'h12a == r_count_27_io_out ? io_r_298_b : _GEN_8487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8491 = 9'h1 == r_count_28_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8492 = 9'h2 == r_count_28_io_out ? io_r_2_b : _GEN_8491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8493 = 9'h3 == r_count_28_io_out ? io_r_3_b : _GEN_8492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8494 = 9'h4 == r_count_28_io_out ? io_r_4_b : _GEN_8493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8495 = 9'h5 == r_count_28_io_out ? io_r_5_b : _GEN_8494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8496 = 9'h6 == r_count_28_io_out ? io_r_6_b : _GEN_8495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8497 = 9'h7 == r_count_28_io_out ? io_r_7_b : _GEN_8496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8498 = 9'h8 == r_count_28_io_out ? io_r_8_b : _GEN_8497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8499 = 9'h9 == r_count_28_io_out ? io_r_9_b : _GEN_8498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8500 = 9'ha == r_count_28_io_out ? io_r_10_b : _GEN_8499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8501 = 9'hb == r_count_28_io_out ? io_r_11_b : _GEN_8500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8502 = 9'hc == r_count_28_io_out ? io_r_12_b : _GEN_8501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8503 = 9'hd == r_count_28_io_out ? io_r_13_b : _GEN_8502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8504 = 9'he == r_count_28_io_out ? io_r_14_b : _GEN_8503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8505 = 9'hf == r_count_28_io_out ? io_r_15_b : _GEN_8504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8506 = 9'h10 == r_count_28_io_out ? io_r_16_b : _GEN_8505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8507 = 9'h11 == r_count_28_io_out ? io_r_17_b : _GEN_8506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8508 = 9'h12 == r_count_28_io_out ? io_r_18_b : _GEN_8507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8509 = 9'h13 == r_count_28_io_out ? io_r_19_b : _GEN_8508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8510 = 9'h14 == r_count_28_io_out ? io_r_20_b : _GEN_8509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8511 = 9'h15 == r_count_28_io_out ? io_r_21_b : _GEN_8510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8512 = 9'h16 == r_count_28_io_out ? io_r_22_b : _GEN_8511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8513 = 9'h17 == r_count_28_io_out ? io_r_23_b : _GEN_8512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8514 = 9'h18 == r_count_28_io_out ? io_r_24_b : _GEN_8513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8515 = 9'h19 == r_count_28_io_out ? io_r_25_b : _GEN_8514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8516 = 9'h1a == r_count_28_io_out ? io_r_26_b : _GEN_8515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8517 = 9'h1b == r_count_28_io_out ? io_r_27_b : _GEN_8516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8518 = 9'h1c == r_count_28_io_out ? io_r_28_b : _GEN_8517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8519 = 9'h1d == r_count_28_io_out ? io_r_29_b : _GEN_8518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8520 = 9'h1e == r_count_28_io_out ? io_r_30_b : _GEN_8519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8521 = 9'h1f == r_count_28_io_out ? io_r_31_b : _GEN_8520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8522 = 9'h20 == r_count_28_io_out ? io_r_32_b : _GEN_8521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8523 = 9'h21 == r_count_28_io_out ? io_r_33_b : _GEN_8522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8524 = 9'h22 == r_count_28_io_out ? io_r_34_b : _GEN_8523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8525 = 9'h23 == r_count_28_io_out ? io_r_35_b : _GEN_8524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8526 = 9'h24 == r_count_28_io_out ? io_r_36_b : _GEN_8525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8527 = 9'h25 == r_count_28_io_out ? io_r_37_b : _GEN_8526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8528 = 9'h26 == r_count_28_io_out ? io_r_38_b : _GEN_8527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8529 = 9'h27 == r_count_28_io_out ? io_r_39_b : _GEN_8528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8530 = 9'h28 == r_count_28_io_out ? io_r_40_b : _GEN_8529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8531 = 9'h29 == r_count_28_io_out ? io_r_41_b : _GEN_8530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8532 = 9'h2a == r_count_28_io_out ? io_r_42_b : _GEN_8531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8533 = 9'h2b == r_count_28_io_out ? io_r_43_b : _GEN_8532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8534 = 9'h2c == r_count_28_io_out ? io_r_44_b : _GEN_8533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8535 = 9'h2d == r_count_28_io_out ? io_r_45_b : _GEN_8534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8536 = 9'h2e == r_count_28_io_out ? io_r_46_b : _GEN_8535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8537 = 9'h2f == r_count_28_io_out ? io_r_47_b : _GEN_8536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8538 = 9'h30 == r_count_28_io_out ? io_r_48_b : _GEN_8537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8539 = 9'h31 == r_count_28_io_out ? io_r_49_b : _GEN_8538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8540 = 9'h32 == r_count_28_io_out ? io_r_50_b : _GEN_8539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8541 = 9'h33 == r_count_28_io_out ? io_r_51_b : _GEN_8540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8542 = 9'h34 == r_count_28_io_out ? io_r_52_b : _GEN_8541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8543 = 9'h35 == r_count_28_io_out ? io_r_53_b : _GEN_8542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8544 = 9'h36 == r_count_28_io_out ? io_r_54_b : _GEN_8543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8545 = 9'h37 == r_count_28_io_out ? io_r_55_b : _GEN_8544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8546 = 9'h38 == r_count_28_io_out ? io_r_56_b : _GEN_8545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8547 = 9'h39 == r_count_28_io_out ? io_r_57_b : _GEN_8546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8548 = 9'h3a == r_count_28_io_out ? io_r_58_b : _GEN_8547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8549 = 9'h3b == r_count_28_io_out ? io_r_59_b : _GEN_8548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8550 = 9'h3c == r_count_28_io_out ? io_r_60_b : _GEN_8549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8551 = 9'h3d == r_count_28_io_out ? io_r_61_b : _GEN_8550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8552 = 9'h3e == r_count_28_io_out ? io_r_62_b : _GEN_8551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8553 = 9'h3f == r_count_28_io_out ? io_r_63_b : _GEN_8552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8554 = 9'h40 == r_count_28_io_out ? io_r_64_b : _GEN_8553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8555 = 9'h41 == r_count_28_io_out ? io_r_65_b : _GEN_8554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8556 = 9'h42 == r_count_28_io_out ? io_r_66_b : _GEN_8555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8557 = 9'h43 == r_count_28_io_out ? io_r_67_b : _GEN_8556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8558 = 9'h44 == r_count_28_io_out ? io_r_68_b : _GEN_8557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8559 = 9'h45 == r_count_28_io_out ? io_r_69_b : _GEN_8558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8560 = 9'h46 == r_count_28_io_out ? io_r_70_b : _GEN_8559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8561 = 9'h47 == r_count_28_io_out ? io_r_71_b : _GEN_8560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8562 = 9'h48 == r_count_28_io_out ? io_r_72_b : _GEN_8561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8563 = 9'h49 == r_count_28_io_out ? io_r_73_b : _GEN_8562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8564 = 9'h4a == r_count_28_io_out ? io_r_74_b : _GEN_8563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8565 = 9'h4b == r_count_28_io_out ? io_r_75_b : _GEN_8564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8566 = 9'h4c == r_count_28_io_out ? io_r_76_b : _GEN_8565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8567 = 9'h4d == r_count_28_io_out ? io_r_77_b : _GEN_8566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8568 = 9'h4e == r_count_28_io_out ? io_r_78_b : _GEN_8567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8569 = 9'h4f == r_count_28_io_out ? io_r_79_b : _GEN_8568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8570 = 9'h50 == r_count_28_io_out ? io_r_80_b : _GEN_8569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8571 = 9'h51 == r_count_28_io_out ? io_r_81_b : _GEN_8570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8572 = 9'h52 == r_count_28_io_out ? io_r_82_b : _GEN_8571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8573 = 9'h53 == r_count_28_io_out ? io_r_83_b : _GEN_8572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8574 = 9'h54 == r_count_28_io_out ? io_r_84_b : _GEN_8573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8575 = 9'h55 == r_count_28_io_out ? io_r_85_b : _GEN_8574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8576 = 9'h56 == r_count_28_io_out ? io_r_86_b : _GEN_8575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8577 = 9'h57 == r_count_28_io_out ? io_r_87_b : _GEN_8576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8578 = 9'h58 == r_count_28_io_out ? io_r_88_b : _GEN_8577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8579 = 9'h59 == r_count_28_io_out ? io_r_89_b : _GEN_8578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8580 = 9'h5a == r_count_28_io_out ? io_r_90_b : _GEN_8579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8581 = 9'h5b == r_count_28_io_out ? io_r_91_b : _GEN_8580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8582 = 9'h5c == r_count_28_io_out ? io_r_92_b : _GEN_8581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8583 = 9'h5d == r_count_28_io_out ? io_r_93_b : _GEN_8582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8584 = 9'h5e == r_count_28_io_out ? io_r_94_b : _GEN_8583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8585 = 9'h5f == r_count_28_io_out ? io_r_95_b : _GEN_8584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8586 = 9'h60 == r_count_28_io_out ? io_r_96_b : _GEN_8585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8587 = 9'h61 == r_count_28_io_out ? io_r_97_b : _GEN_8586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8588 = 9'h62 == r_count_28_io_out ? io_r_98_b : _GEN_8587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8589 = 9'h63 == r_count_28_io_out ? io_r_99_b : _GEN_8588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8590 = 9'h64 == r_count_28_io_out ? io_r_100_b : _GEN_8589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8591 = 9'h65 == r_count_28_io_out ? io_r_101_b : _GEN_8590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8592 = 9'h66 == r_count_28_io_out ? io_r_102_b : _GEN_8591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8593 = 9'h67 == r_count_28_io_out ? io_r_103_b : _GEN_8592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8594 = 9'h68 == r_count_28_io_out ? io_r_104_b : _GEN_8593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8595 = 9'h69 == r_count_28_io_out ? io_r_105_b : _GEN_8594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8596 = 9'h6a == r_count_28_io_out ? io_r_106_b : _GEN_8595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8597 = 9'h6b == r_count_28_io_out ? io_r_107_b : _GEN_8596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8598 = 9'h6c == r_count_28_io_out ? io_r_108_b : _GEN_8597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8599 = 9'h6d == r_count_28_io_out ? io_r_109_b : _GEN_8598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8600 = 9'h6e == r_count_28_io_out ? io_r_110_b : _GEN_8599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8601 = 9'h6f == r_count_28_io_out ? io_r_111_b : _GEN_8600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8602 = 9'h70 == r_count_28_io_out ? io_r_112_b : _GEN_8601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8603 = 9'h71 == r_count_28_io_out ? io_r_113_b : _GEN_8602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8604 = 9'h72 == r_count_28_io_out ? io_r_114_b : _GEN_8603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8605 = 9'h73 == r_count_28_io_out ? io_r_115_b : _GEN_8604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8606 = 9'h74 == r_count_28_io_out ? io_r_116_b : _GEN_8605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8607 = 9'h75 == r_count_28_io_out ? io_r_117_b : _GEN_8606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8608 = 9'h76 == r_count_28_io_out ? io_r_118_b : _GEN_8607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8609 = 9'h77 == r_count_28_io_out ? io_r_119_b : _GEN_8608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8610 = 9'h78 == r_count_28_io_out ? io_r_120_b : _GEN_8609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8611 = 9'h79 == r_count_28_io_out ? io_r_121_b : _GEN_8610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8612 = 9'h7a == r_count_28_io_out ? io_r_122_b : _GEN_8611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8613 = 9'h7b == r_count_28_io_out ? io_r_123_b : _GEN_8612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8614 = 9'h7c == r_count_28_io_out ? io_r_124_b : _GEN_8613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8615 = 9'h7d == r_count_28_io_out ? io_r_125_b : _GEN_8614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8616 = 9'h7e == r_count_28_io_out ? io_r_126_b : _GEN_8615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8617 = 9'h7f == r_count_28_io_out ? io_r_127_b : _GEN_8616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8618 = 9'h80 == r_count_28_io_out ? io_r_128_b : _GEN_8617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8619 = 9'h81 == r_count_28_io_out ? io_r_129_b : _GEN_8618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8620 = 9'h82 == r_count_28_io_out ? io_r_130_b : _GEN_8619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8621 = 9'h83 == r_count_28_io_out ? io_r_131_b : _GEN_8620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8622 = 9'h84 == r_count_28_io_out ? io_r_132_b : _GEN_8621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8623 = 9'h85 == r_count_28_io_out ? io_r_133_b : _GEN_8622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8624 = 9'h86 == r_count_28_io_out ? io_r_134_b : _GEN_8623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8625 = 9'h87 == r_count_28_io_out ? io_r_135_b : _GEN_8624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8626 = 9'h88 == r_count_28_io_out ? io_r_136_b : _GEN_8625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8627 = 9'h89 == r_count_28_io_out ? io_r_137_b : _GEN_8626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8628 = 9'h8a == r_count_28_io_out ? io_r_138_b : _GEN_8627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8629 = 9'h8b == r_count_28_io_out ? io_r_139_b : _GEN_8628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8630 = 9'h8c == r_count_28_io_out ? io_r_140_b : _GEN_8629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8631 = 9'h8d == r_count_28_io_out ? io_r_141_b : _GEN_8630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8632 = 9'h8e == r_count_28_io_out ? io_r_142_b : _GEN_8631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8633 = 9'h8f == r_count_28_io_out ? io_r_143_b : _GEN_8632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8634 = 9'h90 == r_count_28_io_out ? io_r_144_b : _GEN_8633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8635 = 9'h91 == r_count_28_io_out ? io_r_145_b : _GEN_8634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8636 = 9'h92 == r_count_28_io_out ? io_r_146_b : _GEN_8635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8637 = 9'h93 == r_count_28_io_out ? io_r_147_b : _GEN_8636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8638 = 9'h94 == r_count_28_io_out ? io_r_148_b : _GEN_8637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8639 = 9'h95 == r_count_28_io_out ? io_r_149_b : _GEN_8638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8640 = 9'h96 == r_count_28_io_out ? io_r_150_b : _GEN_8639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8641 = 9'h97 == r_count_28_io_out ? io_r_151_b : _GEN_8640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8642 = 9'h98 == r_count_28_io_out ? io_r_152_b : _GEN_8641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8643 = 9'h99 == r_count_28_io_out ? io_r_153_b : _GEN_8642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8644 = 9'h9a == r_count_28_io_out ? io_r_154_b : _GEN_8643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8645 = 9'h9b == r_count_28_io_out ? io_r_155_b : _GEN_8644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8646 = 9'h9c == r_count_28_io_out ? io_r_156_b : _GEN_8645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8647 = 9'h9d == r_count_28_io_out ? io_r_157_b : _GEN_8646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8648 = 9'h9e == r_count_28_io_out ? io_r_158_b : _GEN_8647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8649 = 9'h9f == r_count_28_io_out ? io_r_159_b : _GEN_8648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8650 = 9'ha0 == r_count_28_io_out ? io_r_160_b : _GEN_8649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8651 = 9'ha1 == r_count_28_io_out ? io_r_161_b : _GEN_8650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8652 = 9'ha2 == r_count_28_io_out ? io_r_162_b : _GEN_8651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8653 = 9'ha3 == r_count_28_io_out ? io_r_163_b : _GEN_8652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8654 = 9'ha4 == r_count_28_io_out ? io_r_164_b : _GEN_8653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8655 = 9'ha5 == r_count_28_io_out ? io_r_165_b : _GEN_8654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8656 = 9'ha6 == r_count_28_io_out ? io_r_166_b : _GEN_8655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8657 = 9'ha7 == r_count_28_io_out ? io_r_167_b : _GEN_8656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8658 = 9'ha8 == r_count_28_io_out ? io_r_168_b : _GEN_8657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8659 = 9'ha9 == r_count_28_io_out ? io_r_169_b : _GEN_8658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8660 = 9'haa == r_count_28_io_out ? io_r_170_b : _GEN_8659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8661 = 9'hab == r_count_28_io_out ? io_r_171_b : _GEN_8660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8662 = 9'hac == r_count_28_io_out ? io_r_172_b : _GEN_8661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8663 = 9'had == r_count_28_io_out ? io_r_173_b : _GEN_8662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8664 = 9'hae == r_count_28_io_out ? io_r_174_b : _GEN_8663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8665 = 9'haf == r_count_28_io_out ? io_r_175_b : _GEN_8664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8666 = 9'hb0 == r_count_28_io_out ? io_r_176_b : _GEN_8665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8667 = 9'hb1 == r_count_28_io_out ? io_r_177_b : _GEN_8666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8668 = 9'hb2 == r_count_28_io_out ? io_r_178_b : _GEN_8667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8669 = 9'hb3 == r_count_28_io_out ? io_r_179_b : _GEN_8668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8670 = 9'hb4 == r_count_28_io_out ? io_r_180_b : _GEN_8669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8671 = 9'hb5 == r_count_28_io_out ? io_r_181_b : _GEN_8670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8672 = 9'hb6 == r_count_28_io_out ? io_r_182_b : _GEN_8671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8673 = 9'hb7 == r_count_28_io_out ? io_r_183_b : _GEN_8672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8674 = 9'hb8 == r_count_28_io_out ? io_r_184_b : _GEN_8673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8675 = 9'hb9 == r_count_28_io_out ? io_r_185_b : _GEN_8674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8676 = 9'hba == r_count_28_io_out ? io_r_186_b : _GEN_8675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8677 = 9'hbb == r_count_28_io_out ? io_r_187_b : _GEN_8676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8678 = 9'hbc == r_count_28_io_out ? io_r_188_b : _GEN_8677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8679 = 9'hbd == r_count_28_io_out ? io_r_189_b : _GEN_8678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8680 = 9'hbe == r_count_28_io_out ? io_r_190_b : _GEN_8679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8681 = 9'hbf == r_count_28_io_out ? io_r_191_b : _GEN_8680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8682 = 9'hc0 == r_count_28_io_out ? io_r_192_b : _GEN_8681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8683 = 9'hc1 == r_count_28_io_out ? io_r_193_b : _GEN_8682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8684 = 9'hc2 == r_count_28_io_out ? io_r_194_b : _GEN_8683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8685 = 9'hc3 == r_count_28_io_out ? io_r_195_b : _GEN_8684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8686 = 9'hc4 == r_count_28_io_out ? io_r_196_b : _GEN_8685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8687 = 9'hc5 == r_count_28_io_out ? io_r_197_b : _GEN_8686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8688 = 9'hc6 == r_count_28_io_out ? io_r_198_b : _GEN_8687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8689 = 9'hc7 == r_count_28_io_out ? io_r_199_b : _GEN_8688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8690 = 9'hc8 == r_count_28_io_out ? io_r_200_b : _GEN_8689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8691 = 9'hc9 == r_count_28_io_out ? io_r_201_b : _GEN_8690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8692 = 9'hca == r_count_28_io_out ? io_r_202_b : _GEN_8691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8693 = 9'hcb == r_count_28_io_out ? io_r_203_b : _GEN_8692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8694 = 9'hcc == r_count_28_io_out ? io_r_204_b : _GEN_8693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8695 = 9'hcd == r_count_28_io_out ? io_r_205_b : _GEN_8694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8696 = 9'hce == r_count_28_io_out ? io_r_206_b : _GEN_8695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8697 = 9'hcf == r_count_28_io_out ? io_r_207_b : _GEN_8696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8698 = 9'hd0 == r_count_28_io_out ? io_r_208_b : _GEN_8697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8699 = 9'hd1 == r_count_28_io_out ? io_r_209_b : _GEN_8698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8700 = 9'hd2 == r_count_28_io_out ? io_r_210_b : _GEN_8699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8701 = 9'hd3 == r_count_28_io_out ? io_r_211_b : _GEN_8700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8702 = 9'hd4 == r_count_28_io_out ? io_r_212_b : _GEN_8701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8703 = 9'hd5 == r_count_28_io_out ? io_r_213_b : _GEN_8702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8704 = 9'hd6 == r_count_28_io_out ? io_r_214_b : _GEN_8703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8705 = 9'hd7 == r_count_28_io_out ? io_r_215_b : _GEN_8704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8706 = 9'hd8 == r_count_28_io_out ? io_r_216_b : _GEN_8705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8707 = 9'hd9 == r_count_28_io_out ? io_r_217_b : _GEN_8706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8708 = 9'hda == r_count_28_io_out ? io_r_218_b : _GEN_8707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8709 = 9'hdb == r_count_28_io_out ? io_r_219_b : _GEN_8708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8710 = 9'hdc == r_count_28_io_out ? io_r_220_b : _GEN_8709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8711 = 9'hdd == r_count_28_io_out ? io_r_221_b : _GEN_8710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8712 = 9'hde == r_count_28_io_out ? io_r_222_b : _GEN_8711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8713 = 9'hdf == r_count_28_io_out ? io_r_223_b : _GEN_8712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8714 = 9'he0 == r_count_28_io_out ? io_r_224_b : _GEN_8713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8715 = 9'he1 == r_count_28_io_out ? io_r_225_b : _GEN_8714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8716 = 9'he2 == r_count_28_io_out ? io_r_226_b : _GEN_8715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8717 = 9'he3 == r_count_28_io_out ? io_r_227_b : _GEN_8716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8718 = 9'he4 == r_count_28_io_out ? io_r_228_b : _GEN_8717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8719 = 9'he5 == r_count_28_io_out ? io_r_229_b : _GEN_8718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8720 = 9'he6 == r_count_28_io_out ? io_r_230_b : _GEN_8719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8721 = 9'he7 == r_count_28_io_out ? io_r_231_b : _GEN_8720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8722 = 9'he8 == r_count_28_io_out ? io_r_232_b : _GEN_8721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8723 = 9'he9 == r_count_28_io_out ? io_r_233_b : _GEN_8722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8724 = 9'hea == r_count_28_io_out ? io_r_234_b : _GEN_8723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8725 = 9'heb == r_count_28_io_out ? io_r_235_b : _GEN_8724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8726 = 9'hec == r_count_28_io_out ? io_r_236_b : _GEN_8725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8727 = 9'hed == r_count_28_io_out ? io_r_237_b : _GEN_8726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8728 = 9'hee == r_count_28_io_out ? io_r_238_b : _GEN_8727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8729 = 9'hef == r_count_28_io_out ? io_r_239_b : _GEN_8728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8730 = 9'hf0 == r_count_28_io_out ? io_r_240_b : _GEN_8729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8731 = 9'hf1 == r_count_28_io_out ? io_r_241_b : _GEN_8730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8732 = 9'hf2 == r_count_28_io_out ? io_r_242_b : _GEN_8731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8733 = 9'hf3 == r_count_28_io_out ? io_r_243_b : _GEN_8732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8734 = 9'hf4 == r_count_28_io_out ? io_r_244_b : _GEN_8733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8735 = 9'hf5 == r_count_28_io_out ? io_r_245_b : _GEN_8734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8736 = 9'hf6 == r_count_28_io_out ? io_r_246_b : _GEN_8735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8737 = 9'hf7 == r_count_28_io_out ? io_r_247_b : _GEN_8736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8738 = 9'hf8 == r_count_28_io_out ? io_r_248_b : _GEN_8737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8739 = 9'hf9 == r_count_28_io_out ? io_r_249_b : _GEN_8738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8740 = 9'hfa == r_count_28_io_out ? io_r_250_b : _GEN_8739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8741 = 9'hfb == r_count_28_io_out ? io_r_251_b : _GEN_8740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8742 = 9'hfc == r_count_28_io_out ? io_r_252_b : _GEN_8741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8743 = 9'hfd == r_count_28_io_out ? io_r_253_b : _GEN_8742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8744 = 9'hfe == r_count_28_io_out ? io_r_254_b : _GEN_8743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8745 = 9'hff == r_count_28_io_out ? io_r_255_b : _GEN_8744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8746 = 9'h100 == r_count_28_io_out ? io_r_256_b : _GEN_8745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8747 = 9'h101 == r_count_28_io_out ? io_r_257_b : _GEN_8746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8748 = 9'h102 == r_count_28_io_out ? io_r_258_b : _GEN_8747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8749 = 9'h103 == r_count_28_io_out ? io_r_259_b : _GEN_8748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8750 = 9'h104 == r_count_28_io_out ? io_r_260_b : _GEN_8749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8751 = 9'h105 == r_count_28_io_out ? io_r_261_b : _GEN_8750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8752 = 9'h106 == r_count_28_io_out ? io_r_262_b : _GEN_8751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8753 = 9'h107 == r_count_28_io_out ? io_r_263_b : _GEN_8752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8754 = 9'h108 == r_count_28_io_out ? io_r_264_b : _GEN_8753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8755 = 9'h109 == r_count_28_io_out ? io_r_265_b : _GEN_8754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8756 = 9'h10a == r_count_28_io_out ? io_r_266_b : _GEN_8755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8757 = 9'h10b == r_count_28_io_out ? io_r_267_b : _GEN_8756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8758 = 9'h10c == r_count_28_io_out ? io_r_268_b : _GEN_8757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8759 = 9'h10d == r_count_28_io_out ? io_r_269_b : _GEN_8758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8760 = 9'h10e == r_count_28_io_out ? io_r_270_b : _GEN_8759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8761 = 9'h10f == r_count_28_io_out ? io_r_271_b : _GEN_8760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8762 = 9'h110 == r_count_28_io_out ? io_r_272_b : _GEN_8761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8763 = 9'h111 == r_count_28_io_out ? io_r_273_b : _GEN_8762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8764 = 9'h112 == r_count_28_io_out ? io_r_274_b : _GEN_8763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8765 = 9'h113 == r_count_28_io_out ? io_r_275_b : _GEN_8764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8766 = 9'h114 == r_count_28_io_out ? io_r_276_b : _GEN_8765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8767 = 9'h115 == r_count_28_io_out ? io_r_277_b : _GEN_8766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8768 = 9'h116 == r_count_28_io_out ? io_r_278_b : _GEN_8767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8769 = 9'h117 == r_count_28_io_out ? io_r_279_b : _GEN_8768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8770 = 9'h118 == r_count_28_io_out ? io_r_280_b : _GEN_8769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8771 = 9'h119 == r_count_28_io_out ? io_r_281_b : _GEN_8770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8772 = 9'h11a == r_count_28_io_out ? io_r_282_b : _GEN_8771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8773 = 9'h11b == r_count_28_io_out ? io_r_283_b : _GEN_8772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8774 = 9'h11c == r_count_28_io_out ? io_r_284_b : _GEN_8773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8775 = 9'h11d == r_count_28_io_out ? io_r_285_b : _GEN_8774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8776 = 9'h11e == r_count_28_io_out ? io_r_286_b : _GEN_8775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8777 = 9'h11f == r_count_28_io_out ? io_r_287_b : _GEN_8776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8778 = 9'h120 == r_count_28_io_out ? io_r_288_b : _GEN_8777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8779 = 9'h121 == r_count_28_io_out ? io_r_289_b : _GEN_8778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8780 = 9'h122 == r_count_28_io_out ? io_r_290_b : _GEN_8779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8781 = 9'h123 == r_count_28_io_out ? io_r_291_b : _GEN_8780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8782 = 9'h124 == r_count_28_io_out ? io_r_292_b : _GEN_8781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8783 = 9'h125 == r_count_28_io_out ? io_r_293_b : _GEN_8782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8784 = 9'h126 == r_count_28_io_out ? io_r_294_b : _GEN_8783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8785 = 9'h127 == r_count_28_io_out ? io_r_295_b : _GEN_8784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8786 = 9'h128 == r_count_28_io_out ? io_r_296_b : _GEN_8785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8787 = 9'h129 == r_count_28_io_out ? io_r_297_b : _GEN_8786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8788 = 9'h12a == r_count_28_io_out ? io_r_298_b : _GEN_8787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8791 = 9'h1 == r_count_29_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8792 = 9'h2 == r_count_29_io_out ? io_r_2_b : _GEN_8791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8793 = 9'h3 == r_count_29_io_out ? io_r_3_b : _GEN_8792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8794 = 9'h4 == r_count_29_io_out ? io_r_4_b : _GEN_8793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8795 = 9'h5 == r_count_29_io_out ? io_r_5_b : _GEN_8794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8796 = 9'h6 == r_count_29_io_out ? io_r_6_b : _GEN_8795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8797 = 9'h7 == r_count_29_io_out ? io_r_7_b : _GEN_8796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8798 = 9'h8 == r_count_29_io_out ? io_r_8_b : _GEN_8797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8799 = 9'h9 == r_count_29_io_out ? io_r_9_b : _GEN_8798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8800 = 9'ha == r_count_29_io_out ? io_r_10_b : _GEN_8799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8801 = 9'hb == r_count_29_io_out ? io_r_11_b : _GEN_8800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8802 = 9'hc == r_count_29_io_out ? io_r_12_b : _GEN_8801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8803 = 9'hd == r_count_29_io_out ? io_r_13_b : _GEN_8802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8804 = 9'he == r_count_29_io_out ? io_r_14_b : _GEN_8803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8805 = 9'hf == r_count_29_io_out ? io_r_15_b : _GEN_8804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8806 = 9'h10 == r_count_29_io_out ? io_r_16_b : _GEN_8805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8807 = 9'h11 == r_count_29_io_out ? io_r_17_b : _GEN_8806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8808 = 9'h12 == r_count_29_io_out ? io_r_18_b : _GEN_8807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8809 = 9'h13 == r_count_29_io_out ? io_r_19_b : _GEN_8808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8810 = 9'h14 == r_count_29_io_out ? io_r_20_b : _GEN_8809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8811 = 9'h15 == r_count_29_io_out ? io_r_21_b : _GEN_8810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8812 = 9'h16 == r_count_29_io_out ? io_r_22_b : _GEN_8811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8813 = 9'h17 == r_count_29_io_out ? io_r_23_b : _GEN_8812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8814 = 9'h18 == r_count_29_io_out ? io_r_24_b : _GEN_8813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8815 = 9'h19 == r_count_29_io_out ? io_r_25_b : _GEN_8814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8816 = 9'h1a == r_count_29_io_out ? io_r_26_b : _GEN_8815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8817 = 9'h1b == r_count_29_io_out ? io_r_27_b : _GEN_8816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8818 = 9'h1c == r_count_29_io_out ? io_r_28_b : _GEN_8817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8819 = 9'h1d == r_count_29_io_out ? io_r_29_b : _GEN_8818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8820 = 9'h1e == r_count_29_io_out ? io_r_30_b : _GEN_8819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8821 = 9'h1f == r_count_29_io_out ? io_r_31_b : _GEN_8820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8822 = 9'h20 == r_count_29_io_out ? io_r_32_b : _GEN_8821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8823 = 9'h21 == r_count_29_io_out ? io_r_33_b : _GEN_8822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8824 = 9'h22 == r_count_29_io_out ? io_r_34_b : _GEN_8823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8825 = 9'h23 == r_count_29_io_out ? io_r_35_b : _GEN_8824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8826 = 9'h24 == r_count_29_io_out ? io_r_36_b : _GEN_8825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8827 = 9'h25 == r_count_29_io_out ? io_r_37_b : _GEN_8826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8828 = 9'h26 == r_count_29_io_out ? io_r_38_b : _GEN_8827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8829 = 9'h27 == r_count_29_io_out ? io_r_39_b : _GEN_8828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8830 = 9'h28 == r_count_29_io_out ? io_r_40_b : _GEN_8829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8831 = 9'h29 == r_count_29_io_out ? io_r_41_b : _GEN_8830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8832 = 9'h2a == r_count_29_io_out ? io_r_42_b : _GEN_8831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8833 = 9'h2b == r_count_29_io_out ? io_r_43_b : _GEN_8832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8834 = 9'h2c == r_count_29_io_out ? io_r_44_b : _GEN_8833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8835 = 9'h2d == r_count_29_io_out ? io_r_45_b : _GEN_8834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8836 = 9'h2e == r_count_29_io_out ? io_r_46_b : _GEN_8835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8837 = 9'h2f == r_count_29_io_out ? io_r_47_b : _GEN_8836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8838 = 9'h30 == r_count_29_io_out ? io_r_48_b : _GEN_8837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8839 = 9'h31 == r_count_29_io_out ? io_r_49_b : _GEN_8838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8840 = 9'h32 == r_count_29_io_out ? io_r_50_b : _GEN_8839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8841 = 9'h33 == r_count_29_io_out ? io_r_51_b : _GEN_8840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8842 = 9'h34 == r_count_29_io_out ? io_r_52_b : _GEN_8841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8843 = 9'h35 == r_count_29_io_out ? io_r_53_b : _GEN_8842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8844 = 9'h36 == r_count_29_io_out ? io_r_54_b : _GEN_8843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8845 = 9'h37 == r_count_29_io_out ? io_r_55_b : _GEN_8844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8846 = 9'h38 == r_count_29_io_out ? io_r_56_b : _GEN_8845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8847 = 9'h39 == r_count_29_io_out ? io_r_57_b : _GEN_8846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8848 = 9'h3a == r_count_29_io_out ? io_r_58_b : _GEN_8847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8849 = 9'h3b == r_count_29_io_out ? io_r_59_b : _GEN_8848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8850 = 9'h3c == r_count_29_io_out ? io_r_60_b : _GEN_8849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8851 = 9'h3d == r_count_29_io_out ? io_r_61_b : _GEN_8850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8852 = 9'h3e == r_count_29_io_out ? io_r_62_b : _GEN_8851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8853 = 9'h3f == r_count_29_io_out ? io_r_63_b : _GEN_8852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8854 = 9'h40 == r_count_29_io_out ? io_r_64_b : _GEN_8853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8855 = 9'h41 == r_count_29_io_out ? io_r_65_b : _GEN_8854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8856 = 9'h42 == r_count_29_io_out ? io_r_66_b : _GEN_8855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8857 = 9'h43 == r_count_29_io_out ? io_r_67_b : _GEN_8856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8858 = 9'h44 == r_count_29_io_out ? io_r_68_b : _GEN_8857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8859 = 9'h45 == r_count_29_io_out ? io_r_69_b : _GEN_8858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8860 = 9'h46 == r_count_29_io_out ? io_r_70_b : _GEN_8859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8861 = 9'h47 == r_count_29_io_out ? io_r_71_b : _GEN_8860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8862 = 9'h48 == r_count_29_io_out ? io_r_72_b : _GEN_8861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8863 = 9'h49 == r_count_29_io_out ? io_r_73_b : _GEN_8862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8864 = 9'h4a == r_count_29_io_out ? io_r_74_b : _GEN_8863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8865 = 9'h4b == r_count_29_io_out ? io_r_75_b : _GEN_8864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8866 = 9'h4c == r_count_29_io_out ? io_r_76_b : _GEN_8865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8867 = 9'h4d == r_count_29_io_out ? io_r_77_b : _GEN_8866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8868 = 9'h4e == r_count_29_io_out ? io_r_78_b : _GEN_8867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8869 = 9'h4f == r_count_29_io_out ? io_r_79_b : _GEN_8868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8870 = 9'h50 == r_count_29_io_out ? io_r_80_b : _GEN_8869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8871 = 9'h51 == r_count_29_io_out ? io_r_81_b : _GEN_8870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8872 = 9'h52 == r_count_29_io_out ? io_r_82_b : _GEN_8871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8873 = 9'h53 == r_count_29_io_out ? io_r_83_b : _GEN_8872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8874 = 9'h54 == r_count_29_io_out ? io_r_84_b : _GEN_8873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8875 = 9'h55 == r_count_29_io_out ? io_r_85_b : _GEN_8874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8876 = 9'h56 == r_count_29_io_out ? io_r_86_b : _GEN_8875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8877 = 9'h57 == r_count_29_io_out ? io_r_87_b : _GEN_8876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8878 = 9'h58 == r_count_29_io_out ? io_r_88_b : _GEN_8877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8879 = 9'h59 == r_count_29_io_out ? io_r_89_b : _GEN_8878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8880 = 9'h5a == r_count_29_io_out ? io_r_90_b : _GEN_8879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8881 = 9'h5b == r_count_29_io_out ? io_r_91_b : _GEN_8880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8882 = 9'h5c == r_count_29_io_out ? io_r_92_b : _GEN_8881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8883 = 9'h5d == r_count_29_io_out ? io_r_93_b : _GEN_8882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8884 = 9'h5e == r_count_29_io_out ? io_r_94_b : _GEN_8883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8885 = 9'h5f == r_count_29_io_out ? io_r_95_b : _GEN_8884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8886 = 9'h60 == r_count_29_io_out ? io_r_96_b : _GEN_8885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8887 = 9'h61 == r_count_29_io_out ? io_r_97_b : _GEN_8886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8888 = 9'h62 == r_count_29_io_out ? io_r_98_b : _GEN_8887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8889 = 9'h63 == r_count_29_io_out ? io_r_99_b : _GEN_8888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8890 = 9'h64 == r_count_29_io_out ? io_r_100_b : _GEN_8889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8891 = 9'h65 == r_count_29_io_out ? io_r_101_b : _GEN_8890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8892 = 9'h66 == r_count_29_io_out ? io_r_102_b : _GEN_8891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8893 = 9'h67 == r_count_29_io_out ? io_r_103_b : _GEN_8892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8894 = 9'h68 == r_count_29_io_out ? io_r_104_b : _GEN_8893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8895 = 9'h69 == r_count_29_io_out ? io_r_105_b : _GEN_8894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8896 = 9'h6a == r_count_29_io_out ? io_r_106_b : _GEN_8895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8897 = 9'h6b == r_count_29_io_out ? io_r_107_b : _GEN_8896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8898 = 9'h6c == r_count_29_io_out ? io_r_108_b : _GEN_8897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8899 = 9'h6d == r_count_29_io_out ? io_r_109_b : _GEN_8898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8900 = 9'h6e == r_count_29_io_out ? io_r_110_b : _GEN_8899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8901 = 9'h6f == r_count_29_io_out ? io_r_111_b : _GEN_8900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8902 = 9'h70 == r_count_29_io_out ? io_r_112_b : _GEN_8901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8903 = 9'h71 == r_count_29_io_out ? io_r_113_b : _GEN_8902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8904 = 9'h72 == r_count_29_io_out ? io_r_114_b : _GEN_8903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8905 = 9'h73 == r_count_29_io_out ? io_r_115_b : _GEN_8904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8906 = 9'h74 == r_count_29_io_out ? io_r_116_b : _GEN_8905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8907 = 9'h75 == r_count_29_io_out ? io_r_117_b : _GEN_8906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8908 = 9'h76 == r_count_29_io_out ? io_r_118_b : _GEN_8907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8909 = 9'h77 == r_count_29_io_out ? io_r_119_b : _GEN_8908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8910 = 9'h78 == r_count_29_io_out ? io_r_120_b : _GEN_8909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8911 = 9'h79 == r_count_29_io_out ? io_r_121_b : _GEN_8910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8912 = 9'h7a == r_count_29_io_out ? io_r_122_b : _GEN_8911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8913 = 9'h7b == r_count_29_io_out ? io_r_123_b : _GEN_8912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8914 = 9'h7c == r_count_29_io_out ? io_r_124_b : _GEN_8913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8915 = 9'h7d == r_count_29_io_out ? io_r_125_b : _GEN_8914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8916 = 9'h7e == r_count_29_io_out ? io_r_126_b : _GEN_8915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8917 = 9'h7f == r_count_29_io_out ? io_r_127_b : _GEN_8916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8918 = 9'h80 == r_count_29_io_out ? io_r_128_b : _GEN_8917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8919 = 9'h81 == r_count_29_io_out ? io_r_129_b : _GEN_8918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8920 = 9'h82 == r_count_29_io_out ? io_r_130_b : _GEN_8919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8921 = 9'h83 == r_count_29_io_out ? io_r_131_b : _GEN_8920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8922 = 9'h84 == r_count_29_io_out ? io_r_132_b : _GEN_8921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8923 = 9'h85 == r_count_29_io_out ? io_r_133_b : _GEN_8922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8924 = 9'h86 == r_count_29_io_out ? io_r_134_b : _GEN_8923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8925 = 9'h87 == r_count_29_io_out ? io_r_135_b : _GEN_8924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8926 = 9'h88 == r_count_29_io_out ? io_r_136_b : _GEN_8925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8927 = 9'h89 == r_count_29_io_out ? io_r_137_b : _GEN_8926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8928 = 9'h8a == r_count_29_io_out ? io_r_138_b : _GEN_8927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8929 = 9'h8b == r_count_29_io_out ? io_r_139_b : _GEN_8928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8930 = 9'h8c == r_count_29_io_out ? io_r_140_b : _GEN_8929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8931 = 9'h8d == r_count_29_io_out ? io_r_141_b : _GEN_8930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8932 = 9'h8e == r_count_29_io_out ? io_r_142_b : _GEN_8931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8933 = 9'h8f == r_count_29_io_out ? io_r_143_b : _GEN_8932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8934 = 9'h90 == r_count_29_io_out ? io_r_144_b : _GEN_8933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8935 = 9'h91 == r_count_29_io_out ? io_r_145_b : _GEN_8934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8936 = 9'h92 == r_count_29_io_out ? io_r_146_b : _GEN_8935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8937 = 9'h93 == r_count_29_io_out ? io_r_147_b : _GEN_8936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8938 = 9'h94 == r_count_29_io_out ? io_r_148_b : _GEN_8937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8939 = 9'h95 == r_count_29_io_out ? io_r_149_b : _GEN_8938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8940 = 9'h96 == r_count_29_io_out ? io_r_150_b : _GEN_8939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8941 = 9'h97 == r_count_29_io_out ? io_r_151_b : _GEN_8940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8942 = 9'h98 == r_count_29_io_out ? io_r_152_b : _GEN_8941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8943 = 9'h99 == r_count_29_io_out ? io_r_153_b : _GEN_8942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8944 = 9'h9a == r_count_29_io_out ? io_r_154_b : _GEN_8943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8945 = 9'h9b == r_count_29_io_out ? io_r_155_b : _GEN_8944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8946 = 9'h9c == r_count_29_io_out ? io_r_156_b : _GEN_8945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8947 = 9'h9d == r_count_29_io_out ? io_r_157_b : _GEN_8946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8948 = 9'h9e == r_count_29_io_out ? io_r_158_b : _GEN_8947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8949 = 9'h9f == r_count_29_io_out ? io_r_159_b : _GEN_8948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8950 = 9'ha0 == r_count_29_io_out ? io_r_160_b : _GEN_8949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8951 = 9'ha1 == r_count_29_io_out ? io_r_161_b : _GEN_8950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8952 = 9'ha2 == r_count_29_io_out ? io_r_162_b : _GEN_8951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8953 = 9'ha3 == r_count_29_io_out ? io_r_163_b : _GEN_8952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8954 = 9'ha4 == r_count_29_io_out ? io_r_164_b : _GEN_8953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8955 = 9'ha5 == r_count_29_io_out ? io_r_165_b : _GEN_8954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8956 = 9'ha6 == r_count_29_io_out ? io_r_166_b : _GEN_8955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8957 = 9'ha7 == r_count_29_io_out ? io_r_167_b : _GEN_8956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8958 = 9'ha8 == r_count_29_io_out ? io_r_168_b : _GEN_8957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8959 = 9'ha9 == r_count_29_io_out ? io_r_169_b : _GEN_8958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8960 = 9'haa == r_count_29_io_out ? io_r_170_b : _GEN_8959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8961 = 9'hab == r_count_29_io_out ? io_r_171_b : _GEN_8960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8962 = 9'hac == r_count_29_io_out ? io_r_172_b : _GEN_8961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8963 = 9'had == r_count_29_io_out ? io_r_173_b : _GEN_8962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8964 = 9'hae == r_count_29_io_out ? io_r_174_b : _GEN_8963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8965 = 9'haf == r_count_29_io_out ? io_r_175_b : _GEN_8964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8966 = 9'hb0 == r_count_29_io_out ? io_r_176_b : _GEN_8965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8967 = 9'hb1 == r_count_29_io_out ? io_r_177_b : _GEN_8966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8968 = 9'hb2 == r_count_29_io_out ? io_r_178_b : _GEN_8967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8969 = 9'hb3 == r_count_29_io_out ? io_r_179_b : _GEN_8968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8970 = 9'hb4 == r_count_29_io_out ? io_r_180_b : _GEN_8969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8971 = 9'hb5 == r_count_29_io_out ? io_r_181_b : _GEN_8970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8972 = 9'hb6 == r_count_29_io_out ? io_r_182_b : _GEN_8971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8973 = 9'hb7 == r_count_29_io_out ? io_r_183_b : _GEN_8972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8974 = 9'hb8 == r_count_29_io_out ? io_r_184_b : _GEN_8973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8975 = 9'hb9 == r_count_29_io_out ? io_r_185_b : _GEN_8974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8976 = 9'hba == r_count_29_io_out ? io_r_186_b : _GEN_8975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8977 = 9'hbb == r_count_29_io_out ? io_r_187_b : _GEN_8976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8978 = 9'hbc == r_count_29_io_out ? io_r_188_b : _GEN_8977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8979 = 9'hbd == r_count_29_io_out ? io_r_189_b : _GEN_8978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8980 = 9'hbe == r_count_29_io_out ? io_r_190_b : _GEN_8979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8981 = 9'hbf == r_count_29_io_out ? io_r_191_b : _GEN_8980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8982 = 9'hc0 == r_count_29_io_out ? io_r_192_b : _GEN_8981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8983 = 9'hc1 == r_count_29_io_out ? io_r_193_b : _GEN_8982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8984 = 9'hc2 == r_count_29_io_out ? io_r_194_b : _GEN_8983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8985 = 9'hc3 == r_count_29_io_out ? io_r_195_b : _GEN_8984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8986 = 9'hc4 == r_count_29_io_out ? io_r_196_b : _GEN_8985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8987 = 9'hc5 == r_count_29_io_out ? io_r_197_b : _GEN_8986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8988 = 9'hc6 == r_count_29_io_out ? io_r_198_b : _GEN_8987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8989 = 9'hc7 == r_count_29_io_out ? io_r_199_b : _GEN_8988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8990 = 9'hc8 == r_count_29_io_out ? io_r_200_b : _GEN_8989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8991 = 9'hc9 == r_count_29_io_out ? io_r_201_b : _GEN_8990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8992 = 9'hca == r_count_29_io_out ? io_r_202_b : _GEN_8991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8993 = 9'hcb == r_count_29_io_out ? io_r_203_b : _GEN_8992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8994 = 9'hcc == r_count_29_io_out ? io_r_204_b : _GEN_8993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8995 = 9'hcd == r_count_29_io_out ? io_r_205_b : _GEN_8994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8996 = 9'hce == r_count_29_io_out ? io_r_206_b : _GEN_8995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8997 = 9'hcf == r_count_29_io_out ? io_r_207_b : _GEN_8996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8998 = 9'hd0 == r_count_29_io_out ? io_r_208_b : _GEN_8997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8999 = 9'hd1 == r_count_29_io_out ? io_r_209_b : _GEN_8998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9000 = 9'hd2 == r_count_29_io_out ? io_r_210_b : _GEN_8999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9001 = 9'hd3 == r_count_29_io_out ? io_r_211_b : _GEN_9000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9002 = 9'hd4 == r_count_29_io_out ? io_r_212_b : _GEN_9001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9003 = 9'hd5 == r_count_29_io_out ? io_r_213_b : _GEN_9002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9004 = 9'hd6 == r_count_29_io_out ? io_r_214_b : _GEN_9003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9005 = 9'hd7 == r_count_29_io_out ? io_r_215_b : _GEN_9004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9006 = 9'hd8 == r_count_29_io_out ? io_r_216_b : _GEN_9005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9007 = 9'hd9 == r_count_29_io_out ? io_r_217_b : _GEN_9006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9008 = 9'hda == r_count_29_io_out ? io_r_218_b : _GEN_9007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9009 = 9'hdb == r_count_29_io_out ? io_r_219_b : _GEN_9008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9010 = 9'hdc == r_count_29_io_out ? io_r_220_b : _GEN_9009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9011 = 9'hdd == r_count_29_io_out ? io_r_221_b : _GEN_9010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9012 = 9'hde == r_count_29_io_out ? io_r_222_b : _GEN_9011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9013 = 9'hdf == r_count_29_io_out ? io_r_223_b : _GEN_9012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9014 = 9'he0 == r_count_29_io_out ? io_r_224_b : _GEN_9013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9015 = 9'he1 == r_count_29_io_out ? io_r_225_b : _GEN_9014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9016 = 9'he2 == r_count_29_io_out ? io_r_226_b : _GEN_9015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9017 = 9'he3 == r_count_29_io_out ? io_r_227_b : _GEN_9016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9018 = 9'he4 == r_count_29_io_out ? io_r_228_b : _GEN_9017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9019 = 9'he5 == r_count_29_io_out ? io_r_229_b : _GEN_9018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9020 = 9'he6 == r_count_29_io_out ? io_r_230_b : _GEN_9019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9021 = 9'he7 == r_count_29_io_out ? io_r_231_b : _GEN_9020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9022 = 9'he8 == r_count_29_io_out ? io_r_232_b : _GEN_9021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9023 = 9'he9 == r_count_29_io_out ? io_r_233_b : _GEN_9022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9024 = 9'hea == r_count_29_io_out ? io_r_234_b : _GEN_9023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9025 = 9'heb == r_count_29_io_out ? io_r_235_b : _GEN_9024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9026 = 9'hec == r_count_29_io_out ? io_r_236_b : _GEN_9025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9027 = 9'hed == r_count_29_io_out ? io_r_237_b : _GEN_9026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9028 = 9'hee == r_count_29_io_out ? io_r_238_b : _GEN_9027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9029 = 9'hef == r_count_29_io_out ? io_r_239_b : _GEN_9028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9030 = 9'hf0 == r_count_29_io_out ? io_r_240_b : _GEN_9029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9031 = 9'hf1 == r_count_29_io_out ? io_r_241_b : _GEN_9030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9032 = 9'hf2 == r_count_29_io_out ? io_r_242_b : _GEN_9031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9033 = 9'hf3 == r_count_29_io_out ? io_r_243_b : _GEN_9032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9034 = 9'hf4 == r_count_29_io_out ? io_r_244_b : _GEN_9033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9035 = 9'hf5 == r_count_29_io_out ? io_r_245_b : _GEN_9034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9036 = 9'hf6 == r_count_29_io_out ? io_r_246_b : _GEN_9035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9037 = 9'hf7 == r_count_29_io_out ? io_r_247_b : _GEN_9036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9038 = 9'hf8 == r_count_29_io_out ? io_r_248_b : _GEN_9037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9039 = 9'hf9 == r_count_29_io_out ? io_r_249_b : _GEN_9038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9040 = 9'hfa == r_count_29_io_out ? io_r_250_b : _GEN_9039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9041 = 9'hfb == r_count_29_io_out ? io_r_251_b : _GEN_9040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9042 = 9'hfc == r_count_29_io_out ? io_r_252_b : _GEN_9041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9043 = 9'hfd == r_count_29_io_out ? io_r_253_b : _GEN_9042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9044 = 9'hfe == r_count_29_io_out ? io_r_254_b : _GEN_9043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9045 = 9'hff == r_count_29_io_out ? io_r_255_b : _GEN_9044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9046 = 9'h100 == r_count_29_io_out ? io_r_256_b : _GEN_9045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9047 = 9'h101 == r_count_29_io_out ? io_r_257_b : _GEN_9046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9048 = 9'h102 == r_count_29_io_out ? io_r_258_b : _GEN_9047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9049 = 9'h103 == r_count_29_io_out ? io_r_259_b : _GEN_9048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9050 = 9'h104 == r_count_29_io_out ? io_r_260_b : _GEN_9049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9051 = 9'h105 == r_count_29_io_out ? io_r_261_b : _GEN_9050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9052 = 9'h106 == r_count_29_io_out ? io_r_262_b : _GEN_9051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9053 = 9'h107 == r_count_29_io_out ? io_r_263_b : _GEN_9052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9054 = 9'h108 == r_count_29_io_out ? io_r_264_b : _GEN_9053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9055 = 9'h109 == r_count_29_io_out ? io_r_265_b : _GEN_9054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9056 = 9'h10a == r_count_29_io_out ? io_r_266_b : _GEN_9055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9057 = 9'h10b == r_count_29_io_out ? io_r_267_b : _GEN_9056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9058 = 9'h10c == r_count_29_io_out ? io_r_268_b : _GEN_9057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9059 = 9'h10d == r_count_29_io_out ? io_r_269_b : _GEN_9058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9060 = 9'h10e == r_count_29_io_out ? io_r_270_b : _GEN_9059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9061 = 9'h10f == r_count_29_io_out ? io_r_271_b : _GEN_9060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9062 = 9'h110 == r_count_29_io_out ? io_r_272_b : _GEN_9061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9063 = 9'h111 == r_count_29_io_out ? io_r_273_b : _GEN_9062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9064 = 9'h112 == r_count_29_io_out ? io_r_274_b : _GEN_9063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9065 = 9'h113 == r_count_29_io_out ? io_r_275_b : _GEN_9064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9066 = 9'h114 == r_count_29_io_out ? io_r_276_b : _GEN_9065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9067 = 9'h115 == r_count_29_io_out ? io_r_277_b : _GEN_9066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9068 = 9'h116 == r_count_29_io_out ? io_r_278_b : _GEN_9067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9069 = 9'h117 == r_count_29_io_out ? io_r_279_b : _GEN_9068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9070 = 9'h118 == r_count_29_io_out ? io_r_280_b : _GEN_9069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9071 = 9'h119 == r_count_29_io_out ? io_r_281_b : _GEN_9070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9072 = 9'h11a == r_count_29_io_out ? io_r_282_b : _GEN_9071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9073 = 9'h11b == r_count_29_io_out ? io_r_283_b : _GEN_9072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9074 = 9'h11c == r_count_29_io_out ? io_r_284_b : _GEN_9073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9075 = 9'h11d == r_count_29_io_out ? io_r_285_b : _GEN_9074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9076 = 9'h11e == r_count_29_io_out ? io_r_286_b : _GEN_9075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9077 = 9'h11f == r_count_29_io_out ? io_r_287_b : _GEN_9076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9078 = 9'h120 == r_count_29_io_out ? io_r_288_b : _GEN_9077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9079 = 9'h121 == r_count_29_io_out ? io_r_289_b : _GEN_9078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9080 = 9'h122 == r_count_29_io_out ? io_r_290_b : _GEN_9079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9081 = 9'h123 == r_count_29_io_out ? io_r_291_b : _GEN_9080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9082 = 9'h124 == r_count_29_io_out ? io_r_292_b : _GEN_9081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9083 = 9'h125 == r_count_29_io_out ? io_r_293_b : _GEN_9082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9084 = 9'h126 == r_count_29_io_out ? io_r_294_b : _GEN_9083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9085 = 9'h127 == r_count_29_io_out ? io_r_295_b : _GEN_9084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9086 = 9'h128 == r_count_29_io_out ? io_r_296_b : _GEN_9085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9087 = 9'h129 == r_count_29_io_out ? io_r_297_b : _GEN_9086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9088 = 9'h12a == r_count_29_io_out ? io_r_298_b : _GEN_9087; // @[SWChisel.scala 221:{19,19}]
  SWCell array_0 ( // @[SWChisel.scala 170:39]
    .io_q(array_0_io_q),
    .io_r(array_0_io_r),
    .io_e_i(array_0_io_e_i),
    .io_f_i(array_0_io_f_i),
    .io_ve_i(array_0_io_ve_i),
    .io_vf_i(array_0_io_vf_i),
    .io_vv_i(array_0_io_vv_i),
    .io_e_o(array_0_io_e_o),
    .io_f_o(array_0_io_f_o),
    .io_v_o(array_0_io_v_o)
  );
  SWCell array_1 ( // @[SWChisel.scala 170:39]
    .io_q(array_1_io_q),
    .io_r(array_1_io_r),
    .io_e_i(array_1_io_e_i),
    .io_f_i(array_1_io_f_i),
    .io_ve_i(array_1_io_ve_i),
    .io_vf_i(array_1_io_vf_i),
    .io_vv_i(array_1_io_vv_i),
    .io_e_o(array_1_io_e_o),
    .io_f_o(array_1_io_f_o),
    .io_v_o(array_1_io_v_o)
  );
  SWCell array_2 ( // @[SWChisel.scala 170:39]
    .io_q(array_2_io_q),
    .io_r(array_2_io_r),
    .io_e_i(array_2_io_e_i),
    .io_f_i(array_2_io_f_i),
    .io_ve_i(array_2_io_ve_i),
    .io_vf_i(array_2_io_vf_i),
    .io_vv_i(array_2_io_vv_i),
    .io_e_o(array_2_io_e_o),
    .io_f_o(array_2_io_f_o),
    .io_v_o(array_2_io_v_o)
  );
  SWCell array_3 ( // @[SWChisel.scala 170:39]
    .io_q(array_3_io_q),
    .io_r(array_3_io_r),
    .io_e_i(array_3_io_e_i),
    .io_f_i(array_3_io_f_i),
    .io_ve_i(array_3_io_ve_i),
    .io_vf_i(array_3_io_vf_i),
    .io_vv_i(array_3_io_vv_i),
    .io_e_o(array_3_io_e_o),
    .io_f_o(array_3_io_f_o),
    .io_v_o(array_3_io_v_o)
  );
  SWCell array_4 ( // @[SWChisel.scala 170:39]
    .io_q(array_4_io_q),
    .io_r(array_4_io_r),
    .io_e_i(array_4_io_e_i),
    .io_f_i(array_4_io_f_i),
    .io_ve_i(array_4_io_ve_i),
    .io_vf_i(array_4_io_vf_i),
    .io_vv_i(array_4_io_vv_i),
    .io_e_o(array_4_io_e_o),
    .io_f_o(array_4_io_f_o),
    .io_v_o(array_4_io_v_o)
  );
  SWCell array_5 ( // @[SWChisel.scala 170:39]
    .io_q(array_5_io_q),
    .io_r(array_5_io_r),
    .io_e_i(array_5_io_e_i),
    .io_f_i(array_5_io_f_i),
    .io_ve_i(array_5_io_ve_i),
    .io_vf_i(array_5_io_vf_i),
    .io_vv_i(array_5_io_vv_i),
    .io_e_o(array_5_io_e_o),
    .io_f_o(array_5_io_f_o),
    .io_v_o(array_5_io_v_o)
  );
  SWCell array_6 ( // @[SWChisel.scala 170:39]
    .io_q(array_6_io_q),
    .io_r(array_6_io_r),
    .io_e_i(array_6_io_e_i),
    .io_f_i(array_6_io_f_i),
    .io_ve_i(array_6_io_ve_i),
    .io_vf_i(array_6_io_vf_i),
    .io_vv_i(array_6_io_vv_i),
    .io_e_o(array_6_io_e_o),
    .io_f_o(array_6_io_f_o),
    .io_v_o(array_6_io_v_o)
  );
  SWCell array_7 ( // @[SWChisel.scala 170:39]
    .io_q(array_7_io_q),
    .io_r(array_7_io_r),
    .io_e_i(array_7_io_e_i),
    .io_f_i(array_7_io_f_i),
    .io_ve_i(array_7_io_ve_i),
    .io_vf_i(array_7_io_vf_i),
    .io_vv_i(array_7_io_vv_i),
    .io_e_o(array_7_io_e_o),
    .io_f_o(array_7_io_f_o),
    .io_v_o(array_7_io_v_o)
  );
  SWCell array_8 ( // @[SWChisel.scala 170:39]
    .io_q(array_8_io_q),
    .io_r(array_8_io_r),
    .io_e_i(array_8_io_e_i),
    .io_f_i(array_8_io_f_i),
    .io_ve_i(array_8_io_ve_i),
    .io_vf_i(array_8_io_vf_i),
    .io_vv_i(array_8_io_vv_i),
    .io_e_o(array_8_io_e_o),
    .io_f_o(array_8_io_f_o),
    .io_v_o(array_8_io_v_o)
  );
  SWCell array_9 ( // @[SWChisel.scala 170:39]
    .io_q(array_9_io_q),
    .io_r(array_9_io_r),
    .io_e_i(array_9_io_e_i),
    .io_f_i(array_9_io_f_i),
    .io_ve_i(array_9_io_ve_i),
    .io_vf_i(array_9_io_vf_i),
    .io_vv_i(array_9_io_vv_i),
    .io_e_o(array_9_io_e_o),
    .io_f_o(array_9_io_f_o),
    .io_v_o(array_9_io_v_o)
  );
  SWCell array_10 ( // @[SWChisel.scala 170:39]
    .io_q(array_10_io_q),
    .io_r(array_10_io_r),
    .io_e_i(array_10_io_e_i),
    .io_f_i(array_10_io_f_i),
    .io_ve_i(array_10_io_ve_i),
    .io_vf_i(array_10_io_vf_i),
    .io_vv_i(array_10_io_vv_i),
    .io_e_o(array_10_io_e_o),
    .io_f_o(array_10_io_f_o),
    .io_v_o(array_10_io_v_o)
  );
  SWCell array_11 ( // @[SWChisel.scala 170:39]
    .io_q(array_11_io_q),
    .io_r(array_11_io_r),
    .io_e_i(array_11_io_e_i),
    .io_f_i(array_11_io_f_i),
    .io_ve_i(array_11_io_ve_i),
    .io_vf_i(array_11_io_vf_i),
    .io_vv_i(array_11_io_vv_i),
    .io_e_o(array_11_io_e_o),
    .io_f_o(array_11_io_f_o),
    .io_v_o(array_11_io_v_o)
  );
  SWCell array_12 ( // @[SWChisel.scala 170:39]
    .io_q(array_12_io_q),
    .io_r(array_12_io_r),
    .io_e_i(array_12_io_e_i),
    .io_f_i(array_12_io_f_i),
    .io_ve_i(array_12_io_ve_i),
    .io_vf_i(array_12_io_vf_i),
    .io_vv_i(array_12_io_vv_i),
    .io_e_o(array_12_io_e_o),
    .io_f_o(array_12_io_f_o),
    .io_v_o(array_12_io_v_o)
  );
  SWCell array_13 ( // @[SWChisel.scala 170:39]
    .io_q(array_13_io_q),
    .io_r(array_13_io_r),
    .io_e_i(array_13_io_e_i),
    .io_f_i(array_13_io_f_i),
    .io_ve_i(array_13_io_ve_i),
    .io_vf_i(array_13_io_vf_i),
    .io_vv_i(array_13_io_vv_i),
    .io_e_o(array_13_io_e_o),
    .io_f_o(array_13_io_f_o),
    .io_v_o(array_13_io_v_o)
  );
  SWCell array_14 ( // @[SWChisel.scala 170:39]
    .io_q(array_14_io_q),
    .io_r(array_14_io_r),
    .io_e_i(array_14_io_e_i),
    .io_f_i(array_14_io_f_i),
    .io_ve_i(array_14_io_ve_i),
    .io_vf_i(array_14_io_vf_i),
    .io_vv_i(array_14_io_vv_i),
    .io_e_o(array_14_io_e_o),
    .io_f_o(array_14_io_f_o),
    .io_v_o(array_14_io_v_o)
  );
  SWCell array_15 ( // @[SWChisel.scala 170:39]
    .io_q(array_15_io_q),
    .io_r(array_15_io_r),
    .io_e_i(array_15_io_e_i),
    .io_f_i(array_15_io_f_i),
    .io_ve_i(array_15_io_ve_i),
    .io_vf_i(array_15_io_vf_i),
    .io_vv_i(array_15_io_vv_i),
    .io_e_o(array_15_io_e_o),
    .io_f_o(array_15_io_f_o),
    .io_v_o(array_15_io_v_o)
  );
  SWCell array_16 ( // @[SWChisel.scala 170:39]
    .io_q(array_16_io_q),
    .io_r(array_16_io_r),
    .io_e_i(array_16_io_e_i),
    .io_f_i(array_16_io_f_i),
    .io_ve_i(array_16_io_ve_i),
    .io_vf_i(array_16_io_vf_i),
    .io_vv_i(array_16_io_vv_i),
    .io_e_o(array_16_io_e_o),
    .io_f_o(array_16_io_f_o),
    .io_v_o(array_16_io_v_o)
  );
  SWCell array_17 ( // @[SWChisel.scala 170:39]
    .io_q(array_17_io_q),
    .io_r(array_17_io_r),
    .io_e_i(array_17_io_e_i),
    .io_f_i(array_17_io_f_i),
    .io_ve_i(array_17_io_ve_i),
    .io_vf_i(array_17_io_vf_i),
    .io_vv_i(array_17_io_vv_i),
    .io_e_o(array_17_io_e_o),
    .io_f_o(array_17_io_f_o),
    .io_v_o(array_17_io_v_o)
  );
  SWCell array_18 ( // @[SWChisel.scala 170:39]
    .io_q(array_18_io_q),
    .io_r(array_18_io_r),
    .io_e_i(array_18_io_e_i),
    .io_f_i(array_18_io_f_i),
    .io_ve_i(array_18_io_ve_i),
    .io_vf_i(array_18_io_vf_i),
    .io_vv_i(array_18_io_vv_i),
    .io_e_o(array_18_io_e_o),
    .io_f_o(array_18_io_f_o),
    .io_v_o(array_18_io_v_o)
  );
  SWCell array_19 ( // @[SWChisel.scala 170:39]
    .io_q(array_19_io_q),
    .io_r(array_19_io_r),
    .io_e_i(array_19_io_e_i),
    .io_f_i(array_19_io_f_i),
    .io_ve_i(array_19_io_ve_i),
    .io_vf_i(array_19_io_vf_i),
    .io_vv_i(array_19_io_vv_i),
    .io_e_o(array_19_io_e_o),
    .io_f_o(array_19_io_f_o),
    .io_v_o(array_19_io_v_o)
  );
  SWCell array_20 ( // @[SWChisel.scala 170:39]
    .io_q(array_20_io_q),
    .io_r(array_20_io_r),
    .io_e_i(array_20_io_e_i),
    .io_f_i(array_20_io_f_i),
    .io_ve_i(array_20_io_ve_i),
    .io_vf_i(array_20_io_vf_i),
    .io_vv_i(array_20_io_vv_i),
    .io_e_o(array_20_io_e_o),
    .io_f_o(array_20_io_f_o),
    .io_v_o(array_20_io_v_o)
  );
  SWCell array_21 ( // @[SWChisel.scala 170:39]
    .io_q(array_21_io_q),
    .io_r(array_21_io_r),
    .io_e_i(array_21_io_e_i),
    .io_f_i(array_21_io_f_i),
    .io_ve_i(array_21_io_ve_i),
    .io_vf_i(array_21_io_vf_i),
    .io_vv_i(array_21_io_vv_i),
    .io_e_o(array_21_io_e_o),
    .io_f_o(array_21_io_f_o),
    .io_v_o(array_21_io_v_o)
  );
  SWCell array_22 ( // @[SWChisel.scala 170:39]
    .io_q(array_22_io_q),
    .io_r(array_22_io_r),
    .io_e_i(array_22_io_e_i),
    .io_f_i(array_22_io_f_i),
    .io_ve_i(array_22_io_ve_i),
    .io_vf_i(array_22_io_vf_i),
    .io_vv_i(array_22_io_vv_i),
    .io_e_o(array_22_io_e_o),
    .io_f_o(array_22_io_f_o),
    .io_v_o(array_22_io_v_o)
  );
  SWCell array_23 ( // @[SWChisel.scala 170:39]
    .io_q(array_23_io_q),
    .io_r(array_23_io_r),
    .io_e_i(array_23_io_e_i),
    .io_f_i(array_23_io_f_i),
    .io_ve_i(array_23_io_ve_i),
    .io_vf_i(array_23_io_vf_i),
    .io_vv_i(array_23_io_vv_i),
    .io_e_o(array_23_io_e_o),
    .io_f_o(array_23_io_f_o),
    .io_v_o(array_23_io_v_o)
  );
  SWCell array_24 ( // @[SWChisel.scala 170:39]
    .io_q(array_24_io_q),
    .io_r(array_24_io_r),
    .io_e_i(array_24_io_e_i),
    .io_f_i(array_24_io_f_i),
    .io_ve_i(array_24_io_ve_i),
    .io_vf_i(array_24_io_vf_i),
    .io_vv_i(array_24_io_vv_i),
    .io_e_o(array_24_io_e_o),
    .io_f_o(array_24_io_f_o),
    .io_v_o(array_24_io_v_o)
  );
  SWCell array_25 ( // @[SWChisel.scala 170:39]
    .io_q(array_25_io_q),
    .io_r(array_25_io_r),
    .io_e_i(array_25_io_e_i),
    .io_f_i(array_25_io_f_i),
    .io_ve_i(array_25_io_ve_i),
    .io_vf_i(array_25_io_vf_i),
    .io_vv_i(array_25_io_vv_i),
    .io_e_o(array_25_io_e_o),
    .io_f_o(array_25_io_f_o),
    .io_v_o(array_25_io_v_o)
  );
  SWCell array_26 ( // @[SWChisel.scala 170:39]
    .io_q(array_26_io_q),
    .io_r(array_26_io_r),
    .io_e_i(array_26_io_e_i),
    .io_f_i(array_26_io_f_i),
    .io_ve_i(array_26_io_ve_i),
    .io_vf_i(array_26_io_vf_i),
    .io_vv_i(array_26_io_vv_i),
    .io_e_o(array_26_io_e_o),
    .io_f_o(array_26_io_f_o),
    .io_v_o(array_26_io_v_o)
  );
  SWCell array_27 ( // @[SWChisel.scala 170:39]
    .io_q(array_27_io_q),
    .io_r(array_27_io_r),
    .io_e_i(array_27_io_e_i),
    .io_f_i(array_27_io_f_i),
    .io_ve_i(array_27_io_ve_i),
    .io_vf_i(array_27_io_vf_i),
    .io_vv_i(array_27_io_vv_i),
    .io_e_o(array_27_io_e_o),
    .io_f_o(array_27_io_f_o),
    .io_v_o(array_27_io_v_o)
  );
  SWCell array_28 ( // @[SWChisel.scala 170:39]
    .io_q(array_28_io_q),
    .io_r(array_28_io_r),
    .io_e_i(array_28_io_e_i),
    .io_f_i(array_28_io_f_i),
    .io_ve_i(array_28_io_ve_i),
    .io_vf_i(array_28_io_vf_i),
    .io_vv_i(array_28_io_vv_i),
    .io_e_o(array_28_io_e_o),
    .io_f_o(array_28_io_f_o),
    .io_v_o(array_28_io_v_o)
  );
  SWCell array_29 ( // @[SWChisel.scala 170:39]
    .io_q(array_29_io_q),
    .io_r(array_29_io_r),
    .io_e_i(array_29_io_e_i),
    .io_f_i(array_29_io_f_i),
    .io_ve_i(array_29_io_ve_i),
    .io_vf_i(array_29_io_vf_i),
    .io_vv_i(array_29_io_vv_i),
    .io_e_o(array_29_io_e_o),
    .io_f_o(array_29_io_f_o),
    .io_v_o(array_29_io_v_o)
  );
  MyCounter r_count_0 ( // @[SWChisel.scala 171:41]
    .clock(r_count_0_clock),
    .reset(r_count_0_reset),
    .io_en(r_count_0_io_en),
    .io_out(r_count_0_io_out)
  );
  MyCounter r_count_1 ( // @[SWChisel.scala 171:41]
    .clock(r_count_1_clock),
    .reset(r_count_1_reset),
    .io_en(r_count_1_io_en),
    .io_out(r_count_1_io_out)
  );
  MyCounter r_count_2 ( // @[SWChisel.scala 171:41]
    .clock(r_count_2_clock),
    .reset(r_count_2_reset),
    .io_en(r_count_2_io_en),
    .io_out(r_count_2_io_out)
  );
  MyCounter r_count_3 ( // @[SWChisel.scala 171:41]
    .clock(r_count_3_clock),
    .reset(r_count_3_reset),
    .io_en(r_count_3_io_en),
    .io_out(r_count_3_io_out)
  );
  MyCounter r_count_4 ( // @[SWChisel.scala 171:41]
    .clock(r_count_4_clock),
    .reset(r_count_4_reset),
    .io_en(r_count_4_io_en),
    .io_out(r_count_4_io_out)
  );
  MyCounter r_count_5 ( // @[SWChisel.scala 171:41]
    .clock(r_count_5_clock),
    .reset(r_count_5_reset),
    .io_en(r_count_5_io_en),
    .io_out(r_count_5_io_out)
  );
  MyCounter r_count_6 ( // @[SWChisel.scala 171:41]
    .clock(r_count_6_clock),
    .reset(r_count_6_reset),
    .io_en(r_count_6_io_en),
    .io_out(r_count_6_io_out)
  );
  MyCounter r_count_7 ( // @[SWChisel.scala 171:41]
    .clock(r_count_7_clock),
    .reset(r_count_7_reset),
    .io_en(r_count_7_io_en),
    .io_out(r_count_7_io_out)
  );
  MyCounter r_count_8 ( // @[SWChisel.scala 171:41]
    .clock(r_count_8_clock),
    .reset(r_count_8_reset),
    .io_en(r_count_8_io_en),
    .io_out(r_count_8_io_out)
  );
  MyCounter r_count_9 ( // @[SWChisel.scala 171:41]
    .clock(r_count_9_clock),
    .reset(r_count_9_reset),
    .io_en(r_count_9_io_en),
    .io_out(r_count_9_io_out)
  );
  MyCounter r_count_10 ( // @[SWChisel.scala 171:41]
    .clock(r_count_10_clock),
    .reset(r_count_10_reset),
    .io_en(r_count_10_io_en),
    .io_out(r_count_10_io_out)
  );
  MyCounter r_count_11 ( // @[SWChisel.scala 171:41]
    .clock(r_count_11_clock),
    .reset(r_count_11_reset),
    .io_en(r_count_11_io_en),
    .io_out(r_count_11_io_out)
  );
  MyCounter r_count_12 ( // @[SWChisel.scala 171:41]
    .clock(r_count_12_clock),
    .reset(r_count_12_reset),
    .io_en(r_count_12_io_en),
    .io_out(r_count_12_io_out)
  );
  MyCounter r_count_13 ( // @[SWChisel.scala 171:41]
    .clock(r_count_13_clock),
    .reset(r_count_13_reset),
    .io_en(r_count_13_io_en),
    .io_out(r_count_13_io_out)
  );
  MyCounter r_count_14 ( // @[SWChisel.scala 171:41]
    .clock(r_count_14_clock),
    .reset(r_count_14_reset),
    .io_en(r_count_14_io_en),
    .io_out(r_count_14_io_out)
  );
  MyCounter r_count_15 ( // @[SWChisel.scala 171:41]
    .clock(r_count_15_clock),
    .reset(r_count_15_reset),
    .io_en(r_count_15_io_en),
    .io_out(r_count_15_io_out)
  );
  MyCounter r_count_16 ( // @[SWChisel.scala 171:41]
    .clock(r_count_16_clock),
    .reset(r_count_16_reset),
    .io_en(r_count_16_io_en),
    .io_out(r_count_16_io_out)
  );
  MyCounter r_count_17 ( // @[SWChisel.scala 171:41]
    .clock(r_count_17_clock),
    .reset(r_count_17_reset),
    .io_en(r_count_17_io_en),
    .io_out(r_count_17_io_out)
  );
  MyCounter r_count_18 ( // @[SWChisel.scala 171:41]
    .clock(r_count_18_clock),
    .reset(r_count_18_reset),
    .io_en(r_count_18_io_en),
    .io_out(r_count_18_io_out)
  );
  MyCounter r_count_19 ( // @[SWChisel.scala 171:41]
    .clock(r_count_19_clock),
    .reset(r_count_19_reset),
    .io_en(r_count_19_io_en),
    .io_out(r_count_19_io_out)
  );
  MyCounter r_count_20 ( // @[SWChisel.scala 171:41]
    .clock(r_count_20_clock),
    .reset(r_count_20_reset),
    .io_en(r_count_20_io_en),
    .io_out(r_count_20_io_out)
  );
  MyCounter r_count_21 ( // @[SWChisel.scala 171:41]
    .clock(r_count_21_clock),
    .reset(r_count_21_reset),
    .io_en(r_count_21_io_en),
    .io_out(r_count_21_io_out)
  );
  MyCounter r_count_22 ( // @[SWChisel.scala 171:41]
    .clock(r_count_22_clock),
    .reset(r_count_22_reset),
    .io_en(r_count_22_io_en),
    .io_out(r_count_22_io_out)
  );
  MyCounter r_count_23 ( // @[SWChisel.scala 171:41]
    .clock(r_count_23_clock),
    .reset(r_count_23_reset),
    .io_en(r_count_23_io_en),
    .io_out(r_count_23_io_out)
  );
  MyCounter r_count_24 ( // @[SWChisel.scala 171:41]
    .clock(r_count_24_clock),
    .reset(r_count_24_reset),
    .io_en(r_count_24_io_en),
    .io_out(r_count_24_io_out)
  );
  MyCounter r_count_25 ( // @[SWChisel.scala 171:41]
    .clock(r_count_25_clock),
    .reset(r_count_25_reset),
    .io_en(r_count_25_io_en),
    .io_out(r_count_25_io_out)
  );
  MyCounter r_count_26 ( // @[SWChisel.scala 171:41]
    .clock(r_count_26_clock),
    .reset(r_count_26_reset),
    .io_en(r_count_26_io_en),
    .io_out(r_count_26_io_out)
  );
  MyCounter r_count_27 ( // @[SWChisel.scala 171:41]
    .clock(r_count_27_clock),
    .reset(r_count_27_reset),
    .io_en(r_count_27_io_en),
    .io_out(r_count_27_io_out)
  );
  MyCounter r_count_28 ( // @[SWChisel.scala 171:41]
    .clock(r_count_28_clock),
    .reset(r_count_28_reset),
    .io_en(r_count_28_io_en),
    .io_out(r_count_28_io_out)
  );
  MyCounter r_count_29 ( // @[SWChisel.scala 171:41]
    .clock(r_count_29_clock),
    .reset(r_count_29_reset),
    .io_en(r_count_29_io_en),
    .io_out(r_count_29_io_out)
  );
  MAX max ( // @[SWChisel.scala 174:19]
    .clock(max_clock),
    .reset(max_reset),
    .io_start(max_io_start),
    .io_in(max_io_in),
    .io_done(max_io_done),
    .io_out(max_io_out)
  );
  assign io_result = max_io_out; // @[SWChisel.scala 181:13]
  assign io_done = max_io_done; // @[SWChisel.scala 182:11]
  assign array_0_io_q = io_q_0_b; // @[SWChisel.scala 220:19]
  assign array_0_io_r = 9'h12b == r_count_0_io_out ? io_r_299_b : _GEN_388; // @[SWChisel.scala 221:{19,19}]
  assign array_0_io_e_i = E_0; // @[SWChisel.scala 196:21]
  assign array_0_io_f_i = 16'sh0; // @[SWChisel.scala 198:21]
  assign array_0_io_ve_i = V1_1; // @[SWChisel.scala 197:22]
  assign array_0_io_vf_i = V1_0; // @[SWChisel.scala 199:22]
  assign array_0_io_vv_i = V2_0; // @[SWChisel.scala 200:22]
  assign array_1_io_q = io_q_1_b; // @[SWChisel.scala 220:19]
  assign array_1_io_r = 9'h12b == r_count_1_io_out ? io_r_299_b : _GEN_688; // @[SWChisel.scala 221:{19,19}]
  assign array_1_io_e_i = E_1; // @[SWChisel.scala 196:21]
  assign array_1_io_f_i = F_1; // @[SWChisel.scala 198:21]
  assign array_1_io_ve_i = V1_2; // @[SWChisel.scala 197:22]
  assign array_1_io_vf_i = V1_1; // @[SWChisel.scala 199:22]
  assign array_1_io_vv_i = V2_1; // @[SWChisel.scala 200:22]
  assign array_2_io_q = io_q_2_b; // @[SWChisel.scala 220:19]
  assign array_2_io_r = 9'h12b == r_count_2_io_out ? io_r_299_b : _GEN_988; // @[SWChisel.scala 221:{19,19}]
  assign array_2_io_e_i = E_2; // @[SWChisel.scala 196:21]
  assign array_2_io_f_i = F_2; // @[SWChisel.scala 198:21]
  assign array_2_io_ve_i = V1_3; // @[SWChisel.scala 197:22]
  assign array_2_io_vf_i = V1_2; // @[SWChisel.scala 199:22]
  assign array_2_io_vv_i = V2_2; // @[SWChisel.scala 200:22]
  assign array_3_io_q = io_q_3_b; // @[SWChisel.scala 220:19]
  assign array_3_io_r = 9'h12b == r_count_3_io_out ? io_r_299_b : _GEN_1288; // @[SWChisel.scala 221:{19,19}]
  assign array_3_io_e_i = E_3; // @[SWChisel.scala 196:21]
  assign array_3_io_f_i = F_3; // @[SWChisel.scala 198:21]
  assign array_3_io_ve_i = V1_4; // @[SWChisel.scala 197:22]
  assign array_3_io_vf_i = V1_3; // @[SWChisel.scala 199:22]
  assign array_3_io_vv_i = V2_3; // @[SWChisel.scala 200:22]
  assign array_4_io_q = io_q_4_b; // @[SWChisel.scala 220:19]
  assign array_4_io_r = 9'h12b == r_count_4_io_out ? io_r_299_b : _GEN_1588; // @[SWChisel.scala 221:{19,19}]
  assign array_4_io_e_i = E_4; // @[SWChisel.scala 196:21]
  assign array_4_io_f_i = F_4; // @[SWChisel.scala 198:21]
  assign array_4_io_ve_i = V1_5; // @[SWChisel.scala 197:22]
  assign array_4_io_vf_i = V1_4; // @[SWChisel.scala 199:22]
  assign array_4_io_vv_i = V2_4; // @[SWChisel.scala 200:22]
  assign array_5_io_q = io_q_5_b; // @[SWChisel.scala 220:19]
  assign array_5_io_r = 9'h12b == r_count_5_io_out ? io_r_299_b : _GEN_1888; // @[SWChisel.scala 221:{19,19}]
  assign array_5_io_e_i = E_5; // @[SWChisel.scala 196:21]
  assign array_5_io_f_i = F_5; // @[SWChisel.scala 198:21]
  assign array_5_io_ve_i = V1_6; // @[SWChisel.scala 197:22]
  assign array_5_io_vf_i = V1_5; // @[SWChisel.scala 199:22]
  assign array_5_io_vv_i = V2_5; // @[SWChisel.scala 200:22]
  assign array_6_io_q = io_q_6_b; // @[SWChisel.scala 220:19]
  assign array_6_io_r = 9'h12b == r_count_6_io_out ? io_r_299_b : _GEN_2188; // @[SWChisel.scala 221:{19,19}]
  assign array_6_io_e_i = E_6; // @[SWChisel.scala 196:21]
  assign array_6_io_f_i = F_6; // @[SWChisel.scala 198:21]
  assign array_6_io_ve_i = V1_7; // @[SWChisel.scala 197:22]
  assign array_6_io_vf_i = V1_6; // @[SWChisel.scala 199:22]
  assign array_6_io_vv_i = V2_6; // @[SWChisel.scala 200:22]
  assign array_7_io_q = io_q_7_b; // @[SWChisel.scala 220:19]
  assign array_7_io_r = 9'h12b == r_count_7_io_out ? io_r_299_b : _GEN_2488; // @[SWChisel.scala 221:{19,19}]
  assign array_7_io_e_i = E_7; // @[SWChisel.scala 196:21]
  assign array_7_io_f_i = F_7; // @[SWChisel.scala 198:21]
  assign array_7_io_ve_i = V1_8; // @[SWChisel.scala 197:22]
  assign array_7_io_vf_i = V1_7; // @[SWChisel.scala 199:22]
  assign array_7_io_vv_i = V2_7; // @[SWChisel.scala 200:22]
  assign array_8_io_q = io_q_8_b; // @[SWChisel.scala 220:19]
  assign array_8_io_r = 9'h12b == r_count_8_io_out ? io_r_299_b : _GEN_2788; // @[SWChisel.scala 221:{19,19}]
  assign array_8_io_e_i = E_8; // @[SWChisel.scala 196:21]
  assign array_8_io_f_i = F_8; // @[SWChisel.scala 198:21]
  assign array_8_io_ve_i = V1_9; // @[SWChisel.scala 197:22]
  assign array_8_io_vf_i = V1_8; // @[SWChisel.scala 199:22]
  assign array_8_io_vv_i = V2_8; // @[SWChisel.scala 200:22]
  assign array_9_io_q = io_q_9_b; // @[SWChisel.scala 220:19]
  assign array_9_io_r = 9'h12b == r_count_9_io_out ? io_r_299_b : _GEN_3088; // @[SWChisel.scala 221:{19,19}]
  assign array_9_io_e_i = E_9; // @[SWChisel.scala 196:21]
  assign array_9_io_f_i = F_9; // @[SWChisel.scala 198:21]
  assign array_9_io_ve_i = V1_10; // @[SWChisel.scala 197:22]
  assign array_9_io_vf_i = V1_9; // @[SWChisel.scala 199:22]
  assign array_9_io_vv_i = V2_9; // @[SWChisel.scala 200:22]
  assign array_10_io_q = io_q_10_b; // @[SWChisel.scala 220:19]
  assign array_10_io_r = 9'h12b == r_count_10_io_out ? io_r_299_b : _GEN_3388; // @[SWChisel.scala 221:{19,19}]
  assign array_10_io_e_i = E_10; // @[SWChisel.scala 196:21]
  assign array_10_io_f_i = F_10; // @[SWChisel.scala 198:21]
  assign array_10_io_ve_i = V1_11; // @[SWChisel.scala 197:22]
  assign array_10_io_vf_i = V1_10; // @[SWChisel.scala 199:22]
  assign array_10_io_vv_i = V2_10; // @[SWChisel.scala 200:22]
  assign array_11_io_q = io_q_11_b; // @[SWChisel.scala 220:19]
  assign array_11_io_r = 9'h12b == r_count_11_io_out ? io_r_299_b : _GEN_3688; // @[SWChisel.scala 221:{19,19}]
  assign array_11_io_e_i = E_11; // @[SWChisel.scala 196:21]
  assign array_11_io_f_i = F_11; // @[SWChisel.scala 198:21]
  assign array_11_io_ve_i = V1_12; // @[SWChisel.scala 197:22]
  assign array_11_io_vf_i = V1_11; // @[SWChisel.scala 199:22]
  assign array_11_io_vv_i = V2_11; // @[SWChisel.scala 200:22]
  assign array_12_io_q = io_q_12_b; // @[SWChisel.scala 220:19]
  assign array_12_io_r = 9'h12b == r_count_12_io_out ? io_r_299_b : _GEN_3988; // @[SWChisel.scala 221:{19,19}]
  assign array_12_io_e_i = E_12; // @[SWChisel.scala 196:21]
  assign array_12_io_f_i = F_12; // @[SWChisel.scala 198:21]
  assign array_12_io_ve_i = V1_13; // @[SWChisel.scala 197:22]
  assign array_12_io_vf_i = V1_12; // @[SWChisel.scala 199:22]
  assign array_12_io_vv_i = V2_12; // @[SWChisel.scala 200:22]
  assign array_13_io_q = io_q_13_b; // @[SWChisel.scala 220:19]
  assign array_13_io_r = 9'h12b == r_count_13_io_out ? io_r_299_b : _GEN_4288; // @[SWChisel.scala 221:{19,19}]
  assign array_13_io_e_i = E_13; // @[SWChisel.scala 196:21]
  assign array_13_io_f_i = F_13; // @[SWChisel.scala 198:21]
  assign array_13_io_ve_i = V1_14; // @[SWChisel.scala 197:22]
  assign array_13_io_vf_i = V1_13; // @[SWChisel.scala 199:22]
  assign array_13_io_vv_i = V2_13; // @[SWChisel.scala 200:22]
  assign array_14_io_q = io_q_14_b; // @[SWChisel.scala 220:19]
  assign array_14_io_r = 9'h12b == r_count_14_io_out ? io_r_299_b : _GEN_4588; // @[SWChisel.scala 221:{19,19}]
  assign array_14_io_e_i = E_14; // @[SWChisel.scala 196:21]
  assign array_14_io_f_i = F_14; // @[SWChisel.scala 198:21]
  assign array_14_io_ve_i = V1_15; // @[SWChisel.scala 197:22]
  assign array_14_io_vf_i = V1_14; // @[SWChisel.scala 199:22]
  assign array_14_io_vv_i = V2_14; // @[SWChisel.scala 200:22]
  assign array_15_io_q = io_q_15_b; // @[SWChisel.scala 220:19]
  assign array_15_io_r = 9'h12b == r_count_15_io_out ? io_r_299_b : _GEN_4888; // @[SWChisel.scala 221:{19,19}]
  assign array_15_io_e_i = E_15; // @[SWChisel.scala 196:21]
  assign array_15_io_f_i = F_15; // @[SWChisel.scala 198:21]
  assign array_15_io_ve_i = V1_16; // @[SWChisel.scala 197:22]
  assign array_15_io_vf_i = V1_15; // @[SWChisel.scala 199:22]
  assign array_15_io_vv_i = V2_15; // @[SWChisel.scala 200:22]
  assign array_16_io_q = io_q_16_b; // @[SWChisel.scala 220:19]
  assign array_16_io_r = 9'h12b == r_count_16_io_out ? io_r_299_b : _GEN_5188; // @[SWChisel.scala 221:{19,19}]
  assign array_16_io_e_i = E_16; // @[SWChisel.scala 196:21]
  assign array_16_io_f_i = F_16; // @[SWChisel.scala 198:21]
  assign array_16_io_ve_i = V1_17; // @[SWChisel.scala 197:22]
  assign array_16_io_vf_i = V1_16; // @[SWChisel.scala 199:22]
  assign array_16_io_vv_i = V2_16; // @[SWChisel.scala 200:22]
  assign array_17_io_q = io_q_17_b; // @[SWChisel.scala 220:19]
  assign array_17_io_r = 9'h12b == r_count_17_io_out ? io_r_299_b : _GEN_5488; // @[SWChisel.scala 221:{19,19}]
  assign array_17_io_e_i = E_17; // @[SWChisel.scala 196:21]
  assign array_17_io_f_i = F_17; // @[SWChisel.scala 198:21]
  assign array_17_io_ve_i = V1_18; // @[SWChisel.scala 197:22]
  assign array_17_io_vf_i = V1_17; // @[SWChisel.scala 199:22]
  assign array_17_io_vv_i = V2_17; // @[SWChisel.scala 200:22]
  assign array_18_io_q = io_q_18_b; // @[SWChisel.scala 220:19]
  assign array_18_io_r = 9'h12b == r_count_18_io_out ? io_r_299_b : _GEN_5788; // @[SWChisel.scala 221:{19,19}]
  assign array_18_io_e_i = E_18; // @[SWChisel.scala 196:21]
  assign array_18_io_f_i = F_18; // @[SWChisel.scala 198:21]
  assign array_18_io_ve_i = V1_19; // @[SWChisel.scala 197:22]
  assign array_18_io_vf_i = V1_18; // @[SWChisel.scala 199:22]
  assign array_18_io_vv_i = V2_18; // @[SWChisel.scala 200:22]
  assign array_19_io_q = io_q_19_b; // @[SWChisel.scala 220:19]
  assign array_19_io_r = 9'h12b == r_count_19_io_out ? io_r_299_b : _GEN_6088; // @[SWChisel.scala 221:{19,19}]
  assign array_19_io_e_i = E_19; // @[SWChisel.scala 196:21]
  assign array_19_io_f_i = F_19; // @[SWChisel.scala 198:21]
  assign array_19_io_ve_i = V1_20; // @[SWChisel.scala 197:22]
  assign array_19_io_vf_i = V1_19; // @[SWChisel.scala 199:22]
  assign array_19_io_vv_i = V2_19; // @[SWChisel.scala 200:22]
  assign array_20_io_q = io_q_20_b; // @[SWChisel.scala 220:19]
  assign array_20_io_r = 9'h12b == r_count_20_io_out ? io_r_299_b : _GEN_6388; // @[SWChisel.scala 221:{19,19}]
  assign array_20_io_e_i = E_20; // @[SWChisel.scala 196:21]
  assign array_20_io_f_i = F_20; // @[SWChisel.scala 198:21]
  assign array_20_io_ve_i = V1_21; // @[SWChisel.scala 197:22]
  assign array_20_io_vf_i = V1_20; // @[SWChisel.scala 199:22]
  assign array_20_io_vv_i = V2_20; // @[SWChisel.scala 200:22]
  assign array_21_io_q = io_q_21_b; // @[SWChisel.scala 220:19]
  assign array_21_io_r = 9'h12b == r_count_21_io_out ? io_r_299_b : _GEN_6688; // @[SWChisel.scala 221:{19,19}]
  assign array_21_io_e_i = E_21; // @[SWChisel.scala 196:21]
  assign array_21_io_f_i = F_21; // @[SWChisel.scala 198:21]
  assign array_21_io_ve_i = V1_22; // @[SWChisel.scala 197:22]
  assign array_21_io_vf_i = V1_21; // @[SWChisel.scala 199:22]
  assign array_21_io_vv_i = V2_21; // @[SWChisel.scala 200:22]
  assign array_22_io_q = io_q_22_b; // @[SWChisel.scala 220:19]
  assign array_22_io_r = 9'h12b == r_count_22_io_out ? io_r_299_b : _GEN_6988; // @[SWChisel.scala 221:{19,19}]
  assign array_22_io_e_i = E_22; // @[SWChisel.scala 196:21]
  assign array_22_io_f_i = F_22; // @[SWChisel.scala 198:21]
  assign array_22_io_ve_i = V1_23; // @[SWChisel.scala 197:22]
  assign array_22_io_vf_i = V1_22; // @[SWChisel.scala 199:22]
  assign array_22_io_vv_i = V2_22; // @[SWChisel.scala 200:22]
  assign array_23_io_q = io_q_23_b; // @[SWChisel.scala 220:19]
  assign array_23_io_r = 9'h12b == r_count_23_io_out ? io_r_299_b : _GEN_7288; // @[SWChisel.scala 221:{19,19}]
  assign array_23_io_e_i = E_23; // @[SWChisel.scala 196:21]
  assign array_23_io_f_i = F_23; // @[SWChisel.scala 198:21]
  assign array_23_io_ve_i = V1_24; // @[SWChisel.scala 197:22]
  assign array_23_io_vf_i = V1_23; // @[SWChisel.scala 199:22]
  assign array_23_io_vv_i = V2_23; // @[SWChisel.scala 200:22]
  assign array_24_io_q = io_q_24_b; // @[SWChisel.scala 220:19]
  assign array_24_io_r = 9'h12b == r_count_24_io_out ? io_r_299_b : _GEN_7588; // @[SWChisel.scala 221:{19,19}]
  assign array_24_io_e_i = E_24; // @[SWChisel.scala 196:21]
  assign array_24_io_f_i = F_24; // @[SWChisel.scala 198:21]
  assign array_24_io_ve_i = V1_25; // @[SWChisel.scala 197:22]
  assign array_24_io_vf_i = V1_24; // @[SWChisel.scala 199:22]
  assign array_24_io_vv_i = V2_24; // @[SWChisel.scala 200:22]
  assign array_25_io_q = io_q_25_b; // @[SWChisel.scala 220:19]
  assign array_25_io_r = 9'h12b == r_count_25_io_out ? io_r_299_b : _GEN_7888; // @[SWChisel.scala 221:{19,19}]
  assign array_25_io_e_i = E_25; // @[SWChisel.scala 196:21]
  assign array_25_io_f_i = F_25; // @[SWChisel.scala 198:21]
  assign array_25_io_ve_i = V1_26; // @[SWChisel.scala 197:22]
  assign array_25_io_vf_i = V1_25; // @[SWChisel.scala 199:22]
  assign array_25_io_vv_i = V2_25; // @[SWChisel.scala 200:22]
  assign array_26_io_q = io_q_26_b; // @[SWChisel.scala 220:19]
  assign array_26_io_r = 9'h12b == r_count_26_io_out ? io_r_299_b : _GEN_8188; // @[SWChisel.scala 221:{19,19}]
  assign array_26_io_e_i = E_26; // @[SWChisel.scala 196:21]
  assign array_26_io_f_i = F_26; // @[SWChisel.scala 198:21]
  assign array_26_io_ve_i = V1_27; // @[SWChisel.scala 197:22]
  assign array_26_io_vf_i = V1_26; // @[SWChisel.scala 199:22]
  assign array_26_io_vv_i = V2_26; // @[SWChisel.scala 200:22]
  assign array_27_io_q = io_q_27_b; // @[SWChisel.scala 220:19]
  assign array_27_io_r = 9'h12b == r_count_27_io_out ? io_r_299_b : _GEN_8488; // @[SWChisel.scala 221:{19,19}]
  assign array_27_io_e_i = E_27; // @[SWChisel.scala 196:21]
  assign array_27_io_f_i = F_27; // @[SWChisel.scala 198:21]
  assign array_27_io_ve_i = V1_28; // @[SWChisel.scala 197:22]
  assign array_27_io_vf_i = V1_27; // @[SWChisel.scala 199:22]
  assign array_27_io_vv_i = V2_27; // @[SWChisel.scala 200:22]
  assign array_28_io_q = io_q_28_b; // @[SWChisel.scala 220:19]
  assign array_28_io_r = 9'h12b == r_count_28_io_out ? io_r_299_b : _GEN_8788; // @[SWChisel.scala 221:{19,19}]
  assign array_28_io_e_i = E_28; // @[SWChisel.scala 196:21]
  assign array_28_io_f_i = F_28; // @[SWChisel.scala 198:21]
  assign array_28_io_ve_i = V1_29; // @[SWChisel.scala 197:22]
  assign array_28_io_vf_i = V1_28; // @[SWChisel.scala 199:22]
  assign array_28_io_vv_i = V2_28; // @[SWChisel.scala 200:22]
  assign array_29_io_q = io_q_29_b; // @[SWChisel.scala 220:19]
  assign array_29_io_r = 9'h12b == r_count_29_io_out ? io_r_299_b : _GEN_9088; // @[SWChisel.scala 221:{19,19}]
  assign array_29_io_e_i = E_29; // @[SWChisel.scala 196:21]
  assign array_29_io_f_i = F_29; // @[SWChisel.scala 198:21]
  assign array_29_io_ve_i = V1_30; // @[SWChisel.scala 197:22]
  assign array_29_io_vf_i = V1_29; // @[SWChisel.scala 199:22]
  assign array_29_io_vv_i = V2_29; // @[SWChisel.scala 200:22]
  assign r_count_0_clock = clock;
  assign r_count_0_reset = reset;
  assign r_count_0_io_en = start_reg_0; // @[SWChisel.scala 192:22]
  assign r_count_1_clock = clock;
  assign r_count_1_reset = reset;
  assign r_count_1_io_en = start_reg_1; // @[SWChisel.scala 192:22]
  assign r_count_2_clock = clock;
  assign r_count_2_reset = reset;
  assign r_count_2_io_en = start_reg_2; // @[SWChisel.scala 192:22]
  assign r_count_3_clock = clock;
  assign r_count_3_reset = reset;
  assign r_count_3_io_en = start_reg_3; // @[SWChisel.scala 192:22]
  assign r_count_4_clock = clock;
  assign r_count_4_reset = reset;
  assign r_count_4_io_en = start_reg_4; // @[SWChisel.scala 192:22]
  assign r_count_5_clock = clock;
  assign r_count_5_reset = reset;
  assign r_count_5_io_en = start_reg_5; // @[SWChisel.scala 192:22]
  assign r_count_6_clock = clock;
  assign r_count_6_reset = reset;
  assign r_count_6_io_en = start_reg_6; // @[SWChisel.scala 192:22]
  assign r_count_7_clock = clock;
  assign r_count_7_reset = reset;
  assign r_count_7_io_en = start_reg_7; // @[SWChisel.scala 192:22]
  assign r_count_8_clock = clock;
  assign r_count_8_reset = reset;
  assign r_count_8_io_en = start_reg_8; // @[SWChisel.scala 192:22]
  assign r_count_9_clock = clock;
  assign r_count_9_reset = reset;
  assign r_count_9_io_en = start_reg_9; // @[SWChisel.scala 192:22]
  assign r_count_10_clock = clock;
  assign r_count_10_reset = reset;
  assign r_count_10_io_en = start_reg_10; // @[SWChisel.scala 192:22]
  assign r_count_11_clock = clock;
  assign r_count_11_reset = reset;
  assign r_count_11_io_en = start_reg_11; // @[SWChisel.scala 192:22]
  assign r_count_12_clock = clock;
  assign r_count_12_reset = reset;
  assign r_count_12_io_en = start_reg_12; // @[SWChisel.scala 192:22]
  assign r_count_13_clock = clock;
  assign r_count_13_reset = reset;
  assign r_count_13_io_en = start_reg_13; // @[SWChisel.scala 192:22]
  assign r_count_14_clock = clock;
  assign r_count_14_reset = reset;
  assign r_count_14_io_en = start_reg_14; // @[SWChisel.scala 192:22]
  assign r_count_15_clock = clock;
  assign r_count_15_reset = reset;
  assign r_count_15_io_en = start_reg_15; // @[SWChisel.scala 192:22]
  assign r_count_16_clock = clock;
  assign r_count_16_reset = reset;
  assign r_count_16_io_en = start_reg_16; // @[SWChisel.scala 192:22]
  assign r_count_17_clock = clock;
  assign r_count_17_reset = reset;
  assign r_count_17_io_en = start_reg_17; // @[SWChisel.scala 192:22]
  assign r_count_18_clock = clock;
  assign r_count_18_reset = reset;
  assign r_count_18_io_en = start_reg_18; // @[SWChisel.scala 192:22]
  assign r_count_19_clock = clock;
  assign r_count_19_reset = reset;
  assign r_count_19_io_en = start_reg_19; // @[SWChisel.scala 192:22]
  assign r_count_20_clock = clock;
  assign r_count_20_reset = reset;
  assign r_count_20_io_en = start_reg_20; // @[SWChisel.scala 192:22]
  assign r_count_21_clock = clock;
  assign r_count_21_reset = reset;
  assign r_count_21_io_en = start_reg_21; // @[SWChisel.scala 192:22]
  assign r_count_22_clock = clock;
  assign r_count_22_reset = reset;
  assign r_count_22_io_en = start_reg_22; // @[SWChisel.scala 192:22]
  assign r_count_23_clock = clock;
  assign r_count_23_reset = reset;
  assign r_count_23_io_en = start_reg_23; // @[SWChisel.scala 192:22]
  assign r_count_24_clock = clock;
  assign r_count_24_reset = reset;
  assign r_count_24_io_en = start_reg_24; // @[SWChisel.scala 192:22]
  assign r_count_25_clock = clock;
  assign r_count_25_reset = reset;
  assign r_count_25_io_en = start_reg_25; // @[SWChisel.scala 192:22]
  assign r_count_26_clock = clock;
  assign r_count_26_reset = reset;
  assign r_count_26_io_en = start_reg_26; // @[SWChisel.scala 192:22]
  assign r_count_27_clock = clock;
  assign r_count_27_reset = reset;
  assign r_count_27_io_en = start_reg_27; // @[SWChisel.scala 192:22]
  assign r_count_28_clock = clock;
  assign r_count_28_reset = reset;
  assign r_count_28_io_en = start_reg_28; // @[SWChisel.scala 192:22]
  assign r_count_29_clock = clock;
  assign r_count_29_reset = reset;
  assign r_count_29_io_en = start_reg_29; // @[SWChisel.scala 192:22]
  assign max_clock = clock;
  assign max_reset = reset;
  assign max_io_start = start_reg_29; // @[SWChisel.scala 178:16]
  assign max_io_in = V1_30; // @[SWChisel.scala 177:13]
  always @(posedge clock) begin
    if (reset) begin // @[SWChisel.scala 162:18]
      E_0 <= -16'sh2; // @[SWChisel.scala 162:18]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      E_0 <= array_0_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_1 <= -16'sh3; // @[SWChisel.scala 162:18]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      E_1 <= array_1_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_2 <= -16'sh4; // @[SWChisel.scala 162:18]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      E_2 <= array_2_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_3 <= -16'sh5; // @[SWChisel.scala 162:18]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      E_3 <= array_3_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_4 <= -16'sh6; // @[SWChisel.scala 162:18]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      E_4 <= array_4_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_5 <= -16'sh7; // @[SWChisel.scala 162:18]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      E_5 <= array_5_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_6 <= -16'sh8; // @[SWChisel.scala 162:18]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      E_6 <= array_6_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_7 <= -16'sh9; // @[SWChisel.scala 162:18]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      E_7 <= array_7_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_8 <= -16'sha; // @[SWChisel.scala 162:18]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      E_8 <= array_8_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_9 <= -16'shb; // @[SWChisel.scala 162:18]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      E_9 <= array_9_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_10 <= -16'shc; // @[SWChisel.scala 162:18]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      E_10 <= array_10_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_11 <= -16'shd; // @[SWChisel.scala 162:18]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      E_11 <= array_11_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_12 <= -16'she; // @[SWChisel.scala 162:18]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      E_12 <= array_12_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_13 <= -16'shf; // @[SWChisel.scala 162:18]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      E_13 <= array_13_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_14 <= -16'sh10; // @[SWChisel.scala 162:18]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      E_14 <= array_14_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_15 <= -16'sh11; // @[SWChisel.scala 162:18]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      E_15 <= array_15_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_16 <= -16'sh12; // @[SWChisel.scala 162:18]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      E_16 <= array_16_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_17 <= -16'sh13; // @[SWChisel.scala 162:18]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      E_17 <= array_17_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_18 <= -16'sh14; // @[SWChisel.scala 162:18]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      E_18 <= array_18_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_19 <= -16'sh15; // @[SWChisel.scala 162:18]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      E_19 <= array_19_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_20 <= -16'sh16; // @[SWChisel.scala 162:18]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      E_20 <= array_20_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_21 <= -16'sh17; // @[SWChisel.scala 162:18]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      E_21 <= array_21_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_22 <= -16'sh18; // @[SWChisel.scala 162:18]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      E_22 <= array_22_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_23 <= -16'sh19; // @[SWChisel.scala 162:18]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      E_23 <= array_23_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_24 <= -16'sh1a; // @[SWChisel.scala 162:18]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      E_24 <= array_24_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_25 <= -16'sh1b; // @[SWChisel.scala 162:18]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      E_25 <= array_25_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_26 <= -16'sh1c; // @[SWChisel.scala 162:18]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      E_26 <= array_26_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_27 <= -16'sh1d; // @[SWChisel.scala 162:18]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      E_27 <= array_27_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_28 <= -16'sh1e; // @[SWChisel.scala 162:18]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      E_28 <= array_28_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_29 <= -16'sh1f; // @[SWChisel.scala 162:18]
    end else if (start_reg_29) begin // @[SWChisel.scala 207:25]
      E_29 <= array_29_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_1 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      F_1 <= array_0_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_2 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      F_2 <= array_1_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_3 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      F_3 <= array_2_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_4 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      F_4 <= array_3_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_5 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      F_5 <= array_4_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_6 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      F_6 <= array_5_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_7 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      F_7 <= array_6_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_8 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      F_8 <= array_7_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_9 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      F_9 <= array_8_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_10 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      F_10 <= array_9_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_11 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      F_11 <= array_10_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_12 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      F_12 <= array_11_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_13 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      F_13 <= array_12_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_14 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      F_14 <= array_13_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_15 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      F_15 <= array_14_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_16 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      F_16 <= array_15_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_17 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      F_17 <= array_16_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_18 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      F_18 <= array_17_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_19 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      F_19 <= array_18_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_20 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      F_20 <= array_19_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_21 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      F_21 <= array_20_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_22 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      F_22 <= array_21_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_23 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      F_23 <= array_22_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_24 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      F_24 <= array_23_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_25 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      F_25 <= array_24_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_26 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      F_26 <= array_25_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_27 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      F_27 <= array_26_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_28 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      F_28 <= array_27_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_29 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      F_29 <= array_28_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_0 <= -16'sh1; // @[SWChisel.scala 164:19]
    end else begin
      V1_0 <= 16'sh0; // @[SWChisel.scala 165:9]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_1 <= -16'sh2; // @[SWChisel.scala 164:19]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      V1_1 <= array_0_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_2 <= -16'sh3; // @[SWChisel.scala 164:19]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      V1_2 <= array_1_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_3 <= -16'sh4; // @[SWChisel.scala 164:19]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      V1_3 <= array_2_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_4 <= -16'sh5; // @[SWChisel.scala 164:19]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      V1_4 <= array_3_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_5 <= -16'sh6; // @[SWChisel.scala 164:19]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      V1_5 <= array_4_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_6 <= -16'sh7; // @[SWChisel.scala 164:19]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      V1_6 <= array_5_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_7 <= -16'sh8; // @[SWChisel.scala 164:19]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      V1_7 <= array_6_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_8 <= -16'sh9; // @[SWChisel.scala 164:19]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      V1_8 <= array_7_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_9 <= -16'sha; // @[SWChisel.scala 164:19]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      V1_9 <= array_8_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_10 <= -16'shb; // @[SWChisel.scala 164:19]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      V1_10 <= array_9_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_11 <= -16'shc; // @[SWChisel.scala 164:19]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      V1_11 <= array_10_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_12 <= -16'shd; // @[SWChisel.scala 164:19]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      V1_12 <= array_11_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_13 <= -16'she; // @[SWChisel.scala 164:19]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      V1_13 <= array_12_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_14 <= -16'shf; // @[SWChisel.scala 164:19]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      V1_14 <= array_13_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_15 <= -16'sh10; // @[SWChisel.scala 164:19]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      V1_15 <= array_14_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_16 <= -16'sh11; // @[SWChisel.scala 164:19]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      V1_16 <= array_15_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_17 <= -16'sh12; // @[SWChisel.scala 164:19]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      V1_17 <= array_16_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_18 <= -16'sh13; // @[SWChisel.scala 164:19]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      V1_18 <= array_17_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_19 <= -16'sh14; // @[SWChisel.scala 164:19]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      V1_19 <= array_18_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_20 <= -16'sh15; // @[SWChisel.scala 164:19]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      V1_20 <= array_19_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_21 <= -16'sh16; // @[SWChisel.scala 164:19]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      V1_21 <= array_20_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_22 <= -16'sh17; // @[SWChisel.scala 164:19]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      V1_22 <= array_21_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_23 <= -16'sh18; // @[SWChisel.scala 164:19]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      V1_23 <= array_22_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_24 <= -16'sh19; // @[SWChisel.scala 164:19]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      V1_24 <= array_23_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_25 <= -16'sh1a; // @[SWChisel.scala 164:19]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      V1_25 <= array_24_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_26 <= -16'sh1b; // @[SWChisel.scala 164:19]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      V1_26 <= array_25_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_27 <= -16'sh1c; // @[SWChisel.scala 164:19]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      V1_27 <= array_26_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_28 <= -16'sh1d; // @[SWChisel.scala 164:19]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      V1_28 <= array_27_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_29 <= -16'sh1e; // @[SWChisel.scala 164:19]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      V1_29 <= array_28_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_30 <= -16'sh1f; // @[SWChisel.scala 164:19]
    end else if (start_reg_29) begin // @[SWChisel.scala 207:25]
      V1_30 <= array_29_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_0 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_0 <= V1_0; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_1 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_1 <= V1_1; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_2 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_2 <= V1_2; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_3 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_3 <= V1_3; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_4 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_4 <= V1_4; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_5 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_5 <= V1_5; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_6 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_6 <= V1_6; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_7 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_7 <= V1_7; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_8 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_8 <= V1_8; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_9 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_9 <= V1_9; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_10 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_10 <= V1_10; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_11 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_11 <= V1_11; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_12 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_12 <= V1_12; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_13 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_13 <= V1_13; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_14 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_14 <= V1_14; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_15 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_15 <= V1_15; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_16 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_16 <= V1_16; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_17 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_17 <= V1_17; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_18 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_18 <= V1_18; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_19 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_19 <= V1_19; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_20 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_20 <= V1_20; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_21 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_21 <= V1_21; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_22 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_22 <= V1_22; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_23 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_23 <= V1_23; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_24 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_24 <= V1_24; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_25 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_25 <= V1_25; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_26 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_26 <= V1_26; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_27 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_27 <= V1_27; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_28 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_28 <= V1_28; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_29 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_29 <= V1_29; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_0 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_0 <= io_start; // @[SWChisel.scala 185:16]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_1 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_1 <= start_reg_0; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_2 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_2 <= start_reg_1; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_3 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_3 <= start_reg_2; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_4 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_4 <= start_reg_3; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_5 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_5 <= start_reg_4; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_6 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_6 <= start_reg_5; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_7 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_7 <= start_reg_6; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_8 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_8 <= start_reg_7; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_9 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_9 <= start_reg_8; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_10 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_10 <= start_reg_9; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_11 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_11 <= start_reg_10; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_12 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_12 <= start_reg_11; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_13 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_13 <= start_reg_12; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_14 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_14 <= start_reg_13; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_15 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_15 <= start_reg_14; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_16 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_16 <= start_reg_15; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_17 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_17 <= start_reg_16; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_18 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_18 <= start_reg_17; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_19 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_19 <= start_reg_18; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_20 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_20 <= start_reg_19; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_21 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_21 <= start_reg_20; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_22 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_22 <= start_reg_21; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_23 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_23 <= start_reg_22; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_24 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_24 <= start_reg_23; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_25 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_25 <= start_reg_24; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_26 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_26 <= start_reg_25; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_27 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_27 <= start_reg_26; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_28 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_28 <= start_reg_27; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_29 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_29 <= start_reg_28; // @[SWChisel.scala 187:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  E_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  E_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  E_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  E_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  E_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  E_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  E_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  E_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  E_8 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  E_9 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  E_10 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  E_11 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  E_12 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  E_13 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  E_14 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  E_15 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  E_16 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  E_17 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  E_18 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  E_19 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  E_20 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  E_21 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  E_22 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  E_23 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  E_24 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  E_25 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  E_26 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  E_27 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  E_28 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  E_29 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  F_1 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  F_2 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  F_3 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  F_4 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  F_5 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  F_6 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  F_7 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  F_8 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  F_9 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  F_10 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  F_11 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  F_12 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  F_13 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  F_14 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  F_15 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  F_16 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  F_17 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  F_18 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  F_19 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  F_20 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  F_21 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  F_22 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  F_23 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  F_24 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  F_25 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  F_26 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  F_27 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  F_28 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  F_29 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  V1_0 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  V1_1 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  V1_2 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  V1_3 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  V1_4 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  V1_5 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  V1_6 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  V1_7 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  V1_8 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  V1_9 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  V1_10 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  V1_11 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  V1_12 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  V1_13 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  V1_14 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  V1_15 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  V1_16 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  V1_17 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  V1_18 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  V1_19 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  V1_20 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  V1_21 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  V1_22 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  V1_23 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  V1_24 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  V1_25 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  V1_26 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  V1_27 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  V1_28 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  V1_29 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  V1_30 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  V2_0 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  V2_1 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  V2_2 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  V2_3 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  V2_4 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  V2_5 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  V2_6 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  V2_7 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  V2_8 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  V2_9 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  V2_10 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  V2_11 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  V2_12 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  V2_13 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  V2_14 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  V2_15 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  V2_16 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  V2_17 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  V2_18 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  V2_19 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  V2_20 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  V2_21 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  V2_22 = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  V2_23 = _RAND_113[15:0];
  _RAND_114 = {1{`RANDOM}};
  V2_24 = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  V2_25 = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  V2_26 = _RAND_116[15:0];
  _RAND_117 = {1{`RANDOM}};
  V2_27 = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  V2_28 = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  V2_29 = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  start_reg_0 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  start_reg_1 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  start_reg_2 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  start_reg_3 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  start_reg_4 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  start_reg_5 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  start_reg_6 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  start_reg_7 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  start_reg_8 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  start_reg_9 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  start_reg_10 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  start_reg_11 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  start_reg_12 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  start_reg_13 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  start_reg_14 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  start_reg_15 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  start_reg_16 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  start_reg_17 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  start_reg_18 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  start_reg_19 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  start_reg_20 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  start_reg_21 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  start_reg_22 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  start_reg_23 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  start_reg_24 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  start_reg_25 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  start_reg_26 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  start_reg_27 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  start_reg_28 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  start_reg_29 = _RAND_149[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
