module SWCell(
  input  [1:0]  io_q,
  input  [1:0]  io_r,
  input  [15:0] io_e_i,
  input  [15:0] io_f_i,
  input  [15:0] io_ve_i,
  input  [15:0] io_vf_i,
  input  [15:0] io_vv_i,
  output [15:0] io_e_o,
  output [15:0] io_f_o,
  output [15:0] io_v_o
);
  wire [15:0] _T_2 = $signed(io_ve_i) - 16'sh2; // @[SWChisel.scala 78:17]
  wire [15:0] _T_5 = $signed(io_e_i) - 16'sh1; // @[SWChisel.scala 78:39]
  wire [15:0] e_max = $signed(_T_2) >= $signed(_T_5) ? $signed(_T_2) : $signed(_T_5); // @[SWChisel.scala 78:51 79:11 81:11]
  wire [15:0] _T_9 = $signed(io_vf_i) - 16'sh2; // @[SWChisel.scala 85:17]
  wire [15:0] _T_12 = $signed(io_f_i) - 16'sh1; // @[SWChisel.scala 85:38]
  wire [15:0] f_max = $signed(_T_9) > $signed(_T_12) ? $signed(_T_9) : $signed(_T_12); // @[SWChisel.scala 85:50 86:11 88:11]
  wire [15:0] ef_temp = $signed(e_max) > $signed(f_max) ? $signed(e_max) : $signed(f_max); // @[SWChisel.scala 92:24 93:13 95:13]
  wire [15:0] _v_temp_T_2 = $signed(io_vv_i) + 16'sh2; // @[SWChisel.scala 100:23]
  wire [15:0] _v_temp_T_5 = $signed(io_vv_i) - 16'sh2; // @[SWChisel.scala 102:23]
  wire [15:0] v_temp = io_q == io_r ? $signed(_v_temp_T_2) : $signed(_v_temp_T_5); // @[SWChisel.scala 100:12 102:12 99:24]
  assign io_e_o = $signed(_T_2) >= $signed(_T_5) ? $signed(_T_2) : $signed(_T_5); // @[SWChisel.scala 78:51 79:11 81:11]
  assign io_f_o = $signed(_T_9) > $signed(_T_12) ? $signed(_T_9) : $signed(_T_12); // @[SWChisel.scala 85:50 86:11 88:11]
  assign io_v_o = $signed(v_temp) > $signed(ef_temp) ? $signed(v_temp) : $signed(ef_temp); // @[SWChisel.scala 106:27 107:11 109:11]
endmodule
module MyCounter(
  input        clock,
  input        reset,
  input        io_en,
  output [9:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [9:0] _io_out_T_2 = io_out + 10'h1; // @[SWChisel.scala 155:55]
  reg [9:0] io_out_r; // @[Reg.scala 35:20]
  assign io_out = io_out_r; // @[SWChisel.scala 155:12]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      io_out_r <= 10'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_out < 10'h2ee) begin // @[SWChisel.scala 155:28]
        io_out_r <= _io_out_T_2;
      end else begin
        io_out_r <= 10'h0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_out_r = _RAND_0[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MAX(
  input         clock,
  input         reset,
  input         io_start,
  input  [15:0] io_in,
  output        io_done,
  output [15:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] max; // @[SWChisel.scala 122:20]
  reg [9:0] counter; // @[SWChisel.scala 133:24]
  wire [9:0] _counter_T_1 = counter - 10'h1; // @[SWChisel.scala 135:24]
  assign io_done = counter == 10'h0; // @[SWChisel.scala 141:17]
  assign io_out = max; // @[SWChisel.scala 123:10]
  always @(posedge clock) begin
    if (reset) begin // @[SWChisel.scala 122:20]
      max <= 16'sh8000; // @[SWChisel.scala 122:20]
    end else if ($signed(io_in) > $signed(max)) begin // @[SWChisel.scala 126:22]
      max <= io_in; // @[SWChisel.scala 127:9]
    end
    if (reset) begin // @[SWChisel.scala 133:24]
      counter <= 10'h2ef; // @[SWChisel.scala 133:24]
    end else if (counter == 10'h0) begin // @[SWChisel.scala 141:26]
      counter <= 10'h0; // @[SWChisel.scala 143:13]
    end else if (io_start) begin // @[SWChisel.scala 134:19]
      counter <= _counter_T_1; // @[SWChisel.scala 135:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  max = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  counter = _RAND_1[9:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SW(
  input         clock,
  input         reset,
  input  [1:0]  io_q_0_b,
  input  [1:0]  io_q_1_b,
  input  [1:0]  io_q_2_b,
  input  [1:0]  io_q_3_b,
  input  [1:0]  io_q_4_b,
  input  [1:0]  io_q_5_b,
  input  [1:0]  io_q_6_b,
  input  [1:0]  io_q_7_b,
  input  [1:0]  io_q_8_b,
  input  [1:0]  io_q_9_b,
  input  [1:0]  io_q_10_b,
  input  [1:0]  io_q_11_b,
  input  [1:0]  io_q_12_b,
  input  [1:0]  io_q_13_b,
  input  [1:0]  io_q_14_b,
  input  [1:0]  io_q_15_b,
  input  [1:0]  io_q_16_b,
  input  [1:0]  io_q_17_b,
  input  [1:0]  io_q_18_b,
  input  [1:0]  io_q_19_b,
  input  [1:0]  io_q_20_b,
  input  [1:0]  io_q_21_b,
  input  [1:0]  io_q_22_b,
  input  [1:0]  io_q_23_b,
  input  [1:0]  io_q_24_b,
  input  [1:0]  io_q_25_b,
  input  [1:0]  io_q_26_b,
  input  [1:0]  io_q_27_b,
  input  [1:0]  io_q_28_b,
  input  [1:0]  io_q_29_b,
  input  [1:0]  io_r_0_b,
  input  [1:0]  io_r_1_b,
  input  [1:0]  io_r_2_b,
  input  [1:0]  io_r_3_b,
  input  [1:0]  io_r_4_b,
  input  [1:0]  io_r_5_b,
  input  [1:0]  io_r_6_b,
  input  [1:0]  io_r_7_b,
  input  [1:0]  io_r_8_b,
  input  [1:0]  io_r_9_b,
  input  [1:0]  io_r_10_b,
  input  [1:0]  io_r_11_b,
  input  [1:0]  io_r_12_b,
  input  [1:0]  io_r_13_b,
  input  [1:0]  io_r_14_b,
  input  [1:0]  io_r_15_b,
  input  [1:0]  io_r_16_b,
  input  [1:0]  io_r_17_b,
  input  [1:0]  io_r_18_b,
  input  [1:0]  io_r_19_b,
  input  [1:0]  io_r_20_b,
  input  [1:0]  io_r_21_b,
  input  [1:0]  io_r_22_b,
  input  [1:0]  io_r_23_b,
  input  [1:0]  io_r_24_b,
  input  [1:0]  io_r_25_b,
  input  [1:0]  io_r_26_b,
  input  [1:0]  io_r_27_b,
  input  [1:0]  io_r_28_b,
  input  [1:0]  io_r_29_b,
  input  [1:0]  io_r_30_b,
  input  [1:0]  io_r_31_b,
  input  [1:0]  io_r_32_b,
  input  [1:0]  io_r_33_b,
  input  [1:0]  io_r_34_b,
  input  [1:0]  io_r_35_b,
  input  [1:0]  io_r_36_b,
  input  [1:0]  io_r_37_b,
  input  [1:0]  io_r_38_b,
  input  [1:0]  io_r_39_b,
  input  [1:0]  io_r_40_b,
  input  [1:0]  io_r_41_b,
  input  [1:0]  io_r_42_b,
  input  [1:0]  io_r_43_b,
  input  [1:0]  io_r_44_b,
  input  [1:0]  io_r_45_b,
  input  [1:0]  io_r_46_b,
  input  [1:0]  io_r_47_b,
  input  [1:0]  io_r_48_b,
  input  [1:0]  io_r_49_b,
  input  [1:0]  io_r_50_b,
  input  [1:0]  io_r_51_b,
  input  [1:0]  io_r_52_b,
  input  [1:0]  io_r_53_b,
  input  [1:0]  io_r_54_b,
  input  [1:0]  io_r_55_b,
  input  [1:0]  io_r_56_b,
  input  [1:0]  io_r_57_b,
  input  [1:0]  io_r_58_b,
  input  [1:0]  io_r_59_b,
  input  [1:0]  io_r_60_b,
  input  [1:0]  io_r_61_b,
  input  [1:0]  io_r_62_b,
  input  [1:0]  io_r_63_b,
  input  [1:0]  io_r_64_b,
  input  [1:0]  io_r_65_b,
  input  [1:0]  io_r_66_b,
  input  [1:0]  io_r_67_b,
  input  [1:0]  io_r_68_b,
  input  [1:0]  io_r_69_b,
  input  [1:0]  io_r_70_b,
  input  [1:0]  io_r_71_b,
  input  [1:0]  io_r_72_b,
  input  [1:0]  io_r_73_b,
  input  [1:0]  io_r_74_b,
  input  [1:0]  io_r_75_b,
  input  [1:0]  io_r_76_b,
  input  [1:0]  io_r_77_b,
  input  [1:0]  io_r_78_b,
  input  [1:0]  io_r_79_b,
  input  [1:0]  io_r_80_b,
  input  [1:0]  io_r_81_b,
  input  [1:0]  io_r_82_b,
  input  [1:0]  io_r_83_b,
  input  [1:0]  io_r_84_b,
  input  [1:0]  io_r_85_b,
  input  [1:0]  io_r_86_b,
  input  [1:0]  io_r_87_b,
  input  [1:0]  io_r_88_b,
  input  [1:0]  io_r_89_b,
  input  [1:0]  io_r_90_b,
  input  [1:0]  io_r_91_b,
  input  [1:0]  io_r_92_b,
  input  [1:0]  io_r_93_b,
  input  [1:0]  io_r_94_b,
  input  [1:0]  io_r_95_b,
  input  [1:0]  io_r_96_b,
  input  [1:0]  io_r_97_b,
  input  [1:0]  io_r_98_b,
  input  [1:0]  io_r_99_b,
  input  [1:0]  io_r_100_b,
  input  [1:0]  io_r_101_b,
  input  [1:0]  io_r_102_b,
  input  [1:0]  io_r_103_b,
  input  [1:0]  io_r_104_b,
  input  [1:0]  io_r_105_b,
  input  [1:0]  io_r_106_b,
  input  [1:0]  io_r_107_b,
  input  [1:0]  io_r_108_b,
  input  [1:0]  io_r_109_b,
  input  [1:0]  io_r_110_b,
  input  [1:0]  io_r_111_b,
  input  [1:0]  io_r_112_b,
  input  [1:0]  io_r_113_b,
  input  [1:0]  io_r_114_b,
  input  [1:0]  io_r_115_b,
  input  [1:0]  io_r_116_b,
  input  [1:0]  io_r_117_b,
  input  [1:0]  io_r_118_b,
  input  [1:0]  io_r_119_b,
  input  [1:0]  io_r_120_b,
  input  [1:0]  io_r_121_b,
  input  [1:0]  io_r_122_b,
  input  [1:0]  io_r_123_b,
  input  [1:0]  io_r_124_b,
  input  [1:0]  io_r_125_b,
  input  [1:0]  io_r_126_b,
  input  [1:0]  io_r_127_b,
  input  [1:0]  io_r_128_b,
  input  [1:0]  io_r_129_b,
  input  [1:0]  io_r_130_b,
  input  [1:0]  io_r_131_b,
  input  [1:0]  io_r_132_b,
  input  [1:0]  io_r_133_b,
  input  [1:0]  io_r_134_b,
  input  [1:0]  io_r_135_b,
  input  [1:0]  io_r_136_b,
  input  [1:0]  io_r_137_b,
  input  [1:0]  io_r_138_b,
  input  [1:0]  io_r_139_b,
  input  [1:0]  io_r_140_b,
  input  [1:0]  io_r_141_b,
  input  [1:0]  io_r_142_b,
  input  [1:0]  io_r_143_b,
  input  [1:0]  io_r_144_b,
  input  [1:0]  io_r_145_b,
  input  [1:0]  io_r_146_b,
  input  [1:0]  io_r_147_b,
  input  [1:0]  io_r_148_b,
  input  [1:0]  io_r_149_b,
  input  [1:0]  io_r_150_b,
  input  [1:0]  io_r_151_b,
  input  [1:0]  io_r_152_b,
  input  [1:0]  io_r_153_b,
  input  [1:0]  io_r_154_b,
  input  [1:0]  io_r_155_b,
  input  [1:0]  io_r_156_b,
  input  [1:0]  io_r_157_b,
  input  [1:0]  io_r_158_b,
  input  [1:0]  io_r_159_b,
  input  [1:0]  io_r_160_b,
  input  [1:0]  io_r_161_b,
  input  [1:0]  io_r_162_b,
  input  [1:0]  io_r_163_b,
  input  [1:0]  io_r_164_b,
  input  [1:0]  io_r_165_b,
  input  [1:0]  io_r_166_b,
  input  [1:0]  io_r_167_b,
  input  [1:0]  io_r_168_b,
  input  [1:0]  io_r_169_b,
  input  [1:0]  io_r_170_b,
  input  [1:0]  io_r_171_b,
  input  [1:0]  io_r_172_b,
  input  [1:0]  io_r_173_b,
  input  [1:0]  io_r_174_b,
  input  [1:0]  io_r_175_b,
  input  [1:0]  io_r_176_b,
  input  [1:0]  io_r_177_b,
  input  [1:0]  io_r_178_b,
  input  [1:0]  io_r_179_b,
  input  [1:0]  io_r_180_b,
  input  [1:0]  io_r_181_b,
  input  [1:0]  io_r_182_b,
  input  [1:0]  io_r_183_b,
  input  [1:0]  io_r_184_b,
  input  [1:0]  io_r_185_b,
  input  [1:0]  io_r_186_b,
  input  [1:0]  io_r_187_b,
  input  [1:0]  io_r_188_b,
  input  [1:0]  io_r_189_b,
  input  [1:0]  io_r_190_b,
  input  [1:0]  io_r_191_b,
  input  [1:0]  io_r_192_b,
  input  [1:0]  io_r_193_b,
  input  [1:0]  io_r_194_b,
  input  [1:0]  io_r_195_b,
  input  [1:0]  io_r_196_b,
  input  [1:0]  io_r_197_b,
  input  [1:0]  io_r_198_b,
  input  [1:0]  io_r_199_b,
  input  [1:0]  io_r_200_b,
  input  [1:0]  io_r_201_b,
  input  [1:0]  io_r_202_b,
  input  [1:0]  io_r_203_b,
  input  [1:0]  io_r_204_b,
  input  [1:0]  io_r_205_b,
  input  [1:0]  io_r_206_b,
  input  [1:0]  io_r_207_b,
  input  [1:0]  io_r_208_b,
  input  [1:0]  io_r_209_b,
  input  [1:0]  io_r_210_b,
  input  [1:0]  io_r_211_b,
  input  [1:0]  io_r_212_b,
  input  [1:0]  io_r_213_b,
  input  [1:0]  io_r_214_b,
  input  [1:0]  io_r_215_b,
  input  [1:0]  io_r_216_b,
  input  [1:0]  io_r_217_b,
  input  [1:0]  io_r_218_b,
  input  [1:0]  io_r_219_b,
  input  [1:0]  io_r_220_b,
  input  [1:0]  io_r_221_b,
  input  [1:0]  io_r_222_b,
  input  [1:0]  io_r_223_b,
  input  [1:0]  io_r_224_b,
  input  [1:0]  io_r_225_b,
  input  [1:0]  io_r_226_b,
  input  [1:0]  io_r_227_b,
  input  [1:0]  io_r_228_b,
  input  [1:0]  io_r_229_b,
  input  [1:0]  io_r_230_b,
  input  [1:0]  io_r_231_b,
  input  [1:0]  io_r_232_b,
  input  [1:0]  io_r_233_b,
  input  [1:0]  io_r_234_b,
  input  [1:0]  io_r_235_b,
  input  [1:0]  io_r_236_b,
  input  [1:0]  io_r_237_b,
  input  [1:0]  io_r_238_b,
  input  [1:0]  io_r_239_b,
  input  [1:0]  io_r_240_b,
  input  [1:0]  io_r_241_b,
  input  [1:0]  io_r_242_b,
  input  [1:0]  io_r_243_b,
  input  [1:0]  io_r_244_b,
  input  [1:0]  io_r_245_b,
  input  [1:0]  io_r_246_b,
  input  [1:0]  io_r_247_b,
  input  [1:0]  io_r_248_b,
  input  [1:0]  io_r_249_b,
  input  [1:0]  io_r_250_b,
  input  [1:0]  io_r_251_b,
  input  [1:0]  io_r_252_b,
  input  [1:0]  io_r_253_b,
  input  [1:0]  io_r_254_b,
  input  [1:0]  io_r_255_b,
  input  [1:0]  io_r_256_b,
  input  [1:0]  io_r_257_b,
  input  [1:0]  io_r_258_b,
  input  [1:0]  io_r_259_b,
  input  [1:0]  io_r_260_b,
  input  [1:0]  io_r_261_b,
  input  [1:0]  io_r_262_b,
  input  [1:0]  io_r_263_b,
  input  [1:0]  io_r_264_b,
  input  [1:0]  io_r_265_b,
  input  [1:0]  io_r_266_b,
  input  [1:0]  io_r_267_b,
  input  [1:0]  io_r_268_b,
  input  [1:0]  io_r_269_b,
  input  [1:0]  io_r_270_b,
  input  [1:0]  io_r_271_b,
  input  [1:0]  io_r_272_b,
  input  [1:0]  io_r_273_b,
  input  [1:0]  io_r_274_b,
  input  [1:0]  io_r_275_b,
  input  [1:0]  io_r_276_b,
  input  [1:0]  io_r_277_b,
  input  [1:0]  io_r_278_b,
  input  [1:0]  io_r_279_b,
  input  [1:0]  io_r_280_b,
  input  [1:0]  io_r_281_b,
  input  [1:0]  io_r_282_b,
  input  [1:0]  io_r_283_b,
  input  [1:0]  io_r_284_b,
  input  [1:0]  io_r_285_b,
  input  [1:0]  io_r_286_b,
  input  [1:0]  io_r_287_b,
  input  [1:0]  io_r_288_b,
  input  [1:0]  io_r_289_b,
  input  [1:0]  io_r_290_b,
  input  [1:0]  io_r_291_b,
  input  [1:0]  io_r_292_b,
  input  [1:0]  io_r_293_b,
  input  [1:0]  io_r_294_b,
  input  [1:0]  io_r_295_b,
  input  [1:0]  io_r_296_b,
  input  [1:0]  io_r_297_b,
  input  [1:0]  io_r_298_b,
  input  [1:0]  io_r_299_b,
  input  [1:0]  io_r_300_b,
  input  [1:0]  io_r_301_b,
  input  [1:0]  io_r_302_b,
  input  [1:0]  io_r_303_b,
  input  [1:0]  io_r_304_b,
  input  [1:0]  io_r_305_b,
  input  [1:0]  io_r_306_b,
  input  [1:0]  io_r_307_b,
  input  [1:0]  io_r_308_b,
  input  [1:0]  io_r_309_b,
  input  [1:0]  io_r_310_b,
  input  [1:0]  io_r_311_b,
  input  [1:0]  io_r_312_b,
  input  [1:0]  io_r_313_b,
  input  [1:0]  io_r_314_b,
  input  [1:0]  io_r_315_b,
  input  [1:0]  io_r_316_b,
  input  [1:0]  io_r_317_b,
  input  [1:0]  io_r_318_b,
  input  [1:0]  io_r_319_b,
  input  [1:0]  io_r_320_b,
  input  [1:0]  io_r_321_b,
  input  [1:0]  io_r_322_b,
  input  [1:0]  io_r_323_b,
  input  [1:0]  io_r_324_b,
  input  [1:0]  io_r_325_b,
  input  [1:0]  io_r_326_b,
  input  [1:0]  io_r_327_b,
  input  [1:0]  io_r_328_b,
  input  [1:0]  io_r_329_b,
  input  [1:0]  io_r_330_b,
  input  [1:0]  io_r_331_b,
  input  [1:0]  io_r_332_b,
  input  [1:0]  io_r_333_b,
  input  [1:0]  io_r_334_b,
  input  [1:0]  io_r_335_b,
  input  [1:0]  io_r_336_b,
  input  [1:0]  io_r_337_b,
  input  [1:0]  io_r_338_b,
  input  [1:0]  io_r_339_b,
  input  [1:0]  io_r_340_b,
  input  [1:0]  io_r_341_b,
  input  [1:0]  io_r_342_b,
  input  [1:0]  io_r_343_b,
  input  [1:0]  io_r_344_b,
  input  [1:0]  io_r_345_b,
  input  [1:0]  io_r_346_b,
  input  [1:0]  io_r_347_b,
  input  [1:0]  io_r_348_b,
  input  [1:0]  io_r_349_b,
  input  [1:0]  io_r_350_b,
  input  [1:0]  io_r_351_b,
  input  [1:0]  io_r_352_b,
  input  [1:0]  io_r_353_b,
  input  [1:0]  io_r_354_b,
  input  [1:0]  io_r_355_b,
  input  [1:0]  io_r_356_b,
  input  [1:0]  io_r_357_b,
  input  [1:0]  io_r_358_b,
  input  [1:0]  io_r_359_b,
  input  [1:0]  io_r_360_b,
  input  [1:0]  io_r_361_b,
  input  [1:0]  io_r_362_b,
  input  [1:0]  io_r_363_b,
  input  [1:0]  io_r_364_b,
  input  [1:0]  io_r_365_b,
  input  [1:0]  io_r_366_b,
  input  [1:0]  io_r_367_b,
  input  [1:0]  io_r_368_b,
  input  [1:0]  io_r_369_b,
  input  [1:0]  io_r_370_b,
  input  [1:0]  io_r_371_b,
  input  [1:0]  io_r_372_b,
  input  [1:0]  io_r_373_b,
  input  [1:0]  io_r_374_b,
  input  [1:0]  io_r_375_b,
  input  [1:0]  io_r_376_b,
  input  [1:0]  io_r_377_b,
  input  [1:0]  io_r_378_b,
  input  [1:0]  io_r_379_b,
  input  [1:0]  io_r_380_b,
  input  [1:0]  io_r_381_b,
  input  [1:0]  io_r_382_b,
  input  [1:0]  io_r_383_b,
  input  [1:0]  io_r_384_b,
  input  [1:0]  io_r_385_b,
  input  [1:0]  io_r_386_b,
  input  [1:0]  io_r_387_b,
  input  [1:0]  io_r_388_b,
  input  [1:0]  io_r_389_b,
  input  [1:0]  io_r_390_b,
  input  [1:0]  io_r_391_b,
  input  [1:0]  io_r_392_b,
  input  [1:0]  io_r_393_b,
  input  [1:0]  io_r_394_b,
  input  [1:0]  io_r_395_b,
  input  [1:0]  io_r_396_b,
  input  [1:0]  io_r_397_b,
  input  [1:0]  io_r_398_b,
  input  [1:0]  io_r_399_b,
  input  [1:0]  io_r_400_b,
  input  [1:0]  io_r_401_b,
  input  [1:0]  io_r_402_b,
  input  [1:0]  io_r_403_b,
  input  [1:0]  io_r_404_b,
  input  [1:0]  io_r_405_b,
  input  [1:0]  io_r_406_b,
  input  [1:0]  io_r_407_b,
  input  [1:0]  io_r_408_b,
  input  [1:0]  io_r_409_b,
  input  [1:0]  io_r_410_b,
  input  [1:0]  io_r_411_b,
  input  [1:0]  io_r_412_b,
  input  [1:0]  io_r_413_b,
  input  [1:0]  io_r_414_b,
  input  [1:0]  io_r_415_b,
  input  [1:0]  io_r_416_b,
  input  [1:0]  io_r_417_b,
  input  [1:0]  io_r_418_b,
  input  [1:0]  io_r_419_b,
  input  [1:0]  io_r_420_b,
  input  [1:0]  io_r_421_b,
  input  [1:0]  io_r_422_b,
  input  [1:0]  io_r_423_b,
  input  [1:0]  io_r_424_b,
  input  [1:0]  io_r_425_b,
  input  [1:0]  io_r_426_b,
  input  [1:0]  io_r_427_b,
  input  [1:0]  io_r_428_b,
  input  [1:0]  io_r_429_b,
  input  [1:0]  io_r_430_b,
  input  [1:0]  io_r_431_b,
  input  [1:0]  io_r_432_b,
  input  [1:0]  io_r_433_b,
  input  [1:0]  io_r_434_b,
  input  [1:0]  io_r_435_b,
  input  [1:0]  io_r_436_b,
  input  [1:0]  io_r_437_b,
  input  [1:0]  io_r_438_b,
  input  [1:0]  io_r_439_b,
  input  [1:0]  io_r_440_b,
  input  [1:0]  io_r_441_b,
  input  [1:0]  io_r_442_b,
  input  [1:0]  io_r_443_b,
  input  [1:0]  io_r_444_b,
  input  [1:0]  io_r_445_b,
  input  [1:0]  io_r_446_b,
  input  [1:0]  io_r_447_b,
  input  [1:0]  io_r_448_b,
  input  [1:0]  io_r_449_b,
  input  [1:0]  io_r_450_b,
  input  [1:0]  io_r_451_b,
  input  [1:0]  io_r_452_b,
  input  [1:0]  io_r_453_b,
  input  [1:0]  io_r_454_b,
  input  [1:0]  io_r_455_b,
  input  [1:0]  io_r_456_b,
  input  [1:0]  io_r_457_b,
  input  [1:0]  io_r_458_b,
  input  [1:0]  io_r_459_b,
  input  [1:0]  io_r_460_b,
  input  [1:0]  io_r_461_b,
  input  [1:0]  io_r_462_b,
  input  [1:0]  io_r_463_b,
  input  [1:0]  io_r_464_b,
  input  [1:0]  io_r_465_b,
  input  [1:0]  io_r_466_b,
  input  [1:0]  io_r_467_b,
  input  [1:0]  io_r_468_b,
  input  [1:0]  io_r_469_b,
  input  [1:0]  io_r_470_b,
  input  [1:0]  io_r_471_b,
  input  [1:0]  io_r_472_b,
  input  [1:0]  io_r_473_b,
  input  [1:0]  io_r_474_b,
  input  [1:0]  io_r_475_b,
  input  [1:0]  io_r_476_b,
  input  [1:0]  io_r_477_b,
  input  [1:0]  io_r_478_b,
  input  [1:0]  io_r_479_b,
  input  [1:0]  io_r_480_b,
  input  [1:0]  io_r_481_b,
  input  [1:0]  io_r_482_b,
  input  [1:0]  io_r_483_b,
  input  [1:0]  io_r_484_b,
  input  [1:0]  io_r_485_b,
  input  [1:0]  io_r_486_b,
  input  [1:0]  io_r_487_b,
  input  [1:0]  io_r_488_b,
  input  [1:0]  io_r_489_b,
  input  [1:0]  io_r_490_b,
  input  [1:0]  io_r_491_b,
  input  [1:0]  io_r_492_b,
  input  [1:0]  io_r_493_b,
  input  [1:0]  io_r_494_b,
  input  [1:0]  io_r_495_b,
  input  [1:0]  io_r_496_b,
  input  [1:0]  io_r_497_b,
  input  [1:0]  io_r_498_b,
  input  [1:0]  io_r_499_b,
  input  [1:0]  io_r_500_b,
  input  [1:0]  io_r_501_b,
  input  [1:0]  io_r_502_b,
  input  [1:0]  io_r_503_b,
  input  [1:0]  io_r_504_b,
  input  [1:0]  io_r_505_b,
  input  [1:0]  io_r_506_b,
  input  [1:0]  io_r_507_b,
  input  [1:0]  io_r_508_b,
  input  [1:0]  io_r_509_b,
  input  [1:0]  io_r_510_b,
  input  [1:0]  io_r_511_b,
  input  [1:0]  io_r_512_b,
  input  [1:0]  io_r_513_b,
  input  [1:0]  io_r_514_b,
  input  [1:0]  io_r_515_b,
  input  [1:0]  io_r_516_b,
  input  [1:0]  io_r_517_b,
  input  [1:0]  io_r_518_b,
  input  [1:0]  io_r_519_b,
  input  [1:0]  io_r_520_b,
  input  [1:0]  io_r_521_b,
  input  [1:0]  io_r_522_b,
  input  [1:0]  io_r_523_b,
  input  [1:0]  io_r_524_b,
  input  [1:0]  io_r_525_b,
  input  [1:0]  io_r_526_b,
  input  [1:0]  io_r_527_b,
  input  [1:0]  io_r_528_b,
  input  [1:0]  io_r_529_b,
  input  [1:0]  io_r_530_b,
  input  [1:0]  io_r_531_b,
  input  [1:0]  io_r_532_b,
  input  [1:0]  io_r_533_b,
  input  [1:0]  io_r_534_b,
  input  [1:0]  io_r_535_b,
  input  [1:0]  io_r_536_b,
  input  [1:0]  io_r_537_b,
  input  [1:0]  io_r_538_b,
  input  [1:0]  io_r_539_b,
  input  [1:0]  io_r_540_b,
  input  [1:0]  io_r_541_b,
  input  [1:0]  io_r_542_b,
  input  [1:0]  io_r_543_b,
  input  [1:0]  io_r_544_b,
  input  [1:0]  io_r_545_b,
  input  [1:0]  io_r_546_b,
  input  [1:0]  io_r_547_b,
  input  [1:0]  io_r_548_b,
  input  [1:0]  io_r_549_b,
  input  [1:0]  io_r_550_b,
  input  [1:0]  io_r_551_b,
  input  [1:0]  io_r_552_b,
  input  [1:0]  io_r_553_b,
  input  [1:0]  io_r_554_b,
  input  [1:0]  io_r_555_b,
  input  [1:0]  io_r_556_b,
  input  [1:0]  io_r_557_b,
  input  [1:0]  io_r_558_b,
  input  [1:0]  io_r_559_b,
  input  [1:0]  io_r_560_b,
  input  [1:0]  io_r_561_b,
  input  [1:0]  io_r_562_b,
  input  [1:0]  io_r_563_b,
  input  [1:0]  io_r_564_b,
  input  [1:0]  io_r_565_b,
  input  [1:0]  io_r_566_b,
  input  [1:0]  io_r_567_b,
  input  [1:0]  io_r_568_b,
  input  [1:0]  io_r_569_b,
  input  [1:0]  io_r_570_b,
  input  [1:0]  io_r_571_b,
  input  [1:0]  io_r_572_b,
  input  [1:0]  io_r_573_b,
  input  [1:0]  io_r_574_b,
  input  [1:0]  io_r_575_b,
  input  [1:0]  io_r_576_b,
  input  [1:0]  io_r_577_b,
  input  [1:0]  io_r_578_b,
  input  [1:0]  io_r_579_b,
  input  [1:0]  io_r_580_b,
  input  [1:0]  io_r_581_b,
  input  [1:0]  io_r_582_b,
  input  [1:0]  io_r_583_b,
  input  [1:0]  io_r_584_b,
  input  [1:0]  io_r_585_b,
  input  [1:0]  io_r_586_b,
  input  [1:0]  io_r_587_b,
  input  [1:0]  io_r_588_b,
  input  [1:0]  io_r_589_b,
  input  [1:0]  io_r_590_b,
  input  [1:0]  io_r_591_b,
  input  [1:0]  io_r_592_b,
  input  [1:0]  io_r_593_b,
  input  [1:0]  io_r_594_b,
  input  [1:0]  io_r_595_b,
  input  [1:0]  io_r_596_b,
  input  [1:0]  io_r_597_b,
  input  [1:0]  io_r_598_b,
  input  [1:0]  io_r_599_b,
  input  [1:0]  io_r_600_b,
  input  [1:0]  io_r_601_b,
  input  [1:0]  io_r_602_b,
  input  [1:0]  io_r_603_b,
  input  [1:0]  io_r_604_b,
  input  [1:0]  io_r_605_b,
  input  [1:0]  io_r_606_b,
  input  [1:0]  io_r_607_b,
  input  [1:0]  io_r_608_b,
  input  [1:0]  io_r_609_b,
  input  [1:0]  io_r_610_b,
  input  [1:0]  io_r_611_b,
  input  [1:0]  io_r_612_b,
  input  [1:0]  io_r_613_b,
  input  [1:0]  io_r_614_b,
  input  [1:0]  io_r_615_b,
  input  [1:0]  io_r_616_b,
  input  [1:0]  io_r_617_b,
  input  [1:0]  io_r_618_b,
  input  [1:0]  io_r_619_b,
  input  [1:0]  io_r_620_b,
  input  [1:0]  io_r_621_b,
  input  [1:0]  io_r_622_b,
  input  [1:0]  io_r_623_b,
  input  [1:0]  io_r_624_b,
  input  [1:0]  io_r_625_b,
  input  [1:0]  io_r_626_b,
  input  [1:0]  io_r_627_b,
  input  [1:0]  io_r_628_b,
  input  [1:0]  io_r_629_b,
  input  [1:0]  io_r_630_b,
  input  [1:0]  io_r_631_b,
  input  [1:0]  io_r_632_b,
  input  [1:0]  io_r_633_b,
  input  [1:0]  io_r_634_b,
  input  [1:0]  io_r_635_b,
  input  [1:0]  io_r_636_b,
  input  [1:0]  io_r_637_b,
  input  [1:0]  io_r_638_b,
  input  [1:0]  io_r_639_b,
  input  [1:0]  io_r_640_b,
  input  [1:0]  io_r_641_b,
  input  [1:0]  io_r_642_b,
  input  [1:0]  io_r_643_b,
  input  [1:0]  io_r_644_b,
  input  [1:0]  io_r_645_b,
  input  [1:0]  io_r_646_b,
  input  [1:0]  io_r_647_b,
  input  [1:0]  io_r_648_b,
  input  [1:0]  io_r_649_b,
  input  [1:0]  io_r_650_b,
  input  [1:0]  io_r_651_b,
  input  [1:0]  io_r_652_b,
  input  [1:0]  io_r_653_b,
  input  [1:0]  io_r_654_b,
  input  [1:0]  io_r_655_b,
  input  [1:0]  io_r_656_b,
  input  [1:0]  io_r_657_b,
  input  [1:0]  io_r_658_b,
  input  [1:0]  io_r_659_b,
  input  [1:0]  io_r_660_b,
  input  [1:0]  io_r_661_b,
  input  [1:0]  io_r_662_b,
  input  [1:0]  io_r_663_b,
  input  [1:0]  io_r_664_b,
  input  [1:0]  io_r_665_b,
  input  [1:0]  io_r_666_b,
  input  [1:0]  io_r_667_b,
  input  [1:0]  io_r_668_b,
  input  [1:0]  io_r_669_b,
  input  [1:0]  io_r_670_b,
  input  [1:0]  io_r_671_b,
  input  [1:0]  io_r_672_b,
  input  [1:0]  io_r_673_b,
  input  [1:0]  io_r_674_b,
  input  [1:0]  io_r_675_b,
  input  [1:0]  io_r_676_b,
  input  [1:0]  io_r_677_b,
  input  [1:0]  io_r_678_b,
  input  [1:0]  io_r_679_b,
  input  [1:0]  io_r_680_b,
  input  [1:0]  io_r_681_b,
  input  [1:0]  io_r_682_b,
  input  [1:0]  io_r_683_b,
  input  [1:0]  io_r_684_b,
  input  [1:0]  io_r_685_b,
  input  [1:0]  io_r_686_b,
  input  [1:0]  io_r_687_b,
  input  [1:0]  io_r_688_b,
  input  [1:0]  io_r_689_b,
  input  [1:0]  io_r_690_b,
  input  [1:0]  io_r_691_b,
  input  [1:0]  io_r_692_b,
  input  [1:0]  io_r_693_b,
  input  [1:0]  io_r_694_b,
  input  [1:0]  io_r_695_b,
  input  [1:0]  io_r_696_b,
  input  [1:0]  io_r_697_b,
  input  [1:0]  io_r_698_b,
  input  [1:0]  io_r_699_b,
  input  [1:0]  io_r_700_b,
  input  [1:0]  io_r_701_b,
  input  [1:0]  io_r_702_b,
  input  [1:0]  io_r_703_b,
  input  [1:0]  io_r_704_b,
  input  [1:0]  io_r_705_b,
  input  [1:0]  io_r_706_b,
  input  [1:0]  io_r_707_b,
  input  [1:0]  io_r_708_b,
  input  [1:0]  io_r_709_b,
  input  [1:0]  io_r_710_b,
  input  [1:0]  io_r_711_b,
  input  [1:0]  io_r_712_b,
  input  [1:0]  io_r_713_b,
  input  [1:0]  io_r_714_b,
  input  [1:0]  io_r_715_b,
  input  [1:0]  io_r_716_b,
  input  [1:0]  io_r_717_b,
  input  [1:0]  io_r_718_b,
  input  [1:0]  io_r_719_b,
  input  [1:0]  io_r_720_b,
  input  [1:0]  io_r_721_b,
  input  [1:0]  io_r_722_b,
  input  [1:0]  io_r_723_b,
  input  [1:0]  io_r_724_b,
  input  [1:0]  io_r_725_b,
  input  [1:0]  io_r_726_b,
  input  [1:0]  io_r_727_b,
  input  [1:0]  io_r_728_b,
  input  [1:0]  io_r_729_b,
  input  [1:0]  io_r_730_b,
  input  [1:0]  io_r_731_b,
  input  [1:0]  io_r_732_b,
  input  [1:0]  io_r_733_b,
  input  [1:0]  io_r_734_b,
  input  [1:0]  io_r_735_b,
  input  [1:0]  io_r_736_b,
  input  [1:0]  io_r_737_b,
  input  [1:0]  io_r_738_b,
  input  [1:0]  io_r_739_b,
  input  [1:0]  io_r_740_b,
  input  [1:0]  io_r_741_b,
  input  [1:0]  io_r_742_b,
  input  [1:0]  io_r_743_b,
  input  [1:0]  io_r_744_b,
  input  [1:0]  io_r_745_b,
  input  [1:0]  io_r_746_b,
  input  [1:0]  io_r_747_b,
  input  [1:0]  io_r_748_b,
  input  [1:0]  io_r_749_b,
  input         io_start,
  output [15:0] io_result,
  output        io_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
`endif // RANDOMIZE_REG_INIT
  wire [1:0] array_0_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_0_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_1_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_1_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_2_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_2_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_3_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_3_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_4_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_4_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_5_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_5_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_6_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_6_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_7_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_7_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_8_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_8_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_9_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_9_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_10_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_10_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_11_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_11_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_12_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_12_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_13_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_13_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_14_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_14_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_15_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_15_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_16_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_16_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_17_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_17_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_18_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_18_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_19_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_19_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_20_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_20_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_21_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_21_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_22_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_22_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_23_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_23_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_24_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_24_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_25_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_25_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_26_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_26_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_27_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_27_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_28_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_28_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_29_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_29_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_v_o; // @[SWChisel.scala 170:39]
  wire  r_count_0_clock; // @[SWChisel.scala 171:41]
  wire  r_count_0_reset; // @[SWChisel.scala 171:41]
  wire  r_count_0_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_0_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_1_clock; // @[SWChisel.scala 171:41]
  wire  r_count_1_reset; // @[SWChisel.scala 171:41]
  wire  r_count_1_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_1_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_2_clock; // @[SWChisel.scala 171:41]
  wire  r_count_2_reset; // @[SWChisel.scala 171:41]
  wire  r_count_2_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_2_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_3_clock; // @[SWChisel.scala 171:41]
  wire  r_count_3_reset; // @[SWChisel.scala 171:41]
  wire  r_count_3_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_3_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_4_clock; // @[SWChisel.scala 171:41]
  wire  r_count_4_reset; // @[SWChisel.scala 171:41]
  wire  r_count_4_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_4_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_5_clock; // @[SWChisel.scala 171:41]
  wire  r_count_5_reset; // @[SWChisel.scala 171:41]
  wire  r_count_5_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_5_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_6_clock; // @[SWChisel.scala 171:41]
  wire  r_count_6_reset; // @[SWChisel.scala 171:41]
  wire  r_count_6_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_6_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_7_clock; // @[SWChisel.scala 171:41]
  wire  r_count_7_reset; // @[SWChisel.scala 171:41]
  wire  r_count_7_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_7_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_8_clock; // @[SWChisel.scala 171:41]
  wire  r_count_8_reset; // @[SWChisel.scala 171:41]
  wire  r_count_8_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_8_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_9_clock; // @[SWChisel.scala 171:41]
  wire  r_count_9_reset; // @[SWChisel.scala 171:41]
  wire  r_count_9_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_9_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_10_clock; // @[SWChisel.scala 171:41]
  wire  r_count_10_reset; // @[SWChisel.scala 171:41]
  wire  r_count_10_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_10_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_11_clock; // @[SWChisel.scala 171:41]
  wire  r_count_11_reset; // @[SWChisel.scala 171:41]
  wire  r_count_11_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_11_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_12_clock; // @[SWChisel.scala 171:41]
  wire  r_count_12_reset; // @[SWChisel.scala 171:41]
  wire  r_count_12_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_12_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_13_clock; // @[SWChisel.scala 171:41]
  wire  r_count_13_reset; // @[SWChisel.scala 171:41]
  wire  r_count_13_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_13_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_14_clock; // @[SWChisel.scala 171:41]
  wire  r_count_14_reset; // @[SWChisel.scala 171:41]
  wire  r_count_14_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_14_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_15_clock; // @[SWChisel.scala 171:41]
  wire  r_count_15_reset; // @[SWChisel.scala 171:41]
  wire  r_count_15_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_15_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_16_clock; // @[SWChisel.scala 171:41]
  wire  r_count_16_reset; // @[SWChisel.scala 171:41]
  wire  r_count_16_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_16_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_17_clock; // @[SWChisel.scala 171:41]
  wire  r_count_17_reset; // @[SWChisel.scala 171:41]
  wire  r_count_17_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_17_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_18_clock; // @[SWChisel.scala 171:41]
  wire  r_count_18_reset; // @[SWChisel.scala 171:41]
  wire  r_count_18_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_18_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_19_clock; // @[SWChisel.scala 171:41]
  wire  r_count_19_reset; // @[SWChisel.scala 171:41]
  wire  r_count_19_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_19_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_20_clock; // @[SWChisel.scala 171:41]
  wire  r_count_20_reset; // @[SWChisel.scala 171:41]
  wire  r_count_20_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_20_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_21_clock; // @[SWChisel.scala 171:41]
  wire  r_count_21_reset; // @[SWChisel.scala 171:41]
  wire  r_count_21_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_21_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_22_clock; // @[SWChisel.scala 171:41]
  wire  r_count_22_reset; // @[SWChisel.scala 171:41]
  wire  r_count_22_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_22_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_23_clock; // @[SWChisel.scala 171:41]
  wire  r_count_23_reset; // @[SWChisel.scala 171:41]
  wire  r_count_23_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_23_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_24_clock; // @[SWChisel.scala 171:41]
  wire  r_count_24_reset; // @[SWChisel.scala 171:41]
  wire  r_count_24_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_24_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_25_clock; // @[SWChisel.scala 171:41]
  wire  r_count_25_reset; // @[SWChisel.scala 171:41]
  wire  r_count_25_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_25_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_26_clock; // @[SWChisel.scala 171:41]
  wire  r_count_26_reset; // @[SWChisel.scala 171:41]
  wire  r_count_26_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_26_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_27_clock; // @[SWChisel.scala 171:41]
  wire  r_count_27_reset; // @[SWChisel.scala 171:41]
  wire  r_count_27_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_27_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_28_clock; // @[SWChisel.scala 171:41]
  wire  r_count_28_reset; // @[SWChisel.scala 171:41]
  wire  r_count_28_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_28_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_29_clock; // @[SWChisel.scala 171:41]
  wire  r_count_29_reset; // @[SWChisel.scala 171:41]
  wire  r_count_29_io_en; // @[SWChisel.scala 171:41]
  wire [9:0] r_count_29_io_out; // @[SWChisel.scala 171:41]
  wire  max_clock; // @[SWChisel.scala 174:19]
  wire  max_reset; // @[SWChisel.scala 174:19]
  wire  max_io_start; // @[SWChisel.scala 174:19]
  wire [15:0] max_io_in; // @[SWChisel.scala 174:19]
  wire  max_io_done; // @[SWChisel.scala 174:19]
  wire [15:0] max_io_out; // @[SWChisel.scala 174:19]
  reg [15:0] E_0; // @[SWChisel.scala 162:18]
  reg [15:0] E_1; // @[SWChisel.scala 162:18]
  reg [15:0] E_2; // @[SWChisel.scala 162:18]
  reg [15:0] E_3; // @[SWChisel.scala 162:18]
  reg [15:0] E_4; // @[SWChisel.scala 162:18]
  reg [15:0] E_5; // @[SWChisel.scala 162:18]
  reg [15:0] E_6; // @[SWChisel.scala 162:18]
  reg [15:0] E_7; // @[SWChisel.scala 162:18]
  reg [15:0] E_8; // @[SWChisel.scala 162:18]
  reg [15:0] E_9; // @[SWChisel.scala 162:18]
  reg [15:0] E_10; // @[SWChisel.scala 162:18]
  reg [15:0] E_11; // @[SWChisel.scala 162:18]
  reg [15:0] E_12; // @[SWChisel.scala 162:18]
  reg [15:0] E_13; // @[SWChisel.scala 162:18]
  reg [15:0] E_14; // @[SWChisel.scala 162:18]
  reg [15:0] E_15; // @[SWChisel.scala 162:18]
  reg [15:0] E_16; // @[SWChisel.scala 162:18]
  reg [15:0] E_17; // @[SWChisel.scala 162:18]
  reg [15:0] E_18; // @[SWChisel.scala 162:18]
  reg [15:0] E_19; // @[SWChisel.scala 162:18]
  reg [15:0] E_20; // @[SWChisel.scala 162:18]
  reg [15:0] E_21; // @[SWChisel.scala 162:18]
  reg [15:0] E_22; // @[SWChisel.scala 162:18]
  reg [15:0] E_23; // @[SWChisel.scala 162:18]
  reg [15:0] E_24; // @[SWChisel.scala 162:18]
  reg [15:0] E_25; // @[SWChisel.scala 162:18]
  reg [15:0] E_26; // @[SWChisel.scala 162:18]
  reg [15:0] E_27; // @[SWChisel.scala 162:18]
  reg [15:0] E_28; // @[SWChisel.scala 162:18]
  reg [15:0] E_29; // @[SWChisel.scala 162:18]
  reg [15:0] F_1; // @[SWChisel.scala 163:18]
  reg [15:0] F_2; // @[SWChisel.scala 163:18]
  reg [15:0] F_3; // @[SWChisel.scala 163:18]
  reg [15:0] F_4; // @[SWChisel.scala 163:18]
  reg [15:0] F_5; // @[SWChisel.scala 163:18]
  reg [15:0] F_6; // @[SWChisel.scala 163:18]
  reg [15:0] F_7; // @[SWChisel.scala 163:18]
  reg [15:0] F_8; // @[SWChisel.scala 163:18]
  reg [15:0] F_9; // @[SWChisel.scala 163:18]
  reg [15:0] F_10; // @[SWChisel.scala 163:18]
  reg [15:0] F_11; // @[SWChisel.scala 163:18]
  reg [15:0] F_12; // @[SWChisel.scala 163:18]
  reg [15:0] F_13; // @[SWChisel.scala 163:18]
  reg [15:0] F_14; // @[SWChisel.scala 163:18]
  reg [15:0] F_15; // @[SWChisel.scala 163:18]
  reg [15:0] F_16; // @[SWChisel.scala 163:18]
  reg [15:0] F_17; // @[SWChisel.scala 163:18]
  reg [15:0] F_18; // @[SWChisel.scala 163:18]
  reg [15:0] F_19; // @[SWChisel.scala 163:18]
  reg [15:0] F_20; // @[SWChisel.scala 163:18]
  reg [15:0] F_21; // @[SWChisel.scala 163:18]
  reg [15:0] F_22; // @[SWChisel.scala 163:18]
  reg [15:0] F_23; // @[SWChisel.scala 163:18]
  reg [15:0] F_24; // @[SWChisel.scala 163:18]
  reg [15:0] F_25; // @[SWChisel.scala 163:18]
  reg [15:0] F_26; // @[SWChisel.scala 163:18]
  reg [15:0] F_27; // @[SWChisel.scala 163:18]
  reg [15:0] F_28; // @[SWChisel.scala 163:18]
  reg [15:0] F_29; // @[SWChisel.scala 163:18]
  reg [15:0] V1_0; // @[SWChisel.scala 164:19]
  reg [15:0] V1_1; // @[SWChisel.scala 164:19]
  reg [15:0] V1_2; // @[SWChisel.scala 164:19]
  reg [15:0] V1_3; // @[SWChisel.scala 164:19]
  reg [15:0] V1_4; // @[SWChisel.scala 164:19]
  reg [15:0] V1_5; // @[SWChisel.scala 164:19]
  reg [15:0] V1_6; // @[SWChisel.scala 164:19]
  reg [15:0] V1_7; // @[SWChisel.scala 164:19]
  reg [15:0] V1_8; // @[SWChisel.scala 164:19]
  reg [15:0] V1_9; // @[SWChisel.scala 164:19]
  reg [15:0] V1_10; // @[SWChisel.scala 164:19]
  reg [15:0] V1_11; // @[SWChisel.scala 164:19]
  reg [15:0] V1_12; // @[SWChisel.scala 164:19]
  reg [15:0] V1_13; // @[SWChisel.scala 164:19]
  reg [15:0] V1_14; // @[SWChisel.scala 164:19]
  reg [15:0] V1_15; // @[SWChisel.scala 164:19]
  reg [15:0] V1_16; // @[SWChisel.scala 164:19]
  reg [15:0] V1_17; // @[SWChisel.scala 164:19]
  reg [15:0] V1_18; // @[SWChisel.scala 164:19]
  reg [15:0] V1_19; // @[SWChisel.scala 164:19]
  reg [15:0] V1_20; // @[SWChisel.scala 164:19]
  reg [15:0] V1_21; // @[SWChisel.scala 164:19]
  reg [15:0] V1_22; // @[SWChisel.scala 164:19]
  reg [15:0] V1_23; // @[SWChisel.scala 164:19]
  reg [15:0] V1_24; // @[SWChisel.scala 164:19]
  reg [15:0] V1_25; // @[SWChisel.scala 164:19]
  reg [15:0] V1_26; // @[SWChisel.scala 164:19]
  reg [15:0] V1_27; // @[SWChisel.scala 164:19]
  reg [15:0] V1_28; // @[SWChisel.scala 164:19]
  reg [15:0] V1_29; // @[SWChisel.scala 164:19]
  reg [15:0] V1_30; // @[SWChisel.scala 164:19]
  reg [15:0] V2_0; // @[SWChisel.scala 166:19]
  reg [15:0] V2_1; // @[SWChisel.scala 166:19]
  reg [15:0] V2_2; // @[SWChisel.scala 166:19]
  reg [15:0] V2_3; // @[SWChisel.scala 166:19]
  reg [15:0] V2_4; // @[SWChisel.scala 166:19]
  reg [15:0] V2_5; // @[SWChisel.scala 166:19]
  reg [15:0] V2_6; // @[SWChisel.scala 166:19]
  reg [15:0] V2_7; // @[SWChisel.scala 166:19]
  reg [15:0] V2_8; // @[SWChisel.scala 166:19]
  reg [15:0] V2_9; // @[SWChisel.scala 166:19]
  reg [15:0] V2_10; // @[SWChisel.scala 166:19]
  reg [15:0] V2_11; // @[SWChisel.scala 166:19]
  reg [15:0] V2_12; // @[SWChisel.scala 166:19]
  reg [15:0] V2_13; // @[SWChisel.scala 166:19]
  reg [15:0] V2_14; // @[SWChisel.scala 166:19]
  reg [15:0] V2_15; // @[SWChisel.scala 166:19]
  reg [15:0] V2_16; // @[SWChisel.scala 166:19]
  reg [15:0] V2_17; // @[SWChisel.scala 166:19]
  reg [15:0] V2_18; // @[SWChisel.scala 166:19]
  reg [15:0] V2_19; // @[SWChisel.scala 166:19]
  reg [15:0] V2_20; // @[SWChisel.scala 166:19]
  reg [15:0] V2_21; // @[SWChisel.scala 166:19]
  reg [15:0] V2_22; // @[SWChisel.scala 166:19]
  reg [15:0] V2_23; // @[SWChisel.scala 166:19]
  reg [15:0] V2_24; // @[SWChisel.scala 166:19]
  reg [15:0] V2_25; // @[SWChisel.scala 166:19]
  reg [15:0] V2_26; // @[SWChisel.scala 166:19]
  reg [15:0] V2_27; // @[SWChisel.scala 166:19]
  reg [15:0] V2_28; // @[SWChisel.scala 166:19]
  reg [15:0] V2_29; // @[SWChisel.scala 166:19]
  reg  start_reg_0; // @[SWChisel.scala 167:26]
  reg  start_reg_1; // @[SWChisel.scala 167:26]
  reg  start_reg_2; // @[SWChisel.scala 167:26]
  reg  start_reg_3; // @[SWChisel.scala 167:26]
  reg  start_reg_4; // @[SWChisel.scala 167:26]
  reg  start_reg_5; // @[SWChisel.scala 167:26]
  reg  start_reg_6; // @[SWChisel.scala 167:26]
  reg  start_reg_7; // @[SWChisel.scala 167:26]
  reg  start_reg_8; // @[SWChisel.scala 167:26]
  reg  start_reg_9; // @[SWChisel.scala 167:26]
  reg  start_reg_10; // @[SWChisel.scala 167:26]
  reg  start_reg_11; // @[SWChisel.scala 167:26]
  reg  start_reg_12; // @[SWChisel.scala 167:26]
  reg  start_reg_13; // @[SWChisel.scala 167:26]
  reg  start_reg_14; // @[SWChisel.scala 167:26]
  reg  start_reg_15; // @[SWChisel.scala 167:26]
  reg  start_reg_16; // @[SWChisel.scala 167:26]
  reg  start_reg_17; // @[SWChisel.scala 167:26]
  reg  start_reg_18; // @[SWChisel.scala 167:26]
  reg  start_reg_19; // @[SWChisel.scala 167:26]
  reg  start_reg_20; // @[SWChisel.scala 167:26]
  reg  start_reg_21; // @[SWChisel.scala 167:26]
  reg  start_reg_22; // @[SWChisel.scala 167:26]
  reg  start_reg_23; // @[SWChisel.scala 167:26]
  reg  start_reg_24; // @[SWChisel.scala 167:26]
  reg  start_reg_25; // @[SWChisel.scala 167:26]
  reg  start_reg_26; // @[SWChisel.scala 167:26]
  reg  start_reg_27; // @[SWChisel.scala 167:26]
  reg  start_reg_28; // @[SWChisel.scala 167:26]
  reg  start_reg_29; // @[SWChisel.scala 167:26]
  wire [1:0] _GEN_91 = 10'h1 == r_count_0_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_92 = 10'h2 == r_count_0_io_out ? io_r_2_b : _GEN_91; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_93 = 10'h3 == r_count_0_io_out ? io_r_3_b : _GEN_92; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_94 = 10'h4 == r_count_0_io_out ? io_r_4_b : _GEN_93; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_95 = 10'h5 == r_count_0_io_out ? io_r_5_b : _GEN_94; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_96 = 10'h6 == r_count_0_io_out ? io_r_6_b : _GEN_95; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_97 = 10'h7 == r_count_0_io_out ? io_r_7_b : _GEN_96; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_98 = 10'h8 == r_count_0_io_out ? io_r_8_b : _GEN_97; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_99 = 10'h9 == r_count_0_io_out ? io_r_9_b : _GEN_98; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_100 = 10'ha == r_count_0_io_out ? io_r_10_b : _GEN_99; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_101 = 10'hb == r_count_0_io_out ? io_r_11_b : _GEN_100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_102 = 10'hc == r_count_0_io_out ? io_r_12_b : _GEN_101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_103 = 10'hd == r_count_0_io_out ? io_r_13_b : _GEN_102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_104 = 10'he == r_count_0_io_out ? io_r_14_b : _GEN_103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_105 = 10'hf == r_count_0_io_out ? io_r_15_b : _GEN_104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_106 = 10'h10 == r_count_0_io_out ? io_r_16_b : _GEN_105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_107 = 10'h11 == r_count_0_io_out ? io_r_17_b : _GEN_106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_108 = 10'h12 == r_count_0_io_out ? io_r_18_b : _GEN_107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_109 = 10'h13 == r_count_0_io_out ? io_r_19_b : _GEN_108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_110 = 10'h14 == r_count_0_io_out ? io_r_20_b : _GEN_109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_111 = 10'h15 == r_count_0_io_out ? io_r_21_b : _GEN_110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_112 = 10'h16 == r_count_0_io_out ? io_r_22_b : _GEN_111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_113 = 10'h17 == r_count_0_io_out ? io_r_23_b : _GEN_112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_114 = 10'h18 == r_count_0_io_out ? io_r_24_b : _GEN_113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_115 = 10'h19 == r_count_0_io_out ? io_r_25_b : _GEN_114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_116 = 10'h1a == r_count_0_io_out ? io_r_26_b : _GEN_115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_117 = 10'h1b == r_count_0_io_out ? io_r_27_b : _GEN_116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_118 = 10'h1c == r_count_0_io_out ? io_r_28_b : _GEN_117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_119 = 10'h1d == r_count_0_io_out ? io_r_29_b : _GEN_118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_120 = 10'h1e == r_count_0_io_out ? io_r_30_b : _GEN_119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_121 = 10'h1f == r_count_0_io_out ? io_r_31_b : _GEN_120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_122 = 10'h20 == r_count_0_io_out ? io_r_32_b : _GEN_121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_123 = 10'h21 == r_count_0_io_out ? io_r_33_b : _GEN_122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_124 = 10'h22 == r_count_0_io_out ? io_r_34_b : _GEN_123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_125 = 10'h23 == r_count_0_io_out ? io_r_35_b : _GEN_124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_126 = 10'h24 == r_count_0_io_out ? io_r_36_b : _GEN_125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_127 = 10'h25 == r_count_0_io_out ? io_r_37_b : _GEN_126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_128 = 10'h26 == r_count_0_io_out ? io_r_38_b : _GEN_127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_129 = 10'h27 == r_count_0_io_out ? io_r_39_b : _GEN_128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_130 = 10'h28 == r_count_0_io_out ? io_r_40_b : _GEN_129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_131 = 10'h29 == r_count_0_io_out ? io_r_41_b : _GEN_130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_132 = 10'h2a == r_count_0_io_out ? io_r_42_b : _GEN_131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_133 = 10'h2b == r_count_0_io_out ? io_r_43_b : _GEN_132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_134 = 10'h2c == r_count_0_io_out ? io_r_44_b : _GEN_133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_135 = 10'h2d == r_count_0_io_out ? io_r_45_b : _GEN_134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_136 = 10'h2e == r_count_0_io_out ? io_r_46_b : _GEN_135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_137 = 10'h2f == r_count_0_io_out ? io_r_47_b : _GEN_136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_138 = 10'h30 == r_count_0_io_out ? io_r_48_b : _GEN_137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_139 = 10'h31 == r_count_0_io_out ? io_r_49_b : _GEN_138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_140 = 10'h32 == r_count_0_io_out ? io_r_50_b : _GEN_139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_141 = 10'h33 == r_count_0_io_out ? io_r_51_b : _GEN_140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_142 = 10'h34 == r_count_0_io_out ? io_r_52_b : _GEN_141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_143 = 10'h35 == r_count_0_io_out ? io_r_53_b : _GEN_142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_144 = 10'h36 == r_count_0_io_out ? io_r_54_b : _GEN_143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_145 = 10'h37 == r_count_0_io_out ? io_r_55_b : _GEN_144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_146 = 10'h38 == r_count_0_io_out ? io_r_56_b : _GEN_145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_147 = 10'h39 == r_count_0_io_out ? io_r_57_b : _GEN_146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_148 = 10'h3a == r_count_0_io_out ? io_r_58_b : _GEN_147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_149 = 10'h3b == r_count_0_io_out ? io_r_59_b : _GEN_148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_150 = 10'h3c == r_count_0_io_out ? io_r_60_b : _GEN_149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_151 = 10'h3d == r_count_0_io_out ? io_r_61_b : _GEN_150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_152 = 10'h3e == r_count_0_io_out ? io_r_62_b : _GEN_151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_153 = 10'h3f == r_count_0_io_out ? io_r_63_b : _GEN_152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_154 = 10'h40 == r_count_0_io_out ? io_r_64_b : _GEN_153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_155 = 10'h41 == r_count_0_io_out ? io_r_65_b : _GEN_154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_156 = 10'h42 == r_count_0_io_out ? io_r_66_b : _GEN_155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_157 = 10'h43 == r_count_0_io_out ? io_r_67_b : _GEN_156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_158 = 10'h44 == r_count_0_io_out ? io_r_68_b : _GEN_157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_159 = 10'h45 == r_count_0_io_out ? io_r_69_b : _GEN_158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_160 = 10'h46 == r_count_0_io_out ? io_r_70_b : _GEN_159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_161 = 10'h47 == r_count_0_io_out ? io_r_71_b : _GEN_160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_162 = 10'h48 == r_count_0_io_out ? io_r_72_b : _GEN_161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_163 = 10'h49 == r_count_0_io_out ? io_r_73_b : _GEN_162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_164 = 10'h4a == r_count_0_io_out ? io_r_74_b : _GEN_163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_165 = 10'h4b == r_count_0_io_out ? io_r_75_b : _GEN_164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_166 = 10'h4c == r_count_0_io_out ? io_r_76_b : _GEN_165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_167 = 10'h4d == r_count_0_io_out ? io_r_77_b : _GEN_166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_168 = 10'h4e == r_count_0_io_out ? io_r_78_b : _GEN_167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_169 = 10'h4f == r_count_0_io_out ? io_r_79_b : _GEN_168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_170 = 10'h50 == r_count_0_io_out ? io_r_80_b : _GEN_169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_171 = 10'h51 == r_count_0_io_out ? io_r_81_b : _GEN_170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_172 = 10'h52 == r_count_0_io_out ? io_r_82_b : _GEN_171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_173 = 10'h53 == r_count_0_io_out ? io_r_83_b : _GEN_172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_174 = 10'h54 == r_count_0_io_out ? io_r_84_b : _GEN_173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_175 = 10'h55 == r_count_0_io_out ? io_r_85_b : _GEN_174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_176 = 10'h56 == r_count_0_io_out ? io_r_86_b : _GEN_175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_177 = 10'h57 == r_count_0_io_out ? io_r_87_b : _GEN_176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_178 = 10'h58 == r_count_0_io_out ? io_r_88_b : _GEN_177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_179 = 10'h59 == r_count_0_io_out ? io_r_89_b : _GEN_178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_180 = 10'h5a == r_count_0_io_out ? io_r_90_b : _GEN_179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_181 = 10'h5b == r_count_0_io_out ? io_r_91_b : _GEN_180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_182 = 10'h5c == r_count_0_io_out ? io_r_92_b : _GEN_181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_183 = 10'h5d == r_count_0_io_out ? io_r_93_b : _GEN_182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_184 = 10'h5e == r_count_0_io_out ? io_r_94_b : _GEN_183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_185 = 10'h5f == r_count_0_io_out ? io_r_95_b : _GEN_184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_186 = 10'h60 == r_count_0_io_out ? io_r_96_b : _GEN_185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_187 = 10'h61 == r_count_0_io_out ? io_r_97_b : _GEN_186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_188 = 10'h62 == r_count_0_io_out ? io_r_98_b : _GEN_187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_189 = 10'h63 == r_count_0_io_out ? io_r_99_b : _GEN_188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_190 = 10'h64 == r_count_0_io_out ? io_r_100_b : _GEN_189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_191 = 10'h65 == r_count_0_io_out ? io_r_101_b : _GEN_190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_192 = 10'h66 == r_count_0_io_out ? io_r_102_b : _GEN_191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_193 = 10'h67 == r_count_0_io_out ? io_r_103_b : _GEN_192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_194 = 10'h68 == r_count_0_io_out ? io_r_104_b : _GEN_193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_195 = 10'h69 == r_count_0_io_out ? io_r_105_b : _GEN_194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_196 = 10'h6a == r_count_0_io_out ? io_r_106_b : _GEN_195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_197 = 10'h6b == r_count_0_io_out ? io_r_107_b : _GEN_196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_198 = 10'h6c == r_count_0_io_out ? io_r_108_b : _GEN_197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_199 = 10'h6d == r_count_0_io_out ? io_r_109_b : _GEN_198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_200 = 10'h6e == r_count_0_io_out ? io_r_110_b : _GEN_199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_201 = 10'h6f == r_count_0_io_out ? io_r_111_b : _GEN_200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_202 = 10'h70 == r_count_0_io_out ? io_r_112_b : _GEN_201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_203 = 10'h71 == r_count_0_io_out ? io_r_113_b : _GEN_202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_204 = 10'h72 == r_count_0_io_out ? io_r_114_b : _GEN_203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_205 = 10'h73 == r_count_0_io_out ? io_r_115_b : _GEN_204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_206 = 10'h74 == r_count_0_io_out ? io_r_116_b : _GEN_205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_207 = 10'h75 == r_count_0_io_out ? io_r_117_b : _GEN_206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_208 = 10'h76 == r_count_0_io_out ? io_r_118_b : _GEN_207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_209 = 10'h77 == r_count_0_io_out ? io_r_119_b : _GEN_208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_210 = 10'h78 == r_count_0_io_out ? io_r_120_b : _GEN_209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_211 = 10'h79 == r_count_0_io_out ? io_r_121_b : _GEN_210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_212 = 10'h7a == r_count_0_io_out ? io_r_122_b : _GEN_211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_213 = 10'h7b == r_count_0_io_out ? io_r_123_b : _GEN_212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_214 = 10'h7c == r_count_0_io_out ? io_r_124_b : _GEN_213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_215 = 10'h7d == r_count_0_io_out ? io_r_125_b : _GEN_214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_216 = 10'h7e == r_count_0_io_out ? io_r_126_b : _GEN_215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_217 = 10'h7f == r_count_0_io_out ? io_r_127_b : _GEN_216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_218 = 10'h80 == r_count_0_io_out ? io_r_128_b : _GEN_217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_219 = 10'h81 == r_count_0_io_out ? io_r_129_b : _GEN_218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_220 = 10'h82 == r_count_0_io_out ? io_r_130_b : _GEN_219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_221 = 10'h83 == r_count_0_io_out ? io_r_131_b : _GEN_220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_222 = 10'h84 == r_count_0_io_out ? io_r_132_b : _GEN_221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_223 = 10'h85 == r_count_0_io_out ? io_r_133_b : _GEN_222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_224 = 10'h86 == r_count_0_io_out ? io_r_134_b : _GEN_223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_225 = 10'h87 == r_count_0_io_out ? io_r_135_b : _GEN_224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_226 = 10'h88 == r_count_0_io_out ? io_r_136_b : _GEN_225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_227 = 10'h89 == r_count_0_io_out ? io_r_137_b : _GEN_226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_228 = 10'h8a == r_count_0_io_out ? io_r_138_b : _GEN_227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_229 = 10'h8b == r_count_0_io_out ? io_r_139_b : _GEN_228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_230 = 10'h8c == r_count_0_io_out ? io_r_140_b : _GEN_229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_231 = 10'h8d == r_count_0_io_out ? io_r_141_b : _GEN_230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_232 = 10'h8e == r_count_0_io_out ? io_r_142_b : _GEN_231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_233 = 10'h8f == r_count_0_io_out ? io_r_143_b : _GEN_232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_234 = 10'h90 == r_count_0_io_out ? io_r_144_b : _GEN_233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_235 = 10'h91 == r_count_0_io_out ? io_r_145_b : _GEN_234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_236 = 10'h92 == r_count_0_io_out ? io_r_146_b : _GEN_235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_237 = 10'h93 == r_count_0_io_out ? io_r_147_b : _GEN_236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_238 = 10'h94 == r_count_0_io_out ? io_r_148_b : _GEN_237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_239 = 10'h95 == r_count_0_io_out ? io_r_149_b : _GEN_238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_240 = 10'h96 == r_count_0_io_out ? io_r_150_b : _GEN_239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_241 = 10'h97 == r_count_0_io_out ? io_r_151_b : _GEN_240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_242 = 10'h98 == r_count_0_io_out ? io_r_152_b : _GEN_241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_243 = 10'h99 == r_count_0_io_out ? io_r_153_b : _GEN_242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_244 = 10'h9a == r_count_0_io_out ? io_r_154_b : _GEN_243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_245 = 10'h9b == r_count_0_io_out ? io_r_155_b : _GEN_244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_246 = 10'h9c == r_count_0_io_out ? io_r_156_b : _GEN_245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_247 = 10'h9d == r_count_0_io_out ? io_r_157_b : _GEN_246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_248 = 10'h9e == r_count_0_io_out ? io_r_158_b : _GEN_247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_249 = 10'h9f == r_count_0_io_out ? io_r_159_b : _GEN_248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_250 = 10'ha0 == r_count_0_io_out ? io_r_160_b : _GEN_249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_251 = 10'ha1 == r_count_0_io_out ? io_r_161_b : _GEN_250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_252 = 10'ha2 == r_count_0_io_out ? io_r_162_b : _GEN_251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_253 = 10'ha3 == r_count_0_io_out ? io_r_163_b : _GEN_252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_254 = 10'ha4 == r_count_0_io_out ? io_r_164_b : _GEN_253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_255 = 10'ha5 == r_count_0_io_out ? io_r_165_b : _GEN_254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_256 = 10'ha6 == r_count_0_io_out ? io_r_166_b : _GEN_255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_257 = 10'ha7 == r_count_0_io_out ? io_r_167_b : _GEN_256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_258 = 10'ha8 == r_count_0_io_out ? io_r_168_b : _GEN_257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_259 = 10'ha9 == r_count_0_io_out ? io_r_169_b : _GEN_258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_260 = 10'haa == r_count_0_io_out ? io_r_170_b : _GEN_259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_261 = 10'hab == r_count_0_io_out ? io_r_171_b : _GEN_260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_262 = 10'hac == r_count_0_io_out ? io_r_172_b : _GEN_261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_263 = 10'had == r_count_0_io_out ? io_r_173_b : _GEN_262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_264 = 10'hae == r_count_0_io_out ? io_r_174_b : _GEN_263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_265 = 10'haf == r_count_0_io_out ? io_r_175_b : _GEN_264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_266 = 10'hb0 == r_count_0_io_out ? io_r_176_b : _GEN_265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_267 = 10'hb1 == r_count_0_io_out ? io_r_177_b : _GEN_266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_268 = 10'hb2 == r_count_0_io_out ? io_r_178_b : _GEN_267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_269 = 10'hb3 == r_count_0_io_out ? io_r_179_b : _GEN_268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_270 = 10'hb4 == r_count_0_io_out ? io_r_180_b : _GEN_269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_271 = 10'hb5 == r_count_0_io_out ? io_r_181_b : _GEN_270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_272 = 10'hb6 == r_count_0_io_out ? io_r_182_b : _GEN_271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_273 = 10'hb7 == r_count_0_io_out ? io_r_183_b : _GEN_272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_274 = 10'hb8 == r_count_0_io_out ? io_r_184_b : _GEN_273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_275 = 10'hb9 == r_count_0_io_out ? io_r_185_b : _GEN_274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_276 = 10'hba == r_count_0_io_out ? io_r_186_b : _GEN_275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_277 = 10'hbb == r_count_0_io_out ? io_r_187_b : _GEN_276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_278 = 10'hbc == r_count_0_io_out ? io_r_188_b : _GEN_277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_279 = 10'hbd == r_count_0_io_out ? io_r_189_b : _GEN_278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_280 = 10'hbe == r_count_0_io_out ? io_r_190_b : _GEN_279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_281 = 10'hbf == r_count_0_io_out ? io_r_191_b : _GEN_280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_282 = 10'hc0 == r_count_0_io_out ? io_r_192_b : _GEN_281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_283 = 10'hc1 == r_count_0_io_out ? io_r_193_b : _GEN_282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_284 = 10'hc2 == r_count_0_io_out ? io_r_194_b : _GEN_283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_285 = 10'hc3 == r_count_0_io_out ? io_r_195_b : _GEN_284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_286 = 10'hc4 == r_count_0_io_out ? io_r_196_b : _GEN_285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_287 = 10'hc5 == r_count_0_io_out ? io_r_197_b : _GEN_286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_288 = 10'hc6 == r_count_0_io_out ? io_r_198_b : _GEN_287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_289 = 10'hc7 == r_count_0_io_out ? io_r_199_b : _GEN_288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_290 = 10'hc8 == r_count_0_io_out ? io_r_200_b : _GEN_289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_291 = 10'hc9 == r_count_0_io_out ? io_r_201_b : _GEN_290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_292 = 10'hca == r_count_0_io_out ? io_r_202_b : _GEN_291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_293 = 10'hcb == r_count_0_io_out ? io_r_203_b : _GEN_292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_294 = 10'hcc == r_count_0_io_out ? io_r_204_b : _GEN_293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_295 = 10'hcd == r_count_0_io_out ? io_r_205_b : _GEN_294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_296 = 10'hce == r_count_0_io_out ? io_r_206_b : _GEN_295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_297 = 10'hcf == r_count_0_io_out ? io_r_207_b : _GEN_296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_298 = 10'hd0 == r_count_0_io_out ? io_r_208_b : _GEN_297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_299 = 10'hd1 == r_count_0_io_out ? io_r_209_b : _GEN_298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_300 = 10'hd2 == r_count_0_io_out ? io_r_210_b : _GEN_299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_301 = 10'hd3 == r_count_0_io_out ? io_r_211_b : _GEN_300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_302 = 10'hd4 == r_count_0_io_out ? io_r_212_b : _GEN_301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_303 = 10'hd5 == r_count_0_io_out ? io_r_213_b : _GEN_302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_304 = 10'hd6 == r_count_0_io_out ? io_r_214_b : _GEN_303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_305 = 10'hd7 == r_count_0_io_out ? io_r_215_b : _GEN_304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_306 = 10'hd8 == r_count_0_io_out ? io_r_216_b : _GEN_305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_307 = 10'hd9 == r_count_0_io_out ? io_r_217_b : _GEN_306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_308 = 10'hda == r_count_0_io_out ? io_r_218_b : _GEN_307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_309 = 10'hdb == r_count_0_io_out ? io_r_219_b : _GEN_308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_310 = 10'hdc == r_count_0_io_out ? io_r_220_b : _GEN_309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_311 = 10'hdd == r_count_0_io_out ? io_r_221_b : _GEN_310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_312 = 10'hde == r_count_0_io_out ? io_r_222_b : _GEN_311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_313 = 10'hdf == r_count_0_io_out ? io_r_223_b : _GEN_312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_314 = 10'he0 == r_count_0_io_out ? io_r_224_b : _GEN_313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_315 = 10'he1 == r_count_0_io_out ? io_r_225_b : _GEN_314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_316 = 10'he2 == r_count_0_io_out ? io_r_226_b : _GEN_315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_317 = 10'he3 == r_count_0_io_out ? io_r_227_b : _GEN_316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_318 = 10'he4 == r_count_0_io_out ? io_r_228_b : _GEN_317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_319 = 10'he5 == r_count_0_io_out ? io_r_229_b : _GEN_318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_320 = 10'he6 == r_count_0_io_out ? io_r_230_b : _GEN_319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_321 = 10'he7 == r_count_0_io_out ? io_r_231_b : _GEN_320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_322 = 10'he8 == r_count_0_io_out ? io_r_232_b : _GEN_321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_323 = 10'he9 == r_count_0_io_out ? io_r_233_b : _GEN_322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_324 = 10'hea == r_count_0_io_out ? io_r_234_b : _GEN_323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_325 = 10'heb == r_count_0_io_out ? io_r_235_b : _GEN_324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_326 = 10'hec == r_count_0_io_out ? io_r_236_b : _GEN_325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_327 = 10'hed == r_count_0_io_out ? io_r_237_b : _GEN_326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_328 = 10'hee == r_count_0_io_out ? io_r_238_b : _GEN_327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_329 = 10'hef == r_count_0_io_out ? io_r_239_b : _GEN_328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_330 = 10'hf0 == r_count_0_io_out ? io_r_240_b : _GEN_329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_331 = 10'hf1 == r_count_0_io_out ? io_r_241_b : _GEN_330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_332 = 10'hf2 == r_count_0_io_out ? io_r_242_b : _GEN_331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_333 = 10'hf3 == r_count_0_io_out ? io_r_243_b : _GEN_332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_334 = 10'hf4 == r_count_0_io_out ? io_r_244_b : _GEN_333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_335 = 10'hf5 == r_count_0_io_out ? io_r_245_b : _GEN_334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_336 = 10'hf6 == r_count_0_io_out ? io_r_246_b : _GEN_335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_337 = 10'hf7 == r_count_0_io_out ? io_r_247_b : _GEN_336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_338 = 10'hf8 == r_count_0_io_out ? io_r_248_b : _GEN_337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_339 = 10'hf9 == r_count_0_io_out ? io_r_249_b : _GEN_338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_340 = 10'hfa == r_count_0_io_out ? io_r_250_b : _GEN_339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_341 = 10'hfb == r_count_0_io_out ? io_r_251_b : _GEN_340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_342 = 10'hfc == r_count_0_io_out ? io_r_252_b : _GEN_341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_343 = 10'hfd == r_count_0_io_out ? io_r_253_b : _GEN_342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_344 = 10'hfe == r_count_0_io_out ? io_r_254_b : _GEN_343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_345 = 10'hff == r_count_0_io_out ? io_r_255_b : _GEN_344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_346 = 10'h100 == r_count_0_io_out ? io_r_256_b : _GEN_345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_347 = 10'h101 == r_count_0_io_out ? io_r_257_b : _GEN_346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_348 = 10'h102 == r_count_0_io_out ? io_r_258_b : _GEN_347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_349 = 10'h103 == r_count_0_io_out ? io_r_259_b : _GEN_348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_350 = 10'h104 == r_count_0_io_out ? io_r_260_b : _GEN_349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_351 = 10'h105 == r_count_0_io_out ? io_r_261_b : _GEN_350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_352 = 10'h106 == r_count_0_io_out ? io_r_262_b : _GEN_351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_353 = 10'h107 == r_count_0_io_out ? io_r_263_b : _GEN_352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_354 = 10'h108 == r_count_0_io_out ? io_r_264_b : _GEN_353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_355 = 10'h109 == r_count_0_io_out ? io_r_265_b : _GEN_354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_356 = 10'h10a == r_count_0_io_out ? io_r_266_b : _GEN_355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_357 = 10'h10b == r_count_0_io_out ? io_r_267_b : _GEN_356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_358 = 10'h10c == r_count_0_io_out ? io_r_268_b : _GEN_357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_359 = 10'h10d == r_count_0_io_out ? io_r_269_b : _GEN_358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_360 = 10'h10e == r_count_0_io_out ? io_r_270_b : _GEN_359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_361 = 10'h10f == r_count_0_io_out ? io_r_271_b : _GEN_360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_362 = 10'h110 == r_count_0_io_out ? io_r_272_b : _GEN_361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_363 = 10'h111 == r_count_0_io_out ? io_r_273_b : _GEN_362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_364 = 10'h112 == r_count_0_io_out ? io_r_274_b : _GEN_363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_365 = 10'h113 == r_count_0_io_out ? io_r_275_b : _GEN_364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_366 = 10'h114 == r_count_0_io_out ? io_r_276_b : _GEN_365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_367 = 10'h115 == r_count_0_io_out ? io_r_277_b : _GEN_366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_368 = 10'h116 == r_count_0_io_out ? io_r_278_b : _GEN_367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_369 = 10'h117 == r_count_0_io_out ? io_r_279_b : _GEN_368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_370 = 10'h118 == r_count_0_io_out ? io_r_280_b : _GEN_369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_371 = 10'h119 == r_count_0_io_out ? io_r_281_b : _GEN_370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_372 = 10'h11a == r_count_0_io_out ? io_r_282_b : _GEN_371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_373 = 10'h11b == r_count_0_io_out ? io_r_283_b : _GEN_372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_374 = 10'h11c == r_count_0_io_out ? io_r_284_b : _GEN_373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_375 = 10'h11d == r_count_0_io_out ? io_r_285_b : _GEN_374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_376 = 10'h11e == r_count_0_io_out ? io_r_286_b : _GEN_375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_377 = 10'h11f == r_count_0_io_out ? io_r_287_b : _GEN_376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_378 = 10'h120 == r_count_0_io_out ? io_r_288_b : _GEN_377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_379 = 10'h121 == r_count_0_io_out ? io_r_289_b : _GEN_378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_380 = 10'h122 == r_count_0_io_out ? io_r_290_b : _GEN_379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_381 = 10'h123 == r_count_0_io_out ? io_r_291_b : _GEN_380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_382 = 10'h124 == r_count_0_io_out ? io_r_292_b : _GEN_381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_383 = 10'h125 == r_count_0_io_out ? io_r_293_b : _GEN_382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_384 = 10'h126 == r_count_0_io_out ? io_r_294_b : _GEN_383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_385 = 10'h127 == r_count_0_io_out ? io_r_295_b : _GEN_384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_386 = 10'h128 == r_count_0_io_out ? io_r_296_b : _GEN_385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_387 = 10'h129 == r_count_0_io_out ? io_r_297_b : _GEN_386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_388 = 10'h12a == r_count_0_io_out ? io_r_298_b : _GEN_387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_389 = 10'h12b == r_count_0_io_out ? io_r_299_b : _GEN_388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_390 = 10'h12c == r_count_0_io_out ? io_r_300_b : _GEN_389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_391 = 10'h12d == r_count_0_io_out ? io_r_301_b : _GEN_390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_392 = 10'h12e == r_count_0_io_out ? io_r_302_b : _GEN_391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_393 = 10'h12f == r_count_0_io_out ? io_r_303_b : _GEN_392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_394 = 10'h130 == r_count_0_io_out ? io_r_304_b : _GEN_393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_395 = 10'h131 == r_count_0_io_out ? io_r_305_b : _GEN_394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_396 = 10'h132 == r_count_0_io_out ? io_r_306_b : _GEN_395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_397 = 10'h133 == r_count_0_io_out ? io_r_307_b : _GEN_396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_398 = 10'h134 == r_count_0_io_out ? io_r_308_b : _GEN_397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_399 = 10'h135 == r_count_0_io_out ? io_r_309_b : _GEN_398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_400 = 10'h136 == r_count_0_io_out ? io_r_310_b : _GEN_399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_401 = 10'h137 == r_count_0_io_out ? io_r_311_b : _GEN_400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_402 = 10'h138 == r_count_0_io_out ? io_r_312_b : _GEN_401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_403 = 10'h139 == r_count_0_io_out ? io_r_313_b : _GEN_402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_404 = 10'h13a == r_count_0_io_out ? io_r_314_b : _GEN_403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_405 = 10'h13b == r_count_0_io_out ? io_r_315_b : _GEN_404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_406 = 10'h13c == r_count_0_io_out ? io_r_316_b : _GEN_405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_407 = 10'h13d == r_count_0_io_out ? io_r_317_b : _GEN_406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_408 = 10'h13e == r_count_0_io_out ? io_r_318_b : _GEN_407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_409 = 10'h13f == r_count_0_io_out ? io_r_319_b : _GEN_408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_410 = 10'h140 == r_count_0_io_out ? io_r_320_b : _GEN_409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_411 = 10'h141 == r_count_0_io_out ? io_r_321_b : _GEN_410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_412 = 10'h142 == r_count_0_io_out ? io_r_322_b : _GEN_411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_413 = 10'h143 == r_count_0_io_out ? io_r_323_b : _GEN_412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_414 = 10'h144 == r_count_0_io_out ? io_r_324_b : _GEN_413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_415 = 10'h145 == r_count_0_io_out ? io_r_325_b : _GEN_414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_416 = 10'h146 == r_count_0_io_out ? io_r_326_b : _GEN_415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_417 = 10'h147 == r_count_0_io_out ? io_r_327_b : _GEN_416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_418 = 10'h148 == r_count_0_io_out ? io_r_328_b : _GEN_417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_419 = 10'h149 == r_count_0_io_out ? io_r_329_b : _GEN_418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_420 = 10'h14a == r_count_0_io_out ? io_r_330_b : _GEN_419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_421 = 10'h14b == r_count_0_io_out ? io_r_331_b : _GEN_420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_422 = 10'h14c == r_count_0_io_out ? io_r_332_b : _GEN_421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_423 = 10'h14d == r_count_0_io_out ? io_r_333_b : _GEN_422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_424 = 10'h14e == r_count_0_io_out ? io_r_334_b : _GEN_423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_425 = 10'h14f == r_count_0_io_out ? io_r_335_b : _GEN_424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_426 = 10'h150 == r_count_0_io_out ? io_r_336_b : _GEN_425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_427 = 10'h151 == r_count_0_io_out ? io_r_337_b : _GEN_426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_428 = 10'h152 == r_count_0_io_out ? io_r_338_b : _GEN_427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_429 = 10'h153 == r_count_0_io_out ? io_r_339_b : _GEN_428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_430 = 10'h154 == r_count_0_io_out ? io_r_340_b : _GEN_429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_431 = 10'h155 == r_count_0_io_out ? io_r_341_b : _GEN_430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_432 = 10'h156 == r_count_0_io_out ? io_r_342_b : _GEN_431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_433 = 10'h157 == r_count_0_io_out ? io_r_343_b : _GEN_432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_434 = 10'h158 == r_count_0_io_out ? io_r_344_b : _GEN_433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_435 = 10'h159 == r_count_0_io_out ? io_r_345_b : _GEN_434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_436 = 10'h15a == r_count_0_io_out ? io_r_346_b : _GEN_435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_437 = 10'h15b == r_count_0_io_out ? io_r_347_b : _GEN_436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_438 = 10'h15c == r_count_0_io_out ? io_r_348_b : _GEN_437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_439 = 10'h15d == r_count_0_io_out ? io_r_349_b : _GEN_438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_440 = 10'h15e == r_count_0_io_out ? io_r_350_b : _GEN_439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_441 = 10'h15f == r_count_0_io_out ? io_r_351_b : _GEN_440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_442 = 10'h160 == r_count_0_io_out ? io_r_352_b : _GEN_441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_443 = 10'h161 == r_count_0_io_out ? io_r_353_b : _GEN_442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_444 = 10'h162 == r_count_0_io_out ? io_r_354_b : _GEN_443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_445 = 10'h163 == r_count_0_io_out ? io_r_355_b : _GEN_444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_446 = 10'h164 == r_count_0_io_out ? io_r_356_b : _GEN_445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_447 = 10'h165 == r_count_0_io_out ? io_r_357_b : _GEN_446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_448 = 10'h166 == r_count_0_io_out ? io_r_358_b : _GEN_447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_449 = 10'h167 == r_count_0_io_out ? io_r_359_b : _GEN_448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_450 = 10'h168 == r_count_0_io_out ? io_r_360_b : _GEN_449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_451 = 10'h169 == r_count_0_io_out ? io_r_361_b : _GEN_450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_452 = 10'h16a == r_count_0_io_out ? io_r_362_b : _GEN_451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_453 = 10'h16b == r_count_0_io_out ? io_r_363_b : _GEN_452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_454 = 10'h16c == r_count_0_io_out ? io_r_364_b : _GEN_453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_455 = 10'h16d == r_count_0_io_out ? io_r_365_b : _GEN_454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_456 = 10'h16e == r_count_0_io_out ? io_r_366_b : _GEN_455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_457 = 10'h16f == r_count_0_io_out ? io_r_367_b : _GEN_456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_458 = 10'h170 == r_count_0_io_out ? io_r_368_b : _GEN_457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_459 = 10'h171 == r_count_0_io_out ? io_r_369_b : _GEN_458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_460 = 10'h172 == r_count_0_io_out ? io_r_370_b : _GEN_459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_461 = 10'h173 == r_count_0_io_out ? io_r_371_b : _GEN_460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_462 = 10'h174 == r_count_0_io_out ? io_r_372_b : _GEN_461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_463 = 10'h175 == r_count_0_io_out ? io_r_373_b : _GEN_462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_464 = 10'h176 == r_count_0_io_out ? io_r_374_b : _GEN_463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_465 = 10'h177 == r_count_0_io_out ? io_r_375_b : _GEN_464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_466 = 10'h178 == r_count_0_io_out ? io_r_376_b : _GEN_465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_467 = 10'h179 == r_count_0_io_out ? io_r_377_b : _GEN_466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_468 = 10'h17a == r_count_0_io_out ? io_r_378_b : _GEN_467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_469 = 10'h17b == r_count_0_io_out ? io_r_379_b : _GEN_468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_470 = 10'h17c == r_count_0_io_out ? io_r_380_b : _GEN_469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_471 = 10'h17d == r_count_0_io_out ? io_r_381_b : _GEN_470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_472 = 10'h17e == r_count_0_io_out ? io_r_382_b : _GEN_471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_473 = 10'h17f == r_count_0_io_out ? io_r_383_b : _GEN_472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_474 = 10'h180 == r_count_0_io_out ? io_r_384_b : _GEN_473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_475 = 10'h181 == r_count_0_io_out ? io_r_385_b : _GEN_474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_476 = 10'h182 == r_count_0_io_out ? io_r_386_b : _GEN_475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_477 = 10'h183 == r_count_0_io_out ? io_r_387_b : _GEN_476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_478 = 10'h184 == r_count_0_io_out ? io_r_388_b : _GEN_477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_479 = 10'h185 == r_count_0_io_out ? io_r_389_b : _GEN_478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_480 = 10'h186 == r_count_0_io_out ? io_r_390_b : _GEN_479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_481 = 10'h187 == r_count_0_io_out ? io_r_391_b : _GEN_480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_482 = 10'h188 == r_count_0_io_out ? io_r_392_b : _GEN_481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_483 = 10'h189 == r_count_0_io_out ? io_r_393_b : _GEN_482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_484 = 10'h18a == r_count_0_io_out ? io_r_394_b : _GEN_483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_485 = 10'h18b == r_count_0_io_out ? io_r_395_b : _GEN_484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_486 = 10'h18c == r_count_0_io_out ? io_r_396_b : _GEN_485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_487 = 10'h18d == r_count_0_io_out ? io_r_397_b : _GEN_486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_488 = 10'h18e == r_count_0_io_out ? io_r_398_b : _GEN_487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_489 = 10'h18f == r_count_0_io_out ? io_r_399_b : _GEN_488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_490 = 10'h190 == r_count_0_io_out ? io_r_400_b : _GEN_489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_491 = 10'h191 == r_count_0_io_out ? io_r_401_b : _GEN_490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_492 = 10'h192 == r_count_0_io_out ? io_r_402_b : _GEN_491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_493 = 10'h193 == r_count_0_io_out ? io_r_403_b : _GEN_492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_494 = 10'h194 == r_count_0_io_out ? io_r_404_b : _GEN_493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_495 = 10'h195 == r_count_0_io_out ? io_r_405_b : _GEN_494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_496 = 10'h196 == r_count_0_io_out ? io_r_406_b : _GEN_495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_497 = 10'h197 == r_count_0_io_out ? io_r_407_b : _GEN_496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_498 = 10'h198 == r_count_0_io_out ? io_r_408_b : _GEN_497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_499 = 10'h199 == r_count_0_io_out ? io_r_409_b : _GEN_498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_500 = 10'h19a == r_count_0_io_out ? io_r_410_b : _GEN_499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_501 = 10'h19b == r_count_0_io_out ? io_r_411_b : _GEN_500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_502 = 10'h19c == r_count_0_io_out ? io_r_412_b : _GEN_501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_503 = 10'h19d == r_count_0_io_out ? io_r_413_b : _GEN_502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_504 = 10'h19e == r_count_0_io_out ? io_r_414_b : _GEN_503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_505 = 10'h19f == r_count_0_io_out ? io_r_415_b : _GEN_504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_506 = 10'h1a0 == r_count_0_io_out ? io_r_416_b : _GEN_505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_507 = 10'h1a1 == r_count_0_io_out ? io_r_417_b : _GEN_506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_508 = 10'h1a2 == r_count_0_io_out ? io_r_418_b : _GEN_507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_509 = 10'h1a3 == r_count_0_io_out ? io_r_419_b : _GEN_508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_510 = 10'h1a4 == r_count_0_io_out ? io_r_420_b : _GEN_509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_511 = 10'h1a5 == r_count_0_io_out ? io_r_421_b : _GEN_510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_512 = 10'h1a6 == r_count_0_io_out ? io_r_422_b : _GEN_511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_513 = 10'h1a7 == r_count_0_io_out ? io_r_423_b : _GEN_512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_514 = 10'h1a8 == r_count_0_io_out ? io_r_424_b : _GEN_513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_515 = 10'h1a9 == r_count_0_io_out ? io_r_425_b : _GEN_514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_516 = 10'h1aa == r_count_0_io_out ? io_r_426_b : _GEN_515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_517 = 10'h1ab == r_count_0_io_out ? io_r_427_b : _GEN_516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_518 = 10'h1ac == r_count_0_io_out ? io_r_428_b : _GEN_517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_519 = 10'h1ad == r_count_0_io_out ? io_r_429_b : _GEN_518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_520 = 10'h1ae == r_count_0_io_out ? io_r_430_b : _GEN_519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_521 = 10'h1af == r_count_0_io_out ? io_r_431_b : _GEN_520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_522 = 10'h1b0 == r_count_0_io_out ? io_r_432_b : _GEN_521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_523 = 10'h1b1 == r_count_0_io_out ? io_r_433_b : _GEN_522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_524 = 10'h1b2 == r_count_0_io_out ? io_r_434_b : _GEN_523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_525 = 10'h1b3 == r_count_0_io_out ? io_r_435_b : _GEN_524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_526 = 10'h1b4 == r_count_0_io_out ? io_r_436_b : _GEN_525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_527 = 10'h1b5 == r_count_0_io_out ? io_r_437_b : _GEN_526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_528 = 10'h1b6 == r_count_0_io_out ? io_r_438_b : _GEN_527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_529 = 10'h1b7 == r_count_0_io_out ? io_r_439_b : _GEN_528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_530 = 10'h1b8 == r_count_0_io_out ? io_r_440_b : _GEN_529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_531 = 10'h1b9 == r_count_0_io_out ? io_r_441_b : _GEN_530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_532 = 10'h1ba == r_count_0_io_out ? io_r_442_b : _GEN_531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_533 = 10'h1bb == r_count_0_io_out ? io_r_443_b : _GEN_532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_534 = 10'h1bc == r_count_0_io_out ? io_r_444_b : _GEN_533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_535 = 10'h1bd == r_count_0_io_out ? io_r_445_b : _GEN_534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_536 = 10'h1be == r_count_0_io_out ? io_r_446_b : _GEN_535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_537 = 10'h1bf == r_count_0_io_out ? io_r_447_b : _GEN_536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_538 = 10'h1c0 == r_count_0_io_out ? io_r_448_b : _GEN_537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_539 = 10'h1c1 == r_count_0_io_out ? io_r_449_b : _GEN_538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_540 = 10'h1c2 == r_count_0_io_out ? io_r_450_b : _GEN_539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_541 = 10'h1c3 == r_count_0_io_out ? io_r_451_b : _GEN_540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_542 = 10'h1c4 == r_count_0_io_out ? io_r_452_b : _GEN_541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_543 = 10'h1c5 == r_count_0_io_out ? io_r_453_b : _GEN_542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_544 = 10'h1c6 == r_count_0_io_out ? io_r_454_b : _GEN_543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_545 = 10'h1c7 == r_count_0_io_out ? io_r_455_b : _GEN_544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_546 = 10'h1c8 == r_count_0_io_out ? io_r_456_b : _GEN_545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_547 = 10'h1c9 == r_count_0_io_out ? io_r_457_b : _GEN_546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_548 = 10'h1ca == r_count_0_io_out ? io_r_458_b : _GEN_547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_549 = 10'h1cb == r_count_0_io_out ? io_r_459_b : _GEN_548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_550 = 10'h1cc == r_count_0_io_out ? io_r_460_b : _GEN_549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_551 = 10'h1cd == r_count_0_io_out ? io_r_461_b : _GEN_550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_552 = 10'h1ce == r_count_0_io_out ? io_r_462_b : _GEN_551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_553 = 10'h1cf == r_count_0_io_out ? io_r_463_b : _GEN_552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_554 = 10'h1d0 == r_count_0_io_out ? io_r_464_b : _GEN_553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_555 = 10'h1d1 == r_count_0_io_out ? io_r_465_b : _GEN_554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_556 = 10'h1d2 == r_count_0_io_out ? io_r_466_b : _GEN_555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_557 = 10'h1d3 == r_count_0_io_out ? io_r_467_b : _GEN_556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_558 = 10'h1d4 == r_count_0_io_out ? io_r_468_b : _GEN_557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_559 = 10'h1d5 == r_count_0_io_out ? io_r_469_b : _GEN_558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_560 = 10'h1d6 == r_count_0_io_out ? io_r_470_b : _GEN_559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_561 = 10'h1d7 == r_count_0_io_out ? io_r_471_b : _GEN_560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_562 = 10'h1d8 == r_count_0_io_out ? io_r_472_b : _GEN_561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_563 = 10'h1d9 == r_count_0_io_out ? io_r_473_b : _GEN_562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_564 = 10'h1da == r_count_0_io_out ? io_r_474_b : _GEN_563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_565 = 10'h1db == r_count_0_io_out ? io_r_475_b : _GEN_564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_566 = 10'h1dc == r_count_0_io_out ? io_r_476_b : _GEN_565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_567 = 10'h1dd == r_count_0_io_out ? io_r_477_b : _GEN_566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_568 = 10'h1de == r_count_0_io_out ? io_r_478_b : _GEN_567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_569 = 10'h1df == r_count_0_io_out ? io_r_479_b : _GEN_568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_570 = 10'h1e0 == r_count_0_io_out ? io_r_480_b : _GEN_569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_571 = 10'h1e1 == r_count_0_io_out ? io_r_481_b : _GEN_570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_572 = 10'h1e2 == r_count_0_io_out ? io_r_482_b : _GEN_571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_573 = 10'h1e3 == r_count_0_io_out ? io_r_483_b : _GEN_572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_574 = 10'h1e4 == r_count_0_io_out ? io_r_484_b : _GEN_573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_575 = 10'h1e5 == r_count_0_io_out ? io_r_485_b : _GEN_574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_576 = 10'h1e6 == r_count_0_io_out ? io_r_486_b : _GEN_575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_577 = 10'h1e7 == r_count_0_io_out ? io_r_487_b : _GEN_576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_578 = 10'h1e8 == r_count_0_io_out ? io_r_488_b : _GEN_577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_579 = 10'h1e9 == r_count_0_io_out ? io_r_489_b : _GEN_578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_580 = 10'h1ea == r_count_0_io_out ? io_r_490_b : _GEN_579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_581 = 10'h1eb == r_count_0_io_out ? io_r_491_b : _GEN_580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_582 = 10'h1ec == r_count_0_io_out ? io_r_492_b : _GEN_581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_583 = 10'h1ed == r_count_0_io_out ? io_r_493_b : _GEN_582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_584 = 10'h1ee == r_count_0_io_out ? io_r_494_b : _GEN_583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_585 = 10'h1ef == r_count_0_io_out ? io_r_495_b : _GEN_584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_586 = 10'h1f0 == r_count_0_io_out ? io_r_496_b : _GEN_585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_587 = 10'h1f1 == r_count_0_io_out ? io_r_497_b : _GEN_586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_588 = 10'h1f2 == r_count_0_io_out ? io_r_498_b : _GEN_587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_589 = 10'h1f3 == r_count_0_io_out ? io_r_499_b : _GEN_588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_590 = 10'h1f4 == r_count_0_io_out ? io_r_500_b : _GEN_589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_591 = 10'h1f5 == r_count_0_io_out ? io_r_501_b : _GEN_590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_592 = 10'h1f6 == r_count_0_io_out ? io_r_502_b : _GEN_591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_593 = 10'h1f7 == r_count_0_io_out ? io_r_503_b : _GEN_592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_594 = 10'h1f8 == r_count_0_io_out ? io_r_504_b : _GEN_593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_595 = 10'h1f9 == r_count_0_io_out ? io_r_505_b : _GEN_594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_596 = 10'h1fa == r_count_0_io_out ? io_r_506_b : _GEN_595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_597 = 10'h1fb == r_count_0_io_out ? io_r_507_b : _GEN_596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_598 = 10'h1fc == r_count_0_io_out ? io_r_508_b : _GEN_597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_599 = 10'h1fd == r_count_0_io_out ? io_r_509_b : _GEN_598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_600 = 10'h1fe == r_count_0_io_out ? io_r_510_b : _GEN_599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_601 = 10'h1ff == r_count_0_io_out ? io_r_511_b : _GEN_600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_602 = 10'h200 == r_count_0_io_out ? io_r_512_b : _GEN_601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_603 = 10'h201 == r_count_0_io_out ? io_r_513_b : _GEN_602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_604 = 10'h202 == r_count_0_io_out ? io_r_514_b : _GEN_603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_605 = 10'h203 == r_count_0_io_out ? io_r_515_b : _GEN_604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_606 = 10'h204 == r_count_0_io_out ? io_r_516_b : _GEN_605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_607 = 10'h205 == r_count_0_io_out ? io_r_517_b : _GEN_606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_608 = 10'h206 == r_count_0_io_out ? io_r_518_b : _GEN_607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_609 = 10'h207 == r_count_0_io_out ? io_r_519_b : _GEN_608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_610 = 10'h208 == r_count_0_io_out ? io_r_520_b : _GEN_609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_611 = 10'h209 == r_count_0_io_out ? io_r_521_b : _GEN_610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_612 = 10'h20a == r_count_0_io_out ? io_r_522_b : _GEN_611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_613 = 10'h20b == r_count_0_io_out ? io_r_523_b : _GEN_612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_614 = 10'h20c == r_count_0_io_out ? io_r_524_b : _GEN_613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_615 = 10'h20d == r_count_0_io_out ? io_r_525_b : _GEN_614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_616 = 10'h20e == r_count_0_io_out ? io_r_526_b : _GEN_615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_617 = 10'h20f == r_count_0_io_out ? io_r_527_b : _GEN_616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_618 = 10'h210 == r_count_0_io_out ? io_r_528_b : _GEN_617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_619 = 10'h211 == r_count_0_io_out ? io_r_529_b : _GEN_618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_620 = 10'h212 == r_count_0_io_out ? io_r_530_b : _GEN_619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_621 = 10'h213 == r_count_0_io_out ? io_r_531_b : _GEN_620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_622 = 10'h214 == r_count_0_io_out ? io_r_532_b : _GEN_621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_623 = 10'h215 == r_count_0_io_out ? io_r_533_b : _GEN_622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_624 = 10'h216 == r_count_0_io_out ? io_r_534_b : _GEN_623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_625 = 10'h217 == r_count_0_io_out ? io_r_535_b : _GEN_624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_626 = 10'h218 == r_count_0_io_out ? io_r_536_b : _GEN_625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_627 = 10'h219 == r_count_0_io_out ? io_r_537_b : _GEN_626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_628 = 10'h21a == r_count_0_io_out ? io_r_538_b : _GEN_627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_629 = 10'h21b == r_count_0_io_out ? io_r_539_b : _GEN_628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_630 = 10'h21c == r_count_0_io_out ? io_r_540_b : _GEN_629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_631 = 10'h21d == r_count_0_io_out ? io_r_541_b : _GEN_630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_632 = 10'h21e == r_count_0_io_out ? io_r_542_b : _GEN_631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_633 = 10'h21f == r_count_0_io_out ? io_r_543_b : _GEN_632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_634 = 10'h220 == r_count_0_io_out ? io_r_544_b : _GEN_633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_635 = 10'h221 == r_count_0_io_out ? io_r_545_b : _GEN_634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_636 = 10'h222 == r_count_0_io_out ? io_r_546_b : _GEN_635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_637 = 10'h223 == r_count_0_io_out ? io_r_547_b : _GEN_636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_638 = 10'h224 == r_count_0_io_out ? io_r_548_b : _GEN_637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_639 = 10'h225 == r_count_0_io_out ? io_r_549_b : _GEN_638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_640 = 10'h226 == r_count_0_io_out ? io_r_550_b : _GEN_639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_641 = 10'h227 == r_count_0_io_out ? io_r_551_b : _GEN_640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_642 = 10'h228 == r_count_0_io_out ? io_r_552_b : _GEN_641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_643 = 10'h229 == r_count_0_io_out ? io_r_553_b : _GEN_642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_644 = 10'h22a == r_count_0_io_out ? io_r_554_b : _GEN_643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_645 = 10'h22b == r_count_0_io_out ? io_r_555_b : _GEN_644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_646 = 10'h22c == r_count_0_io_out ? io_r_556_b : _GEN_645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_647 = 10'h22d == r_count_0_io_out ? io_r_557_b : _GEN_646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_648 = 10'h22e == r_count_0_io_out ? io_r_558_b : _GEN_647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_649 = 10'h22f == r_count_0_io_out ? io_r_559_b : _GEN_648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_650 = 10'h230 == r_count_0_io_out ? io_r_560_b : _GEN_649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_651 = 10'h231 == r_count_0_io_out ? io_r_561_b : _GEN_650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_652 = 10'h232 == r_count_0_io_out ? io_r_562_b : _GEN_651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_653 = 10'h233 == r_count_0_io_out ? io_r_563_b : _GEN_652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_654 = 10'h234 == r_count_0_io_out ? io_r_564_b : _GEN_653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_655 = 10'h235 == r_count_0_io_out ? io_r_565_b : _GEN_654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_656 = 10'h236 == r_count_0_io_out ? io_r_566_b : _GEN_655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_657 = 10'h237 == r_count_0_io_out ? io_r_567_b : _GEN_656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_658 = 10'h238 == r_count_0_io_out ? io_r_568_b : _GEN_657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_659 = 10'h239 == r_count_0_io_out ? io_r_569_b : _GEN_658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_660 = 10'h23a == r_count_0_io_out ? io_r_570_b : _GEN_659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_661 = 10'h23b == r_count_0_io_out ? io_r_571_b : _GEN_660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_662 = 10'h23c == r_count_0_io_out ? io_r_572_b : _GEN_661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_663 = 10'h23d == r_count_0_io_out ? io_r_573_b : _GEN_662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_664 = 10'h23e == r_count_0_io_out ? io_r_574_b : _GEN_663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_665 = 10'h23f == r_count_0_io_out ? io_r_575_b : _GEN_664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_666 = 10'h240 == r_count_0_io_out ? io_r_576_b : _GEN_665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_667 = 10'h241 == r_count_0_io_out ? io_r_577_b : _GEN_666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_668 = 10'h242 == r_count_0_io_out ? io_r_578_b : _GEN_667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_669 = 10'h243 == r_count_0_io_out ? io_r_579_b : _GEN_668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_670 = 10'h244 == r_count_0_io_out ? io_r_580_b : _GEN_669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_671 = 10'h245 == r_count_0_io_out ? io_r_581_b : _GEN_670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_672 = 10'h246 == r_count_0_io_out ? io_r_582_b : _GEN_671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_673 = 10'h247 == r_count_0_io_out ? io_r_583_b : _GEN_672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_674 = 10'h248 == r_count_0_io_out ? io_r_584_b : _GEN_673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_675 = 10'h249 == r_count_0_io_out ? io_r_585_b : _GEN_674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_676 = 10'h24a == r_count_0_io_out ? io_r_586_b : _GEN_675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_677 = 10'h24b == r_count_0_io_out ? io_r_587_b : _GEN_676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_678 = 10'h24c == r_count_0_io_out ? io_r_588_b : _GEN_677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_679 = 10'h24d == r_count_0_io_out ? io_r_589_b : _GEN_678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_680 = 10'h24e == r_count_0_io_out ? io_r_590_b : _GEN_679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_681 = 10'h24f == r_count_0_io_out ? io_r_591_b : _GEN_680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_682 = 10'h250 == r_count_0_io_out ? io_r_592_b : _GEN_681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_683 = 10'h251 == r_count_0_io_out ? io_r_593_b : _GEN_682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_684 = 10'h252 == r_count_0_io_out ? io_r_594_b : _GEN_683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_685 = 10'h253 == r_count_0_io_out ? io_r_595_b : _GEN_684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_686 = 10'h254 == r_count_0_io_out ? io_r_596_b : _GEN_685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_687 = 10'h255 == r_count_0_io_out ? io_r_597_b : _GEN_686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_688 = 10'h256 == r_count_0_io_out ? io_r_598_b : _GEN_687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_689 = 10'h257 == r_count_0_io_out ? io_r_599_b : _GEN_688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_690 = 10'h258 == r_count_0_io_out ? io_r_600_b : _GEN_689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_691 = 10'h259 == r_count_0_io_out ? io_r_601_b : _GEN_690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_692 = 10'h25a == r_count_0_io_out ? io_r_602_b : _GEN_691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_693 = 10'h25b == r_count_0_io_out ? io_r_603_b : _GEN_692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_694 = 10'h25c == r_count_0_io_out ? io_r_604_b : _GEN_693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_695 = 10'h25d == r_count_0_io_out ? io_r_605_b : _GEN_694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_696 = 10'h25e == r_count_0_io_out ? io_r_606_b : _GEN_695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_697 = 10'h25f == r_count_0_io_out ? io_r_607_b : _GEN_696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_698 = 10'h260 == r_count_0_io_out ? io_r_608_b : _GEN_697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_699 = 10'h261 == r_count_0_io_out ? io_r_609_b : _GEN_698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_700 = 10'h262 == r_count_0_io_out ? io_r_610_b : _GEN_699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_701 = 10'h263 == r_count_0_io_out ? io_r_611_b : _GEN_700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_702 = 10'h264 == r_count_0_io_out ? io_r_612_b : _GEN_701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_703 = 10'h265 == r_count_0_io_out ? io_r_613_b : _GEN_702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_704 = 10'h266 == r_count_0_io_out ? io_r_614_b : _GEN_703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_705 = 10'h267 == r_count_0_io_out ? io_r_615_b : _GEN_704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_706 = 10'h268 == r_count_0_io_out ? io_r_616_b : _GEN_705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_707 = 10'h269 == r_count_0_io_out ? io_r_617_b : _GEN_706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_708 = 10'h26a == r_count_0_io_out ? io_r_618_b : _GEN_707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_709 = 10'h26b == r_count_0_io_out ? io_r_619_b : _GEN_708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_710 = 10'h26c == r_count_0_io_out ? io_r_620_b : _GEN_709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_711 = 10'h26d == r_count_0_io_out ? io_r_621_b : _GEN_710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_712 = 10'h26e == r_count_0_io_out ? io_r_622_b : _GEN_711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_713 = 10'h26f == r_count_0_io_out ? io_r_623_b : _GEN_712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_714 = 10'h270 == r_count_0_io_out ? io_r_624_b : _GEN_713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_715 = 10'h271 == r_count_0_io_out ? io_r_625_b : _GEN_714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_716 = 10'h272 == r_count_0_io_out ? io_r_626_b : _GEN_715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_717 = 10'h273 == r_count_0_io_out ? io_r_627_b : _GEN_716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_718 = 10'h274 == r_count_0_io_out ? io_r_628_b : _GEN_717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_719 = 10'h275 == r_count_0_io_out ? io_r_629_b : _GEN_718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_720 = 10'h276 == r_count_0_io_out ? io_r_630_b : _GEN_719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_721 = 10'h277 == r_count_0_io_out ? io_r_631_b : _GEN_720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_722 = 10'h278 == r_count_0_io_out ? io_r_632_b : _GEN_721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_723 = 10'h279 == r_count_0_io_out ? io_r_633_b : _GEN_722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_724 = 10'h27a == r_count_0_io_out ? io_r_634_b : _GEN_723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_725 = 10'h27b == r_count_0_io_out ? io_r_635_b : _GEN_724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_726 = 10'h27c == r_count_0_io_out ? io_r_636_b : _GEN_725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_727 = 10'h27d == r_count_0_io_out ? io_r_637_b : _GEN_726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_728 = 10'h27e == r_count_0_io_out ? io_r_638_b : _GEN_727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_729 = 10'h27f == r_count_0_io_out ? io_r_639_b : _GEN_728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_730 = 10'h280 == r_count_0_io_out ? io_r_640_b : _GEN_729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_731 = 10'h281 == r_count_0_io_out ? io_r_641_b : _GEN_730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_732 = 10'h282 == r_count_0_io_out ? io_r_642_b : _GEN_731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_733 = 10'h283 == r_count_0_io_out ? io_r_643_b : _GEN_732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_734 = 10'h284 == r_count_0_io_out ? io_r_644_b : _GEN_733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_735 = 10'h285 == r_count_0_io_out ? io_r_645_b : _GEN_734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_736 = 10'h286 == r_count_0_io_out ? io_r_646_b : _GEN_735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_737 = 10'h287 == r_count_0_io_out ? io_r_647_b : _GEN_736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_738 = 10'h288 == r_count_0_io_out ? io_r_648_b : _GEN_737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_739 = 10'h289 == r_count_0_io_out ? io_r_649_b : _GEN_738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_740 = 10'h28a == r_count_0_io_out ? io_r_650_b : _GEN_739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_741 = 10'h28b == r_count_0_io_out ? io_r_651_b : _GEN_740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_742 = 10'h28c == r_count_0_io_out ? io_r_652_b : _GEN_741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_743 = 10'h28d == r_count_0_io_out ? io_r_653_b : _GEN_742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_744 = 10'h28e == r_count_0_io_out ? io_r_654_b : _GEN_743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_745 = 10'h28f == r_count_0_io_out ? io_r_655_b : _GEN_744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_746 = 10'h290 == r_count_0_io_out ? io_r_656_b : _GEN_745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_747 = 10'h291 == r_count_0_io_out ? io_r_657_b : _GEN_746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_748 = 10'h292 == r_count_0_io_out ? io_r_658_b : _GEN_747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_749 = 10'h293 == r_count_0_io_out ? io_r_659_b : _GEN_748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_750 = 10'h294 == r_count_0_io_out ? io_r_660_b : _GEN_749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_751 = 10'h295 == r_count_0_io_out ? io_r_661_b : _GEN_750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_752 = 10'h296 == r_count_0_io_out ? io_r_662_b : _GEN_751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_753 = 10'h297 == r_count_0_io_out ? io_r_663_b : _GEN_752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_754 = 10'h298 == r_count_0_io_out ? io_r_664_b : _GEN_753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_755 = 10'h299 == r_count_0_io_out ? io_r_665_b : _GEN_754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_756 = 10'h29a == r_count_0_io_out ? io_r_666_b : _GEN_755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_757 = 10'h29b == r_count_0_io_out ? io_r_667_b : _GEN_756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_758 = 10'h29c == r_count_0_io_out ? io_r_668_b : _GEN_757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_759 = 10'h29d == r_count_0_io_out ? io_r_669_b : _GEN_758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_760 = 10'h29e == r_count_0_io_out ? io_r_670_b : _GEN_759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_761 = 10'h29f == r_count_0_io_out ? io_r_671_b : _GEN_760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_762 = 10'h2a0 == r_count_0_io_out ? io_r_672_b : _GEN_761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_763 = 10'h2a1 == r_count_0_io_out ? io_r_673_b : _GEN_762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_764 = 10'h2a2 == r_count_0_io_out ? io_r_674_b : _GEN_763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_765 = 10'h2a3 == r_count_0_io_out ? io_r_675_b : _GEN_764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_766 = 10'h2a4 == r_count_0_io_out ? io_r_676_b : _GEN_765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_767 = 10'h2a5 == r_count_0_io_out ? io_r_677_b : _GEN_766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_768 = 10'h2a6 == r_count_0_io_out ? io_r_678_b : _GEN_767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_769 = 10'h2a7 == r_count_0_io_out ? io_r_679_b : _GEN_768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_770 = 10'h2a8 == r_count_0_io_out ? io_r_680_b : _GEN_769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_771 = 10'h2a9 == r_count_0_io_out ? io_r_681_b : _GEN_770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_772 = 10'h2aa == r_count_0_io_out ? io_r_682_b : _GEN_771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_773 = 10'h2ab == r_count_0_io_out ? io_r_683_b : _GEN_772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_774 = 10'h2ac == r_count_0_io_out ? io_r_684_b : _GEN_773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_775 = 10'h2ad == r_count_0_io_out ? io_r_685_b : _GEN_774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_776 = 10'h2ae == r_count_0_io_out ? io_r_686_b : _GEN_775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_777 = 10'h2af == r_count_0_io_out ? io_r_687_b : _GEN_776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_778 = 10'h2b0 == r_count_0_io_out ? io_r_688_b : _GEN_777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_779 = 10'h2b1 == r_count_0_io_out ? io_r_689_b : _GEN_778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_780 = 10'h2b2 == r_count_0_io_out ? io_r_690_b : _GEN_779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_781 = 10'h2b3 == r_count_0_io_out ? io_r_691_b : _GEN_780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_782 = 10'h2b4 == r_count_0_io_out ? io_r_692_b : _GEN_781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_783 = 10'h2b5 == r_count_0_io_out ? io_r_693_b : _GEN_782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_784 = 10'h2b6 == r_count_0_io_out ? io_r_694_b : _GEN_783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_785 = 10'h2b7 == r_count_0_io_out ? io_r_695_b : _GEN_784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_786 = 10'h2b8 == r_count_0_io_out ? io_r_696_b : _GEN_785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_787 = 10'h2b9 == r_count_0_io_out ? io_r_697_b : _GEN_786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_788 = 10'h2ba == r_count_0_io_out ? io_r_698_b : _GEN_787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_789 = 10'h2bb == r_count_0_io_out ? io_r_699_b : _GEN_788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_790 = 10'h2bc == r_count_0_io_out ? io_r_700_b : _GEN_789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_791 = 10'h2bd == r_count_0_io_out ? io_r_701_b : _GEN_790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_792 = 10'h2be == r_count_0_io_out ? io_r_702_b : _GEN_791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_793 = 10'h2bf == r_count_0_io_out ? io_r_703_b : _GEN_792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_794 = 10'h2c0 == r_count_0_io_out ? io_r_704_b : _GEN_793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_795 = 10'h2c1 == r_count_0_io_out ? io_r_705_b : _GEN_794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_796 = 10'h2c2 == r_count_0_io_out ? io_r_706_b : _GEN_795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_797 = 10'h2c3 == r_count_0_io_out ? io_r_707_b : _GEN_796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_798 = 10'h2c4 == r_count_0_io_out ? io_r_708_b : _GEN_797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_799 = 10'h2c5 == r_count_0_io_out ? io_r_709_b : _GEN_798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_800 = 10'h2c6 == r_count_0_io_out ? io_r_710_b : _GEN_799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_801 = 10'h2c7 == r_count_0_io_out ? io_r_711_b : _GEN_800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_802 = 10'h2c8 == r_count_0_io_out ? io_r_712_b : _GEN_801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_803 = 10'h2c9 == r_count_0_io_out ? io_r_713_b : _GEN_802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_804 = 10'h2ca == r_count_0_io_out ? io_r_714_b : _GEN_803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_805 = 10'h2cb == r_count_0_io_out ? io_r_715_b : _GEN_804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_806 = 10'h2cc == r_count_0_io_out ? io_r_716_b : _GEN_805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_807 = 10'h2cd == r_count_0_io_out ? io_r_717_b : _GEN_806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_808 = 10'h2ce == r_count_0_io_out ? io_r_718_b : _GEN_807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_809 = 10'h2cf == r_count_0_io_out ? io_r_719_b : _GEN_808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_810 = 10'h2d0 == r_count_0_io_out ? io_r_720_b : _GEN_809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_811 = 10'h2d1 == r_count_0_io_out ? io_r_721_b : _GEN_810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_812 = 10'h2d2 == r_count_0_io_out ? io_r_722_b : _GEN_811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_813 = 10'h2d3 == r_count_0_io_out ? io_r_723_b : _GEN_812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_814 = 10'h2d4 == r_count_0_io_out ? io_r_724_b : _GEN_813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_815 = 10'h2d5 == r_count_0_io_out ? io_r_725_b : _GEN_814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_816 = 10'h2d6 == r_count_0_io_out ? io_r_726_b : _GEN_815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_817 = 10'h2d7 == r_count_0_io_out ? io_r_727_b : _GEN_816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_818 = 10'h2d8 == r_count_0_io_out ? io_r_728_b : _GEN_817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_819 = 10'h2d9 == r_count_0_io_out ? io_r_729_b : _GEN_818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_820 = 10'h2da == r_count_0_io_out ? io_r_730_b : _GEN_819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_821 = 10'h2db == r_count_0_io_out ? io_r_731_b : _GEN_820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_822 = 10'h2dc == r_count_0_io_out ? io_r_732_b : _GEN_821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_823 = 10'h2dd == r_count_0_io_out ? io_r_733_b : _GEN_822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_824 = 10'h2de == r_count_0_io_out ? io_r_734_b : _GEN_823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_825 = 10'h2df == r_count_0_io_out ? io_r_735_b : _GEN_824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_826 = 10'h2e0 == r_count_0_io_out ? io_r_736_b : _GEN_825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_827 = 10'h2e1 == r_count_0_io_out ? io_r_737_b : _GEN_826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_828 = 10'h2e2 == r_count_0_io_out ? io_r_738_b : _GEN_827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_829 = 10'h2e3 == r_count_0_io_out ? io_r_739_b : _GEN_828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_830 = 10'h2e4 == r_count_0_io_out ? io_r_740_b : _GEN_829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_831 = 10'h2e5 == r_count_0_io_out ? io_r_741_b : _GEN_830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_832 = 10'h2e6 == r_count_0_io_out ? io_r_742_b : _GEN_831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_833 = 10'h2e7 == r_count_0_io_out ? io_r_743_b : _GEN_832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_834 = 10'h2e8 == r_count_0_io_out ? io_r_744_b : _GEN_833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_835 = 10'h2e9 == r_count_0_io_out ? io_r_745_b : _GEN_834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_836 = 10'h2ea == r_count_0_io_out ? io_r_746_b : _GEN_835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_837 = 10'h2eb == r_count_0_io_out ? io_r_747_b : _GEN_836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_838 = 10'h2ec == r_count_0_io_out ? io_r_748_b : _GEN_837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_841 = 10'h1 == r_count_1_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_842 = 10'h2 == r_count_1_io_out ? io_r_2_b : _GEN_841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_843 = 10'h3 == r_count_1_io_out ? io_r_3_b : _GEN_842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_844 = 10'h4 == r_count_1_io_out ? io_r_4_b : _GEN_843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_845 = 10'h5 == r_count_1_io_out ? io_r_5_b : _GEN_844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_846 = 10'h6 == r_count_1_io_out ? io_r_6_b : _GEN_845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_847 = 10'h7 == r_count_1_io_out ? io_r_7_b : _GEN_846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_848 = 10'h8 == r_count_1_io_out ? io_r_8_b : _GEN_847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_849 = 10'h9 == r_count_1_io_out ? io_r_9_b : _GEN_848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_850 = 10'ha == r_count_1_io_out ? io_r_10_b : _GEN_849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_851 = 10'hb == r_count_1_io_out ? io_r_11_b : _GEN_850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_852 = 10'hc == r_count_1_io_out ? io_r_12_b : _GEN_851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_853 = 10'hd == r_count_1_io_out ? io_r_13_b : _GEN_852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_854 = 10'he == r_count_1_io_out ? io_r_14_b : _GEN_853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_855 = 10'hf == r_count_1_io_out ? io_r_15_b : _GEN_854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_856 = 10'h10 == r_count_1_io_out ? io_r_16_b : _GEN_855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_857 = 10'h11 == r_count_1_io_out ? io_r_17_b : _GEN_856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_858 = 10'h12 == r_count_1_io_out ? io_r_18_b : _GEN_857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_859 = 10'h13 == r_count_1_io_out ? io_r_19_b : _GEN_858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_860 = 10'h14 == r_count_1_io_out ? io_r_20_b : _GEN_859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_861 = 10'h15 == r_count_1_io_out ? io_r_21_b : _GEN_860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_862 = 10'h16 == r_count_1_io_out ? io_r_22_b : _GEN_861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_863 = 10'h17 == r_count_1_io_out ? io_r_23_b : _GEN_862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_864 = 10'h18 == r_count_1_io_out ? io_r_24_b : _GEN_863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_865 = 10'h19 == r_count_1_io_out ? io_r_25_b : _GEN_864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_866 = 10'h1a == r_count_1_io_out ? io_r_26_b : _GEN_865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_867 = 10'h1b == r_count_1_io_out ? io_r_27_b : _GEN_866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_868 = 10'h1c == r_count_1_io_out ? io_r_28_b : _GEN_867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_869 = 10'h1d == r_count_1_io_out ? io_r_29_b : _GEN_868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_870 = 10'h1e == r_count_1_io_out ? io_r_30_b : _GEN_869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_871 = 10'h1f == r_count_1_io_out ? io_r_31_b : _GEN_870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_872 = 10'h20 == r_count_1_io_out ? io_r_32_b : _GEN_871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_873 = 10'h21 == r_count_1_io_out ? io_r_33_b : _GEN_872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_874 = 10'h22 == r_count_1_io_out ? io_r_34_b : _GEN_873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_875 = 10'h23 == r_count_1_io_out ? io_r_35_b : _GEN_874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_876 = 10'h24 == r_count_1_io_out ? io_r_36_b : _GEN_875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_877 = 10'h25 == r_count_1_io_out ? io_r_37_b : _GEN_876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_878 = 10'h26 == r_count_1_io_out ? io_r_38_b : _GEN_877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_879 = 10'h27 == r_count_1_io_out ? io_r_39_b : _GEN_878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_880 = 10'h28 == r_count_1_io_out ? io_r_40_b : _GEN_879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_881 = 10'h29 == r_count_1_io_out ? io_r_41_b : _GEN_880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_882 = 10'h2a == r_count_1_io_out ? io_r_42_b : _GEN_881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_883 = 10'h2b == r_count_1_io_out ? io_r_43_b : _GEN_882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_884 = 10'h2c == r_count_1_io_out ? io_r_44_b : _GEN_883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_885 = 10'h2d == r_count_1_io_out ? io_r_45_b : _GEN_884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_886 = 10'h2e == r_count_1_io_out ? io_r_46_b : _GEN_885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_887 = 10'h2f == r_count_1_io_out ? io_r_47_b : _GEN_886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_888 = 10'h30 == r_count_1_io_out ? io_r_48_b : _GEN_887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_889 = 10'h31 == r_count_1_io_out ? io_r_49_b : _GEN_888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_890 = 10'h32 == r_count_1_io_out ? io_r_50_b : _GEN_889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_891 = 10'h33 == r_count_1_io_out ? io_r_51_b : _GEN_890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_892 = 10'h34 == r_count_1_io_out ? io_r_52_b : _GEN_891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_893 = 10'h35 == r_count_1_io_out ? io_r_53_b : _GEN_892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_894 = 10'h36 == r_count_1_io_out ? io_r_54_b : _GEN_893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_895 = 10'h37 == r_count_1_io_out ? io_r_55_b : _GEN_894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_896 = 10'h38 == r_count_1_io_out ? io_r_56_b : _GEN_895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_897 = 10'h39 == r_count_1_io_out ? io_r_57_b : _GEN_896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_898 = 10'h3a == r_count_1_io_out ? io_r_58_b : _GEN_897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_899 = 10'h3b == r_count_1_io_out ? io_r_59_b : _GEN_898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_900 = 10'h3c == r_count_1_io_out ? io_r_60_b : _GEN_899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_901 = 10'h3d == r_count_1_io_out ? io_r_61_b : _GEN_900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_902 = 10'h3e == r_count_1_io_out ? io_r_62_b : _GEN_901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_903 = 10'h3f == r_count_1_io_out ? io_r_63_b : _GEN_902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_904 = 10'h40 == r_count_1_io_out ? io_r_64_b : _GEN_903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_905 = 10'h41 == r_count_1_io_out ? io_r_65_b : _GEN_904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_906 = 10'h42 == r_count_1_io_out ? io_r_66_b : _GEN_905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_907 = 10'h43 == r_count_1_io_out ? io_r_67_b : _GEN_906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_908 = 10'h44 == r_count_1_io_out ? io_r_68_b : _GEN_907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_909 = 10'h45 == r_count_1_io_out ? io_r_69_b : _GEN_908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_910 = 10'h46 == r_count_1_io_out ? io_r_70_b : _GEN_909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_911 = 10'h47 == r_count_1_io_out ? io_r_71_b : _GEN_910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_912 = 10'h48 == r_count_1_io_out ? io_r_72_b : _GEN_911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_913 = 10'h49 == r_count_1_io_out ? io_r_73_b : _GEN_912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_914 = 10'h4a == r_count_1_io_out ? io_r_74_b : _GEN_913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_915 = 10'h4b == r_count_1_io_out ? io_r_75_b : _GEN_914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_916 = 10'h4c == r_count_1_io_out ? io_r_76_b : _GEN_915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_917 = 10'h4d == r_count_1_io_out ? io_r_77_b : _GEN_916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_918 = 10'h4e == r_count_1_io_out ? io_r_78_b : _GEN_917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_919 = 10'h4f == r_count_1_io_out ? io_r_79_b : _GEN_918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_920 = 10'h50 == r_count_1_io_out ? io_r_80_b : _GEN_919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_921 = 10'h51 == r_count_1_io_out ? io_r_81_b : _GEN_920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_922 = 10'h52 == r_count_1_io_out ? io_r_82_b : _GEN_921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_923 = 10'h53 == r_count_1_io_out ? io_r_83_b : _GEN_922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_924 = 10'h54 == r_count_1_io_out ? io_r_84_b : _GEN_923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_925 = 10'h55 == r_count_1_io_out ? io_r_85_b : _GEN_924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_926 = 10'h56 == r_count_1_io_out ? io_r_86_b : _GEN_925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_927 = 10'h57 == r_count_1_io_out ? io_r_87_b : _GEN_926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_928 = 10'h58 == r_count_1_io_out ? io_r_88_b : _GEN_927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_929 = 10'h59 == r_count_1_io_out ? io_r_89_b : _GEN_928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_930 = 10'h5a == r_count_1_io_out ? io_r_90_b : _GEN_929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_931 = 10'h5b == r_count_1_io_out ? io_r_91_b : _GEN_930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_932 = 10'h5c == r_count_1_io_out ? io_r_92_b : _GEN_931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_933 = 10'h5d == r_count_1_io_out ? io_r_93_b : _GEN_932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_934 = 10'h5e == r_count_1_io_out ? io_r_94_b : _GEN_933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_935 = 10'h5f == r_count_1_io_out ? io_r_95_b : _GEN_934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_936 = 10'h60 == r_count_1_io_out ? io_r_96_b : _GEN_935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_937 = 10'h61 == r_count_1_io_out ? io_r_97_b : _GEN_936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_938 = 10'h62 == r_count_1_io_out ? io_r_98_b : _GEN_937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_939 = 10'h63 == r_count_1_io_out ? io_r_99_b : _GEN_938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_940 = 10'h64 == r_count_1_io_out ? io_r_100_b : _GEN_939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_941 = 10'h65 == r_count_1_io_out ? io_r_101_b : _GEN_940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_942 = 10'h66 == r_count_1_io_out ? io_r_102_b : _GEN_941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_943 = 10'h67 == r_count_1_io_out ? io_r_103_b : _GEN_942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_944 = 10'h68 == r_count_1_io_out ? io_r_104_b : _GEN_943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_945 = 10'h69 == r_count_1_io_out ? io_r_105_b : _GEN_944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_946 = 10'h6a == r_count_1_io_out ? io_r_106_b : _GEN_945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_947 = 10'h6b == r_count_1_io_out ? io_r_107_b : _GEN_946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_948 = 10'h6c == r_count_1_io_out ? io_r_108_b : _GEN_947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_949 = 10'h6d == r_count_1_io_out ? io_r_109_b : _GEN_948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_950 = 10'h6e == r_count_1_io_out ? io_r_110_b : _GEN_949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_951 = 10'h6f == r_count_1_io_out ? io_r_111_b : _GEN_950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_952 = 10'h70 == r_count_1_io_out ? io_r_112_b : _GEN_951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_953 = 10'h71 == r_count_1_io_out ? io_r_113_b : _GEN_952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_954 = 10'h72 == r_count_1_io_out ? io_r_114_b : _GEN_953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_955 = 10'h73 == r_count_1_io_out ? io_r_115_b : _GEN_954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_956 = 10'h74 == r_count_1_io_out ? io_r_116_b : _GEN_955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_957 = 10'h75 == r_count_1_io_out ? io_r_117_b : _GEN_956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_958 = 10'h76 == r_count_1_io_out ? io_r_118_b : _GEN_957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_959 = 10'h77 == r_count_1_io_out ? io_r_119_b : _GEN_958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_960 = 10'h78 == r_count_1_io_out ? io_r_120_b : _GEN_959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_961 = 10'h79 == r_count_1_io_out ? io_r_121_b : _GEN_960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_962 = 10'h7a == r_count_1_io_out ? io_r_122_b : _GEN_961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_963 = 10'h7b == r_count_1_io_out ? io_r_123_b : _GEN_962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_964 = 10'h7c == r_count_1_io_out ? io_r_124_b : _GEN_963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_965 = 10'h7d == r_count_1_io_out ? io_r_125_b : _GEN_964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_966 = 10'h7e == r_count_1_io_out ? io_r_126_b : _GEN_965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_967 = 10'h7f == r_count_1_io_out ? io_r_127_b : _GEN_966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_968 = 10'h80 == r_count_1_io_out ? io_r_128_b : _GEN_967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_969 = 10'h81 == r_count_1_io_out ? io_r_129_b : _GEN_968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_970 = 10'h82 == r_count_1_io_out ? io_r_130_b : _GEN_969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_971 = 10'h83 == r_count_1_io_out ? io_r_131_b : _GEN_970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_972 = 10'h84 == r_count_1_io_out ? io_r_132_b : _GEN_971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_973 = 10'h85 == r_count_1_io_out ? io_r_133_b : _GEN_972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_974 = 10'h86 == r_count_1_io_out ? io_r_134_b : _GEN_973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_975 = 10'h87 == r_count_1_io_out ? io_r_135_b : _GEN_974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_976 = 10'h88 == r_count_1_io_out ? io_r_136_b : _GEN_975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_977 = 10'h89 == r_count_1_io_out ? io_r_137_b : _GEN_976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_978 = 10'h8a == r_count_1_io_out ? io_r_138_b : _GEN_977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_979 = 10'h8b == r_count_1_io_out ? io_r_139_b : _GEN_978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_980 = 10'h8c == r_count_1_io_out ? io_r_140_b : _GEN_979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_981 = 10'h8d == r_count_1_io_out ? io_r_141_b : _GEN_980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_982 = 10'h8e == r_count_1_io_out ? io_r_142_b : _GEN_981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_983 = 10'h8f == r_count_1_io_out ? io_r_143_b : _GEN_982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_984 = 10'h90 == r_count_1_io_out ? io_r_144_b : _GEN_983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_985 = 10'h91 == r_count_1_io_out ? io_r_145_b : _GEN_984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_986 = 10'h92 == r_count_1_io_out ? io_r_146_b : _GEN_985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_987 = 10'h93 == r_count_1_io_out ? io_r_147_b : _GEN_986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_988 = 10'h94 == r_count_1_io_out ? io_r_148_b : _GEN_987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_989 = 10'h95 == r_count_1_io_out ? io_r_149_b : _GEN_988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_990 = 10'h96 == r_count_1_io_out ? io_r_150_b : _GEN_989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_991 = 10'h97 == r_count_1_io_out ? io_r_151_b : _GEN_990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_992 = 10'h98 == r_count_1_io_out ? io_r_152_b : _GEN_991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_993 = 10'h99 == r_count_1_io_out ? io_r_153_b : _GEN_992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_994 = 10'h9a == r_count_1_io_out ? io_r_154_b : _GEN_993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_995 = 10'h9b == r_count_1_io_out ? io_r_155_b : _GEN_994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_996 = 10'h9c == r_count_1_io_out ? io_r_156_b : _GEN_995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_997 = 10'h9d == r_count_1_io_out ? io_r_157_b : _GEN_996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_998 = 10'h9e == r_count_1_io_out ? io_r_158_b : _GEN_997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_999 = 10'h9f == r_count_1_io_out ? io_r_159_b : _GEN_998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1000 = 10'ha0 == r_count_1_io_out ? io_r_160_b : _GEN_999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1001 = 10'ha1 == r_count_1_io_out ? io_r_161_b : _GEN_1000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1002 = 10'ha2 == r_count_1_io_out ? io_r_162_b : _GEN_1001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1003 = 10'ha3 == r_count_1_io_out ? io_r_163_b : _GEN_1002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1004 = 10'ha4 == r_count_1_io_out ? io_r_164_b : _GEN_1003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1005 = 10'ha5 == r_count_1_io_out ? io_r_165_b : _GEN_1004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1006 = 10'ha6 == r_count_1_io_out ? io_r_166_b : _GEN_1005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1007 = 10'ha7 == r_count_1_io_out ? io_r_167_b : _GEN_1006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1008 = 10'ha8 == r_count_1_io_out ? io_r_168_b : _GEN_1007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1009 = 10'ha9 == r_count_1_io_out ? io_r_169_b : _GEN_1008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1010 = 10'haa == r_count_1_io_out ? io_r_170_b : _GEN_1009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1011 = 10'hab == r_count_1_io_out ? io_r_171_b : _GEN_1010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1012 = 10'hac == r_count_1_io_out ? io_r_172_b : _GEN_1011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1013 = 10'had == r_count_1_io_out ? io_r_173_b : _GEN_1012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1014 = 10'hae == r_count_1_io_out ? io_r_174_b : _GEN_1013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1015 = 10'haf == r_count_1_io_out ? io_r_175_b : _GEN_1014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1016 = 10'hb0 == r_count_1_io_out ? io_r_176_b : _GEN_1015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1017 = 10'hb1 == r_count_1_io_out ? io_r_177_b : _GEN_1016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1018 = 10'hb2 == r_count_1_io_out ? io_r_178_b : _GEN_1017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1019 = 10'hb3 == r_count_1_io_out ? io_r_179_b : _GEN_1018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1020 = 10'hb4 == r_count_1_io_out ? io_r_180_b : _GEN_1019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1021 = 10'hb5 == r_count_1_io_out ? io_r_181_b : _GEN_1020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1022 = 10'hb6 == r_count_1_io_out ? io_r_182_b : _GEN_1021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1023 = 10'hb7 == r_count_1_io_out ? io_r_183_b : _GEN_1022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1024 = 10'hb8 == r_count_1_io_out ? io_r_184_b : _GEN_1023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1025 = 10'hb9 == r_count_1_io_out ? io_r_185_b : _GEN_1024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1026 = 10'hba == r_count_1_io_out ? io_r_186_b : _GEN_1025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1027 = 10'hbb == r_count_1_io_out ? io_r_187_b : _GEN_1026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1028 = 10'hbc == r_count_1_io_out ? io_r_188_b : _GEN_1027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1029 = 10'hbd == r_count_1_io_out ? io_r_189_b : _GEN_1028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1030 = 10'hbe == r_count_1_io_out ? io_r_190_b : _GEN_1029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1031 = 10'hbf == r_count_1_io_out ? io_r_191_b : _GEN_1030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1032 = 10'hc0 == r_count_1_io_out ? io_r_192_b : _GEN_1031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1033 = 10'hc1 == r_count_1_io_out ? io_r_193_b : _GEN_1032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1034 = 10'hc2 == r_count_1_io_out ? io_r_194_b : _GEN_1033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1035 = 10'hc3 == r_count_1_io_out ? io_r_195_b : _GEN_1034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1036 = 10'hc4 == r_count_1_io_out ? io_r_196_b : _GEN_1035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1037 = 10'hc5 == r_count_1_io_out ? io_r_197_b : _GEN_1036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1038 = 10'hc6 == r_count_1_io_out ? io_r_198_b : _GEN_1037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1039 = 10'hc7 == r_count_1_io_out ? io_r_199_b : _GEN_1038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1040 = 10'hc8 == r_count_1_io_out ? io_r_200_b : _GEN_1039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1041 = 10'hc9 == r_count_1_io_out ? io_r_201_b : _GEN_1040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1042 = 10'hca == r_count_1_io_out ? io_r_202_b : _GEN_1041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1043 = 10'hcb == r_count_1_io_out ? io_r_203_b : _GEN_1042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1044 = 10'hcc == r_count_1_io_out ? io_r_204_b : _GEN_1043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1045 = 10'hcd == r_count_1_io_out ? io_r_205_b : _GEN_1044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1046 = 10'hce == r_count_1_io_out ? io_r_206_b : _GEN_1045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1047 = 10'hcf == r_count_1_io_out ? io_r_207_b : _GEN_1046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1048 = 10'hd0 == r_count_1_io_out ? io_r_208_b : _GEN_1047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1049 = 10'hd1 == r_count_1_io_out ? io_r_209_b : _GEN_1048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1050 = 10'hd2 == r_count_1_io_out ? io_r_210_b : _GEN_1049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1051 = 10'hd3 == r_count_1_io_out ? io_r_211_b : _GEN_1050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1052 = 10'hd4 == r_count_1_io_out ? io_r_212_b : _GEN_1051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1053 = 10'hd5 == r_count_1_io_out ? io_r_213_b : _GEN_1052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1054 = 10'hd6 == r_count_1_io_out ? io_r_214_b : _GEN_1053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1055 = 10'hd7 == r_count_1_io_out ? io_r_215_b : _GEN_1054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1056 = 10'hd8 == r_count_1_io_out ? io_r_216_b : _GEN_1055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1057 = 10'hd9 == r_count_1_io_out ? io_r_217_b : _GEN_1056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1058 = 10'hda == r_count_1_io_out ? io_r_218_b : _GEN_1057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1059 = 10'hdb == r_count_1_io_out ? io_r_219_b : _GEN_1058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1060 = 10'hdc == r_count_1_io_out ? io_r_220_b : _GEN_1059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1061 = 10'hdd == r_count_1_io_out ? io_r_221_b : _GEN_1060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1062 = 10'hde == r_count_1_io_out ? io_r_222_b : _GEN_1061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1063 = 10'hdf == r_count_1_io_out ? io_r_223_b : _GEN_1062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1064 = 10'he0 == r_count_1_io_out ? io_r_224_b : _GEN_1063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1065 = 10'he1 == r_count_1_io_out ? io_r_225_b : _GEN_1064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1066 = 10'he2 == r_count_1_io_out ? io_r_226_b : _GEN_1065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1067 = 10'he3 == r_count_1_io_out ? io_r_227_b : _GEN_1066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1068 = 10'he4 == r_count_1_io_out ? io_r_228_b : _GEN_1067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1069 = 10'he5 == r_count_1_io_out ? io_r_229_b : _GEN_1068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1070 = 10'he6 == r_count_1_io_out ? io_r_230_b : _GEN_1069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1071 = 10'he7 == r_count_1_io_out ? io_r_231_b : _GEN_1070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1072 = 10'he8 == r_count_1_io_out ? io_r_232_b : _GEN_1071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1073 = 10'he9 == r_count_1_io_out ? io_r_233_b : _GEN_1072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1074 = 10'hea == r_count_1_io_out ? io_r_234_b : _GEN_1073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1075 = 10'heb == r_count_1_io_out ? io_r_235_b : _GEN_1074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1076 = 10'hec == r_count_1_io_out ? io_r_236_b : _GEN_1075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1077 = 10'hed == r_count_1_io_out ? io_r_237_b : _GEN_1076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1078 = 10'hee == r_count_1_io_out ? io_r_238_b : _GEN_1077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1079 = 10'hef == r_count_1_io_out ? io_r_239_b : _GEN_1078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1080 = 10'hf0 == r_count_1_io_out ? io_r_240_b : _GEN_1079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1081 = 10'hf1 == r_count_1_io_out ? io_r_241_b : _GEN_1080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1082 = 10'hf2 == r_count_1_io_out ? io_r_242_b : _GEN_1081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1083 = 10'hf3 == r_count_1_io_out ? io_r_243_b : _GEN_1082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1084 = 10'hf4 == r_count_1_io_out ? io_r_244_b : _GEN_1083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1085 = 10'hf5 == r_count_1_io_out ? io_r_245_b : _GEN_1084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1086 = 10'hf6 == r_count_1_io_out ? io_r_246_b : _GEN_1085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1087 = 10'hf7 == r_count_1_io_out ? io_r_247_b : _GEN_1086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1088 = 10'hf8 == r_count_1_io_out ? io_r_248_b : _GEN_1087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1089 = 10'hf9 == r_count_1_io_out ? io_r_249_b : _GEN_1088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1090 = 10'hfa == r_count_1_io_out ? io_r_250_b : _GEN_1089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1091 = 10'hfb == r_count_1_io_out ? io_r_251_b : _GEN_1090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1092 = 10'hfc == r_count_1_io_out ? io_r_252_b : _GEN_1091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1093 = 10'hfd == r_count_1_io_out ? io_r_253_b : _GEN_1092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1094 = 10'hfe == r_count_1_io_out ? io_r_254_b : _GEN_1093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1095 = 10'hff == r_count_1_io_out ? io_r_255_b : _GEN_1094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1096 = 10'h100 == r_count_1_io_out ? io_r_256_b : _GEN_1095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1097 = 10'h101 == r_count_1_io_out ? io_r_257_b : _GEN_1096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1098 = 10'h102 == r_count_1_io_out ? io_r_258_b : _GEN_1097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1099 = 10'h103 == r_count_1_io_out ? io_r_259_b : _GEN_1098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1100 = 10'h104 == r_count_1_io_out ? io_r_260_b : _GEN_1099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1101 = 10'h105 == r_count_1_io_out ? io_r_261_b : _GEN_1100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1102 = 10'h106 == r_count_1_io_out ? io_r_262_b : _GEN_1101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1103 = 10'h107 == r_count_1_io_out ? io_r_263_b : _GEN_1102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1104 = 10'h108 == r_count_1_io_out ? io_r_264_b : _GEN_1103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1105 = 10'h109 == r_count_1_io_out ? io_r_265_b : _GEN_1104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1106 = 10'h10a == r_count_1_io_out ? io_r_266_b : _GEN_1105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1107 = 10'h10b == r_count_1_io_out ? io_r_267_b : _GEN_1106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1108 = 10'h10c == r_count_1_io_out ? io_r_268_b : _GEN_1107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1109 = 10'h10d == r_count_1_io_out ? io_r_269_b : _GEN_1108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1110 = 10'h10e == r_count_1_io_out ? io_r_270_b : _GEN_1109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1111 = 10'h10f == r_count_1_io_out ? io_r_271_b : _GEN_1110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1112 = 10'h110 == r_count_1_io_out ? io_r_272_b : _GEN_1111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1113 = 10'h111 == r_count_1_io_out ? io_r_273_b : _GEN_1112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1114 = 10'h112 == r_count_1_io_out ? io_r_274_b : _GEN_1113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1115 = 10'h113 == r_count_1_io_out ? io_r_275_b : _GEN_1114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1116 = 10'h114 == r_count_1_io_out ? io_r_276_b : _GEN_1115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1117 = 10'h115 == r_count_1_io_out ? io_r_277_b : _GEN_1116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1118 = 10'h116 == r_count_1_io_out ? io_r_278_b : _GEN_1117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1119 = 10'h117 == r_count_1_io_out ? io_r_279_b : _GEN_1118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1120 = 10'h118 == r_count_1_io_out ? io_r_280_b : _GEN_1119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1121 = 10'h119 == r_count_1_io_out ? io_r_281_b : _GEN_1120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1122 = 10'h11a == r_count_1_io_out ? io_r_282_b : _GEN_1121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1123 = 10'h11b == r_count_1_io_out ? io_r_283_b : _GEN_1122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1124 = 10'h11c == r_count_1_io_out ? io_r_284_b : _GEN_1123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1125 = 10'h11d == r_count_1_io_out ? io_r_285_b : _GEN_1124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1126 = 10'h11e == r_count_1_io_out ? io_r_286_b : _GEN_1125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1127 = 10'h11f == r_count_1_io_out ? io_r_287_b : _GEN_1126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1128 = 10'h120 == r_count_1_io_out ? io_r_288_b : _GEN_1127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1129 = 10'h121 == r_count_1_io_out ? io_r_289_b : _GEN_1128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1130 = 10'h122 == r_count_1_io_out ? io_r_290_b : _GEN_1129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1131 = 10'h123 == r_count_1_io_out ? io_r_291_b : _GEN_1130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1132 = 10'h124 == r_count_1_io_out ? io_r_292_b : _GEN_1131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1133 = 10'h125 == r_count_1_io_out ? io_r_293_b : _GEN_1132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1134 = 10'h126 == r_count_1_io_out ? io_r_294_b : _GEN_1133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1135 = 10'h127 == r_count_1_io_out ? io_r_295_b : _GEN_1134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1136 = 10'h128 == r_count_1_io_out ? io_r_296_b : _GEN_1135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1137 = 10'h129 == r_count_1_io_out ? io_r_297_b : _GEN_1136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1138 = 10'h12a == r_count_1_io_out ? io_r_298_b : _GEN_1137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1139 = 10'h12b == r_count_1_io_out ? io_r_299_b : _GEN_1138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1140 = 10'h12c == r_count_1_io_out ? io_r_300_b : _GEN_1139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1141 = 10'h12d == r_count_1_io_out ? io_r_301_b : _GEN_1140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1142 = 10'h12e == r_count_1_io_out ? io_r_302_b : _GEN_1141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1143 = 10'h12f == r_count_1_io_out ? io_r_303_b : _GEN_1142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1144 = 10'h130 == r_count_1_io_out ? io_r_304_b : _GEN_1143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1145 = 10'h131 == r_count_1_io_out ? io_r_305_b : _GEN_1144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1146 = 10'h132 == r_count_1_io_out ? io_r_306_b : _GEN_1145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1147 = 10'h133 == r_count_1_io_out ? io_r_307_b : _GEN_1146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1148 = 10'h134 == r_count_1_io_out ? io_r_308_b : _GEN_1147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1149 = 10'h135 == r_count_1_io_out ? io_r_309_b : _GEN_1148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1150 = 10'h136 == r_count_1_io_out ? io_r_310_b : _GEN_1149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1151 = 10'h137 == r_count_1_io_out ? io_r_311_b : _GEN_1150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1152 = 10'h138 == r_count_1_io_out ? io_r_312_b : _GEN_1151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1153 = 10'h139 == r_count_1_io_out ? io_r_313_b : _GEN_1152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1154 = 10'h13a == r_count_1_io_out ? io_r_314_b : _GEN_1153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1155 = 10'h13b == r_count_1_io_out ? io_r_315_b : _GEN_1154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1156 = 10'h13c == r_count_1_io_out ? io_r_316_b : _GEN_1155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1157 = 10'h13d == r_count_1_io_out ? io_r_317_b : _GEN_1156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1158 = 10'h13e == r_count_1_io_out ? io_r_318_b : _GEN_1157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1159 = 10'h13f == r_count_1_io_out ? io_r_319_b : _GEN_1158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1160 = 10'h140 == r_count_1_io_out ? io_r_320_b : _GEN_1159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1161 = 10'h141 == r_count_1_io_out ? io_r_321_b : _GEN_1160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1162 = 10'h142 == r_count_1_io_out ? io_r_322_b : _GEN_1161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1163 = 10'h143 == r_count_1_io_out ? io_r_323_b : _GEN_1162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1164 = 10'h144 == r_count_1_io_out ? io_r_324_b : _GEN_1163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1165 = 10'h145 == r_count_1_io_out ? io_r_325_b : _GEN_1164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1166 = 10'h146 == r_count_1_io_out ? io_r_326_b : _GEN_1165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1167 = 10'h147 == r_count_1_io_out ? io_r_327_b : _GEN_1166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1168 = 10'h148 == r_count_1_io_out ? io_r_328_b : _GEN_1167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1169 = 10'h149 == r_count_1_io_out ? io_r_329_b : _GEN_1168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1170 = 10'h14a == r_count_1_io_out ? io_r_330_b : _GEN_1169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1171 = 10'h14b == r_count_1_io_out ? io_r_331_b : _GEN_1170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1172 = 10'h14c == r_count_1_io_out ? io_r_332_b : _GEN_1171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1173 = 10'h14d == r_count_1_io_out ? io_r_333_b : _GEN_1172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1174 = 10'h14e == r_count_1_io_out ? io_r_334_b : _GEN_1173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1175 = 10'h14f == r_count_1_io_out ? io_r_335_b : _GEN_1174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1176 = 10'h150 == r_count_1_io_out ? io_r_336_b : _GEN_1175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1177 = 10'h151 == r_count_1_io_out ? io_r_337_b : _GEN_1176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1178 = 10'h152 == r_count_1_io_out ? io_r_338_b : _GEN_1177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1179 = 10'h153 == r_count_1_io_out ? io_r_339_b : _GEN_1178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1180 = 10'h154 == r_count_1_io_out ? io_r_340_b : _GEN_1179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1181 = 10'h155 == r_count_1_io_out ? io_r_341_b : _GEN_1180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1182 = 10'h156 == r_count_1_io_out ? io_r_342_b : _GEN_1181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1183 = 10'h157 == r_count_1_io_out ? io_r_343_b : _GEN_1182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1184 = 10'h158 == r_count_1_io_out ? io_r_344_b : _GEN_1183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1185 = 10'h159 == r_count_1_io_out ? io_r_345_b : _GEN_1184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1186 = 10'h15a == r_count_1_io_out ? io_r_346_b : _GEN_1185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1187 = 10'h15b == r_count_1_io_out ? io_r_347_b : _GEN_1186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1188 = 10'h15c == r_count_1_io_out ? io_r_348_b : _GEN_1187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1189 = 10'h15d == r_count_1_io_out ? io_r_349_b : _GEN_1188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1190 = 10'h15e == r_count_1_io_out ? io_r_350_b : _GEN_1189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1191 = 10'h15f == r_count_1_io_out ? io_r_351_b : _GEN_1190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1192 = 10'h160 == r_count_1_io_out ? io_r_352_b : _GEN_1191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1193 = 10'h161 == r_count_1_io_out ? io_r_353_b : _GEN_1192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1194 = 10'h162 == r_count_1_io_out ? io_r_354_b : _GEN_1193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1195 = 10'h163 == r_count_1_io_out ? io_r_355_b : _GEN_1194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1196 = 10'h164 == r_count_1_io_out ? io_r_356_b : _GEN_1195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1197 = 10'h165 == r_count_1_io_out ? io_r_357_b : _GEN_1196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1198 = 10'h166 == r_count_1_io_out ? io_r_358_b : _GEN_1197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1199 = 10'h167 == r_count_1_io_out ? io_r_359_b : _GEN_1198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1200 = 10'h168 == r_count_1_io_out ? io_r_360_b : _GEN_1199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1201 = 10'h169 == r_count_1_io_out ? io_r_361_b : _GEN_1200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1202 = 10'h16a == r_count_1_io_out ? io_r_362_b : _GEN_1201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1203 = 10'h16b == r_count_1_io_out ? io_r_363_b : _GEN_1202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1204 = 10'h16c == r_count_1_io_out ? io_r_364_b : _GEN_1203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1205 = 10'h16d == r_count_1_io_out ? io_r_365_b : _GEN_1204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1206 = 10'h16e == r_count_1_io_out ? io_r_366_b : _GEN_1205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1207 = 10'h16f == r_count_1_io_out ? io_r_367_b : _GEN_1206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1208 = 10'h170 == r_count_1_io_out ? io_r_368_b : _GEN_1207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1209 = 10'h171 == r_count_1_io_out ? io_r_369_b : _GEN_1208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1210 = 10'h172 == r_count_1_io_out ? io_r_370_b : _GEN_1209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1211 = 10'h173 == r_count_1_io_out ? io_r_371_b : _GEN_1210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1212 = 10'h174 == r_count_1_io_out ? io_r_372_b : _GEN_1211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1213 = 10'h175 == r_count_1_io_out ? io_r_373_b : _GEN_1212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1214 = 10'h176 == r_count_1_io_out ? io_r_374_b : _GEN_1213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1215 = 10'h177 == r_count_1_io_out ? io_r_375_b : _GEN_1214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1216 = 10'h178 == r_count_1_io_out ? io_r_376_b : _GEN_1215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1217 = 10'h179 == r_count_1_io_out ? io_r_377_b : _GEN_1216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1218 = 10'h17a == r_count_1_io_out ? io_r_378_b : _GEN_1217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1219 = 10'h17b == r_count_1_io_out ? io_r_379_b : _GEN_1218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1220 = 10'h17c == r_count_1_io_out ? io_r_380_b : _GEN_1219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1221 = 10'h17d == r_count_1_io_out ? io_r_381_b : _GEN_1220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1222 = 10'h17e == r_count_1_io_out ? io_r_382_b : _GEN_1221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1223 = 10'h17f == r_count_1_io_out ? io_r_383_b : _GEN_1222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1224 = 10'h180 == r_count_1_io_out ? io_r_384_b : _GEN_1223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1225 = 10'h181 == r_count_1_io_out ? io_r_385_b : _GEN_1224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1226 = 10'h182 == r_count_1_io_out ? io_r_386_b : _GEN_1225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1227 = 10'h183 == r_count_1_io_out ? io_r_387_b : _GEN_1226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1228 = 10'h184 == r_count_1_io_out ? io_r_388_b : _GEN_1227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1229 = 10'h185 == r_count_1_io_out ? io_r_389_b : _GEN_1228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1230 = 10'h186 == r_count_1_io_out ? io_r_390_b : _GEN_1229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1231 = 10'h187 == r_count_1_io_out ? io_r_391_b : _GEN_1230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1232 = 10'h188 == r_count_1_io_out ? io_r_392_b : _GEN_1231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1233 = 10'h189 == r_count_1_io_out ? io_r_393_b : _GEN_1232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1234 = 10'h18a == r_count_1_io_out ? io_r_394_b : _GEN_1233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1235 = 10'h18b == r_count_1_io_out ? io_r_395_b : _GEN_1234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1236 = 10'h18c == r_count_1_io_out ? io_r_396_b : _GEN_1235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1237 = 10'h18d == r_count_1_io_out ? io_r_397_b : _GEN_1236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1238 = 10'h18e == r_count_1_io_out ? io_r_398_b : _GEN_1237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1239 = 10'h18f == r_count_1_io_out ? io_r_399_b : _GEN_1238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1240 = 10'h190 == r_count_1_io_out ? io_r_400_b : _GEN_1239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1241 = 10'h191 == r_count_1_io_out ? io_r_401_b : _GEN_1240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1242 = 10'h192 == r_count_1_io_out ? io_r_402_b : _GEN_1241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1243 = 10'h193 == r_count_1_io_out ? io_r_403_b : _GEN_1242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1244 = 10'h194 == r_count_1_io_out ? io_r_404_b : _GEN_1243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1245 = 10'h195 == r_count_1_io_out ? io_r_405_b : _GEN_1244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1246 = 10'h196 == r_count_1_io_out ? io_r_406_b : _GEN_1245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1247 = 10'h197 == r_count_1_io_out ? io_r_407_b : _GEN_1246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1248 = 10'h198 == r_count_1_io_out ? io_r_408_b : _GEN_1247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1249 = 10'h199 == r_count_1_io_out ? io_r_409_b : _GEN_1248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1250 = 10'h19a == r_count_1_io_out ? io_r_410_b : _GEN_1249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1251 = 10'h19b == r_count_1_io_out ? io_r_411_b : _GEN_1250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1252 = 10'h19c == r_count_1_io_out ? io_r_412_b : _GEN_1251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1253 = 10'h19d == r_count_1_io_out ? io_r_413_b : _GEN_1252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1254 = 10'h19e == r_count_1_io_out ? io_r_414_b : _GEN_1253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1255 = 10'h19f == r_count_1_io_out ? io_r_415_b : _GEN_1254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1256 = 10'h1a0 == r_count_1_io_out ? io_r_416_b : _GEN_1255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1257 = 10'h1a1 == r_count_1_io_out ? io_r_417_b : _GEN_1256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1258 = 10'h1a2 == r_count_1_io_out ? io_r_418_b : _GEN_1257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1259 = 10'h1a3 == r_count_1_io_out ? io_r_419_b : _GEN_1258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1260 = 10'h1a4 == r_count_1_io_out ? io_r_420_b : _GEN_1259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1261 = 10'h1a5 == r_count_1_io_out ? io_r_421_b : _GEN_1260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1262 = 10'h1a6 == r_count_1_io_out ? io_r_422_b : _GEN_1261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1263 = 10'h1a7 == r_count_1_io_out ? io_r_423_b : _GEN_1262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1264 = 10'h1a8 == r_count_1_io_out ? io_r_424_b : _GEN_1263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1265 = 10'h1a9 == r_count_1_io_out ? io_r_425_b : _GEN_1264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1266 = 10'h1aa == r_count_1_io_out ? io_r_426_b : _GEN_1265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1267 = 10'h1ab == r_count_1_io_out ? io_r_427_b : _GEN_1266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1268 = 10'h1ac == r_count_1_io_out ? io_r_428_b : _GEN_1267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1269 = 10'h1ad == r_count_1_io_out ? io_r_429_b : _GEN_1268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1270 = 10'h1ae == r_count_1_io_out ? io_r_430_b : _GEN_1269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1271 = 10'h1af == r_count_1_io_out ? io_r_431_b : _GEN_1270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1272 = 10'h1b0 == r_count_1_io_out ? io_r_432_b : _GEN_1271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1273 = 10'h1b1 == r_count_1_io_out ? io_r_433_b : _GEN_1272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1274 = 10'h1b2 == r_count_1_io_out ? io_r_434_b : _GEN_1273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1275 = 10'h1b3 == r_count_1_io_out ? io_r_435_b : _GEN_1274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1276 = 10'h1b4 == r_count_1_io_out ? io_r_436_b : _GEN_1275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1277 = 10'h1b5 == r_count_1_io_out ? io_r_437_b : _GEN_1276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1278 = 10'h1b6 == r_count_1_io_out ? io_r_438_b : _GEN_1277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1279 = 10'h1b7 == r_count_1_io_out ? io_r_439_b : _GEN_1278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1280 = 10'h1b8 == r_count_1_io_out ? io_r_440_b : _GEN_1279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1281 = 10'h1b9 == r_count_1_io_out ? io_r_441_b : _GEN_1280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1282 = 10'h1ba == r_count_1_io_out ? io_r_442_b : _GEN_1281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1283 = 10'h1bb == r_count_1_io_out ? io_r_443_b : _GEN_1282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1284 = 10'h1bc == r_count_1_io_out ? io_r_444_b : _GEN_1283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1285 = 10'h1bd == r_count_1_io_out ? io_r_445_b : _GEN_1284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1286 = 10'h1be == r_count_1_io_out ? io_r_446_b : _GEN_1285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1287 = 10'h1bf == r_count_1_io_out ? io_r_447_b : _GEN_1286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1288 = 10'h1c0 == r_count_1_io_out ? io_r_448_b : _GEN_1287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1289 = 10'h1c1 == r_count_1_io_out ? io_r_449_b : _GEN_1288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1290 = 10'h1c2 == r_count_1_io_out ? io_r_450_b : _GEN_1289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1291 = 10'h1c3 == r_count_1_io_out ? io_r_451_b : _GEN_1290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1292 = 10'h1c4 == r_count_1_io_out ? io_r_452_b : _GEN_1291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1293 = 10'h1c5 == r_count_1_io_out ? io_r_453_b : _GEN_1292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1294 = 10'h1c6 == r_count_1_io_out ? io_r_454_b : _GEN_1293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1295 = 10'h1c7 == r_count_1_io_out ? io_r_455_b : _GEN_1294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1296 = 10'h1c8 == r_count_1_io_out ? io_r_456_b : _GEN_1295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1297 = 10'h1c9 == r_count_1_io_out ? io_r_457_b : _GEN_1296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1298 = 10'h1ca == r_count_1_io_out ? io_r_458_b : _GEN_1297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1299 = 10'h1cb == r_count_1_io_out ? io_r_459_b : _GEN_1298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1300 = 10'h1cc == r_count_1_io_out ? io_r_460_b : _GEN_1299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1301 = 10'h1cd == r_count_1_io_out ? io_r_461_b : _GEN_1300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1302 = 10'h1ce == r_count_1_io_out ? io_r_462_b : _GEN_1301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1303 = 10'h1cf == r_count_1_io_out ? io_r_463_b : _GEN_1302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1304 = 10'h1d0 == r_count_1_io_out ? io_r_464_b : _GEN_1303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1305 = 10'h1d1 == r_count_1_io_out ? io_r_465_b : _GEN_1304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1306 = 10'h1d2 == r_count_1_io_out ? io_r_466_b : _GEN_1305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1307 = 10'h1d3 == r_count_1_io_out ? io_r_467_b : _GEN_1306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1308 = 10'h1d4 == r_count_1_io_out ? io_r_468_b : _GEN_1307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1309 = 10'h1d5 == r_count_1_io_out ? io_r_469_b : _GEN_1308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1310 = 10'h1d6 == r_count_1_io_out ? io_r_470_b : _GEN_1309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1311 = 10'h1d7 == r_count_1_io_out ? io_r_471_b : _GEN_1310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1312 = 10'h1d8 == r_count_1_io_out ? io_r_472_b : _GEN_1311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1313 = 10'h1d9 == r_count_1_io_out ? io_r_473_b : _GEN_1312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1314 = 10'h1da == r_count_1_io_out ? io_r_474_b : _GEN_1313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1315 = 10'h1db == r_count_1_io_out ? io_r_475_b : _GEN_1314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1316 = 10'h1dc == r_count_1_io_out ? io_r_476_b : _GEN_1315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1317 = 10'h1dd == r_count_1_io_out ? io_r_477_b : _GEN_1316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1318 = 10'h1de == r_count_1_io_out ? io_r_478_b : _GEN_1317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1319 = 10'h1df == r_count_1_io_out ? io_r_479_b : _GEN_1318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1320 = 10'h1e0 == r_count_1_io_out ? io_r_480_b : _GEN_1319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1321 = 10'h1e1 == r_count_1_io_out ? io_r_481_b : _GEN_1320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1322 = 10'h1e2 == r_count_1_io_out ? io_r_482_b : _GEN_1321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1323 = 10'h1e3 == r_count_1_io_out ? io_r_483_b : _GEN_1322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1324 = 10'h1e4 == r_count_1_io_out ? io_r_484_b : _GEN_1323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1325 = 10'h1e5 == r_count_1_io_out ? io_r_485_b : _GEN_1324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1326 = 10'h1e6 == r_count_1_io_out ? io_r_486_b : _GEN_1325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1327 = 10'h1e7 == r_count_1_io_out ? io_r_487_b : _GEN_1326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1328 = 10'h1e8 == r_count_1_io_out ? io_r_488_b : _GEN_1327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1329 = 10'h1e9 == r_count_1_io_out ? io_r_489_b : _GEN_1328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1330 = 10'h1ea == r_count_1_io_out ? io_r_490_b : _GEN_1329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1331 = 10'h1eb == r_count_1_io_out ? io_r_491_b : _GEN_1330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1332 = 10'h1ec == r_count_1_io_out ? io_r_492_b : _GEN_1331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1333 = 10'h1ed == r_count_1_io_out ? io_r_493_b : _GEN_1332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1334 = 10'h1ee == r_count_1_io_out ? io_r_494_b : _GEN_1333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1335 = 10'h1ef == r_count_1_io_out ? io_r_495_b : _GEN_1334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1336 = 10'h1f0 == r_count_1_io_out ? io_r_496_b : _GEN_1335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1337 = 10'h1f1 == r_count_1_io_out ? io_r_497_b : _GEN_1336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1338 = 10'h1f2 == r_count_1_io_out ? io_r_498_b : _GEN_1337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1339 = 10'h1f3 == r_count_1_io_out ? io_r_499_b : _GEN_1338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1340 = 10'h1f4 == r_count_1_io_out ? io_r_500_b : _GEN_1339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1341 = 10'h1f5 == r_count_1_io_out ? io_r_501_b : _GEN_1340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1342 = 10'h1f6 == r_count_1_io_out ? io_r_502_b : _GEN_1341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1343 = 10'h1f7 == r_count_1_io_out ? io_r_503_b : _GEN_1342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1344 = 10'h1f8 == r_count_1_io_out ? io_r_504_b : _GEN_1343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1345 = 10'h1f9 == r_count_1_io_out ? io_r_505_b : _GEN_1344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1346 = 10'h1fa == r_count_1_io_out ? io_r_506_b : _GEN_1345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1347 = 10'h1fb == r_count_1_io_out ? io_r_507_b : _GEN_1346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1348 = 10'h1fc == r_count_1_io_out ? io_r_508_b : _GEN_1347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1349 = 10'h1fd == r_count_1_io_out ? io_r_509_b : _GEN_1348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1350 = 10'h1fe == r_count_1_io_out ? io_r_510_b : _GEN_1349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1351 = 10'h1ff == r_count_1_io_out ? io_r_511_b : _GEN_1350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1352 = 10'h200 == r_count_1_io_out ? io_r_512_b : _GEN_1351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1353 = 10'h201 == r_count_1_io_out ? io_r_513_b : _GEN_1352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1354 = 10'h202 == r_count_1_io_out ? io_r_514_b : _GEN_1353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1355 = 10'h203 == r_count_1_io_out ? io_r_515_b : _GEN_1354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1356 = 10'h204 == r_count_1_io_out ? io_r_516_b : _GEN_1355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1357 = 10'h205 == r_count_1_io_out ? io_r_517_b : _GEN_1356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1358 = 10'h206 == r_count_1_io_out ? io_r_518_b : _GEN_1357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1359 = 10'h207 == r_count_1_io_out ? io_r_519_b : _GEN_1358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1360 = 10'h208 == r_count_1_io_out ? io_r_520_b : _GEN_1359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1361 = 10'h209 == r_count_1_io_out ? io_r_521_b : _GEN_1360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1362 = 10'h20a == r_count_1_io_out ? io_r_522_b : _GEN_1361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1363 = 10'h20b == r_count_1_io_out ? io_r_523_b : _GEN_1362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1364 = 10'h20c == r_count_1_io_out ? io_r_524_b : _GEN_1363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1365 = 10'h20d == r_count_1_io_out ? io_r_525_b : _GEN_1364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1366 = 10'h20e == r_count_1_io_out ? io_r_526_b : _GEN_1365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1367 = 10'h20f == r_count_1_io_out ? io_r_527_b : _GEN_1366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1368 = 10'h210 == r_count_1_io_out ? io_r_528_b : _GEN_1367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1369 = 10'h211 == r_count_1_io_out ? io_r_529_b : _GEN_1368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1370 = 10'h212 == r_count_1_io_out ? io_r_530_b : _GEN_1369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1371 = 10'h213 == r_count_1_io_out ? io_r_531_b : _GEN_1370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1372 = 10'h214 == r_count_1_io_out ? io_r_532_b : _GEN_1371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1373 = 10'h215 == r_count_1_io_out ? io_r_533_b : _GEN_1372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1374 = 10'h216 == r_count_1_io_out ? io_r_534_b : _GEN_1373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1375 = 10'h217 == r_count_1_io_out ? io_r_535_b : _GEN_1374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1376 = 10'h218 == r_count_1_io_out ? io_r_536_b : _GEN_1375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1377 = 10'h219 == r_count_1_io_out ? io_r_537_b : _GEN_1376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1378 = 10'h21a == r_count_1_io_out ? io_r_538_b : _GEN_1377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1379 = 10'h21b == r_count_1_io_out ? io_r_539_b : _GEN_1378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1380 = 10'h21c == r_count_1_io_out ? io_r_540_b : _GEN_1379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1381 = 10'h21d == r_count_1_io_out ? io_r_541_b : _GEN_1380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1382 = 10'h21e == r_count_1_io_out ? io_r_542_b : _GEN_1381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1383 = 10'h21f == r_count_1_io_out ? io_r_543_b : _GEN_1382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1384 = 10'h220 == r_count_1_io_out ? io_r_544_b : _GEN_1383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1385 = 10'h221 == r_count_1_io_out ? io_r_545_b : _GEN_1384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1386 = 10'h222 == r_count_1_io_out ? io_r_546_b : _GEN_1385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1387 = 10'h223 == r_count_1_io_out ? io_r_547_b : _GEN_1386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1388 = 10'h224 == r_count_1_io_out ? io_r_548_b : _GEN_1387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1389 = 10'h225 == r_count_1_io_out ? io_r_549_b : _GEN_1388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1390 = 10'h226 == r_count_1_io_out ? io_r_550_b : _GEN_1389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1391 = 10'h227 == r_count_1_io_out ? io_r_551_b : _GEN_1390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1392 = 10'h228 == r_count_1_io_out ? io_r_552_b : _GEN_1391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1393 = 10'h229 == r_count_1_io_out ? io_r_553_b : _GEN_1392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1394 = 10'h22a == r_count_1_io_out ? io_r_554_b : _GEN_1393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1395 = 10'h22b == r_count_1_io_out ? io_r_555_b : _GEN_1394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1396 = 10'h22c == r_count_1_io_out ? io_r_556_b : _GEN_1395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1397 = 10'h22d == r_count_1_io_out ? io_r_557_b : _GEN_1396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1398 = 10'h22e == r_count_1_io_out ? io_r_558_b : _GEN_1397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1399 = 10'h22f == r_count_1_io_out ? io_r_559_b : _GEN_1398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1400 = 10'h230 == r_count_1_io_out ? io_r_560_b : _GEN_1399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1401 = 10'h231 == r_count_1_io_out ? io_r_561_b : _GEN_1400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1402 = 10'h232 == r_count_1_io_out ? io_r_562_b : _GEN_1401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1403 = 10'h233 == r_count_1_io_out ? io_r_563_b : _GEN_1402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1404 = 10'h234 == r_count_1_io_out ? io_r_564_b : _GEN_1403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1405 = 10'h235 == r_count_1_io_out ? io_r_565_b : _GEN_1404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1406 = 10'h236 == r_count_1_io_out ? io_r_566_b : _GEN_1405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1407 = 10'h237 == r_count_1_io_out ? io_r_567_b : _GEN_1406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1408 = 10'h238 == r_count_1_io_out ? io_r_568_b : _GEN_1407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1409 = 10'h239 == r_count_1_io_out ? io_r_569_b : _GEN_1408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1410 = 10'h23a == r_count_1_io_out ? io_r_570_b : _GEN_1409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1411 = 10'h23b == r_count_1_io_out ? io_r_571_b : _GEN_1410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1412 = 10'h23c == r_count_1_io_out ? io_r_572_b : _GEN_1411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1413 = 10'h23d == r_count_1_io_out ? io_r_573_b : _GEN_1412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1414 = 10'h23e == r_count_1_io_out ? io_r_574_b : _GEN_1413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1415 = 10'h23f == r_count_1_io_out ? io_r_575_b : _GEN_1414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1416 = 10'h240 == r_count_1_io_out ? io_r_576_b : _GEN_1415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1417 = 10'h241 == r_count_1_io_out ? io_r_577_b : _GEN_1416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1418 = 10'h242 == r_count_1_io_out ? io_r_578_b : _GEN_1417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1419 = 10'h243 == r_count_1_io_out ? io_r_579_b : _GEN_1418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1420 = 10'h244 == r_count_1_io_out ? io_r_580_b : _GEN_1419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1421 = 10'h245 == r_count_1_io_out ? io_r_581_b : _GEN_1420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1422 = 10'h246 == r_count_1_io_out ? io_r_582_b : _GEN_1421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1423 = 10'h247 == r_count_1_io_out ? io_r_583_b : _GEN_1422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1424 = 10'h248 == r_count_1_io_out ? io_r_584_b : _GEN_1423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1425 = 10'h249 == r_count_1_io_out ? io_r_585_b : _GEN_1424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1426 = 10'h24a == r_count_1_io_out ? io_r_586_b : _GEN_1425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1427 = 10'h24b == r_count_1_io_out ? io_r_587_b : _GEN_1426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1428 = 10'h24c == r_count_1_io_out ? io_r_588_b : _GEN_1427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1429 = 10'h24d == r_count_1_io_out ? io_r_589_b : _GEN_1428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1430 = 10'h24e == r_count_1_io_out ? io_r_590_b : _GEN_1429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1431 = 10'h24f == r_count_1_io_out ? io_r_591_b : _GEN_1430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1432 = 10'h250 == r_count_1_io_out ? io_r_592_b : _GEN_1431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1433 = 10'h251 == r_count_1_io_out ? io_r_593_b : _GEN_1432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1434 = 10'h252 == r_count_1_io_out ? io_r_594_b : _GEN_1433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1435 = 10'h253 == r_count_1_io_out ? io_r_595_b : _GEN_1434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1436 = 10'h254 == r_count_1_io_out ? io_r_596_b : _GEN_1435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1437 = 10'h255 == r_count_1_io_out ? io_r_597_b : _GEN_1436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1438 = 10'h256 == r_count_1_io_out ? io_r_598_b : _GEN_1437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1439 = 10'h257 == r_count_1_io_out ? io_r_599_b : _GEN_1438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1440 = 10'h258 == r_count_1_io_out ? io_r_600_b : _GEN_1439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1441 = 10'h259 == r_count_1_io_out ? io_r_601_b : _GEN_1440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1442 = 10'h25a == r_count_1_io_out ? io_r_602_b : _GEN_1441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1443 = 10'h25b == r_count_1_io_out ? io_r_603_b : _GEN_1442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1444 = 10'h25c == r_count_1_io_out ? io_r_604_b : _GEN_1443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1445 = 10'h25d == r_count_1_io_out ? io_r_605_b : _GEN_1444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1446 = 10'h25e == r_count_1_io_out ? io_r_606_b : _GEN_1445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1447 = 10'h25f == r_count_1_io_out ? io_r_607_b : _GEN_1446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1448 = 10'h260 == r_count_1_io_out ? io_r_608_b : _GEN_1447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1449 = 10'h261 == r_count_1_io_out ? io_r_609_b : _GEN_1448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1450 = 10'h262 == r_count_1_io_out ? io_r_610_b : _GEN_1449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1451 = 10'h263 == r_count_1_io_out ? io_r_611_b : _GEN_1450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1452 = 10'h264 == r_count_1_io_out ? io_r_612_b : _GEN_1451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1453 = 10'h265 == r_count_1_io_out ? io_r_613_b : _GEN_1452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1454 = 10'h266 == r_count_1_io_out ? io_r_614_b : _GEN_1453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1455 = 10'h267 == r_count_1_io_out ? io_r_615_b : _GEN_1454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1456 = 10'h268 == r_count_1_io_out ? io_r_616_b : _GEN_1455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1457 = 10'h269 == r_count_1_io_out ? io_r_617_b : _GEN_1456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1458 = 10'h26a == r_count_1_io_out ? io_r_618_b : _GEN_1457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1459 = 10'h26b == r_count_1_io_out ? io_r_619_b : _GEN_1458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1460 = 10'h26c == r_count_1_io_out ? io_r_620_b : _GEN_1459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1461 = 10'h26d == r_count_1_io_out ? io_r_621_b : _GEN_1460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1462 = 10'h26e == r_count_1_io_out ? io_r_622_b : _GEN_1461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1463 = 10'h26f == r_count_1_io_out ? io_r_623_b : _GEN_1462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1464 = 10'h270 == r_count_1_io_out ? io_r_624_b : _GEN_1463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1465 = 10'h271 == r_count_1_io_out ? io_r_625_b : _GEN_1464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1466 = 10'h272 == r_count_1_io_out ? io_r_626_b : _GEN_1465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1467 = 10'h273 == r_count_1_io_out ? io_r_627_b : _GEN_1466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1468 = 10'h274 == r_count_1_io_out ? io_r_628_b : _GEN_1467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1469 = 10'h275 == r_count_1_io_out ? io_r_629_b : _GEN_1468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1470 = 10'h276 == r_count_1_io_out ? io_r_630_b : _GEN_1469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1471 = 10'h277 == r_count_1_io_out ? io_r_631_b : _GEN_1470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1472 = 10'h278 == r_count_1_io_out ? io_r_632_b : _GEN_1471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1473 = 10'h279 == r_count_1_io_out ? io_r_633_b : _GEN_1472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1474 = 10'h27a == r_count_1_io_out ? io_r_634_b : _GEN_1473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1475 = 10'h27b == r_count_1_io_out ? io_r_635_b : _GEN_1474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1476 = 10'h27c == r_count_1_io_out ? io_r_636_b : _GEN_1475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1477 = 10'h27d == r_count_1_io_out ? io_r_637_b : _GEN_1476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1478 = 10'h27e == r_count_1_io_out ? io_r_638_b : _GEN_1477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1479 = 10'h27f == r_count_1_io_out ? io_r_639_b : _GEN_1478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1480 = 10'h280 == r_count_1_io_out ? io_r_640_b : _GEN_1479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1481 = 10'h281 == r_count_1_io_out ? io_r_641_b : _GEN_1480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1482 = 10'h282 == r_count_1_io_out ? io_r_642_b : _GEN_1481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1483 = 10'h283 == r_count_1_io_out ? io_r_643_b : _GEN_1482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1484 = 10'h284 == r_count_1_io_out ? io_r_644_b : _GEN_1483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1485 = 10'h285 == r_count_1_io_out ? io_r_645_b : _GEN_1484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1486 = 10'h286 == r_count_1_io_out ? io_r_646_b : _GEN_1485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1487 = 10'h287 == r_count_1_io_out ? io_r_647_b : _GEN_1486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1488 = 10'h288 == r_count_1_io_out ? io_r_648_b : _GEN_1487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1489 = 10'h289 == r_count_1_io_out ? io_r_649_b : _GEN_1488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1490 = 10'h28a == r_count_1_io_out ? io_r_650_b : _GEN_1489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1491 = 10'h28b == r_count_1_io_out ? io_r_651_b : _GEN_1490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1492 = 10'h28c == r_count_1_io_out ? io_r_652_b : _GEN_1491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1493 = 10'h28d == r_count_1_io_out ? io_r_653_b : _GEN_1492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1494 = 10'h28e == r_count_1_io_out ? io_r_654_b : _GEN_1493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1495 = 10'h28f == r_count_1_io_out ? io_r_655_b : _GEN_1494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1496 = 10'h290 == r_count_1_io_out ? io_r_656_b : _GEN_1495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1497 = 10'h291 == r_count_1_io_out ? io_r_657_b : _GEN_1496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1498 = 10'h292 == r_count_1_io_out ? io_r_658_b : _GEN_1497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1499 = 10'h293 == r_count_1_io_out ? io_r_659_b : _GEN_1498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1500 = 10'h294 == r_count_1_io_out ? io_r_660_b : _GEN_1499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1501 = 10'h295 == r_count_1_io_out ? io_r_661_b : _GEN_1500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1502 = 10'h296 == r_count_1_io_out ? io_r_662_b : _GEN_1501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1503 = 10'h297 == r_count_1_io_out ? io_r_663_b : _GEN_1502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1504 = 10'h298 == r_count_1_io_out ? io_r_664_b : _GEN_1503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1505 = 10'h299 == r_count_1_io_out ? io_r_665_b : _GEN_1504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1506 = 10'h29a == r_count_1_io_out ? io_r_666_b : _GEN_1505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1507 = 10'h29b == r_count_1_io_out ? io_r_667_b : _GEN_1506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1508 = 10'h29c == r_count_1_io_out ? io_r_668_b : _GEN_1507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1509 = 10'h29d == r_count_1_io_out ? io_r_669_b : _GEN_1508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1510 = 10'h29e == r_count_1_io_out ? io_r_670_b : _GEN_1509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1511 = 10'h29f == r_count_1_io_out ? io_r_671_b : _GEN_1510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1512 = 10'h2a0 == r_count_1_io_out ? io_r_672_b : _GEN_1511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1513 = 10'h2a1 == r_count_1_io_out ? io_r_673_b : _GEN_1512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1514 = 10'h2a2 == r_count_1_io_out ? io_r_674_b : _GEN_1513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1515 = 10'h2a3 == r_count_1_io_out ? io_r_675_b : _GEN_1514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1516 = 10'h2a4 == r_count_1_io_out ? io_r_676_b : _GEN_1515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1517 = 10'h2a5 == r_count_1_io_out ? io_r_677_b : _GEN_1516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1518 = 10'h2a6 == r_count_1_io_out ? io_r_678_b : _GEN_1517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1519 = 10'h2a7 == r_count_1_io_out ? io_r_679_b : _GEN_1518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1520 = 10'h2a8 == r_count_1_io_out ? io_r_680_b : _GEN_1519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1521 = 10'h2a9 == r_count_1_io_out ? io_r_681_b : _GEN_1520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1522 = 10'h2aa == r_count_1_io_out ? io_r_682_b : _GEN_1521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1523 = 10'h2ab == r_count_1_io_out ? io_r_683_b : _GEN_1522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1524 = 10'h2ac == r_count_1_io_out ? io_r_684_b : _GEN_1523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1525 = 10'h2ad == r_count_1_io_out ? io_r_685_b : _GEN_1524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1526 = 10'h2ae == r_count_1_io_out ? io_r_686_b : _GEN_1525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1527 = 10'h2af == r_count_1_io_out ? io_r_687_b : _GEN_1526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1528 = 10'h2b0 == r_count_1_io_out ? io_r_688_b : _GEN_1527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1529 = 10'h2b1 == r_count_1_io_out ? io_r_689_b : _GEN_1528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1530 = 10'h2b2 == r_count_1_io_out ? io_r_690_b : _GEN_1529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1531 = 10'h2b3 == r_count_1_io_out ? io_r_691_b : _GEN_1530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1532 = 10'h2b4 == r_count_1_io_out ? io_r_692_b : _GEN_1531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1533 = 10'h2b5 == r_count_1_io_out ? io_r_693_b : _GEN_1532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1534 = 10'h2b6 == r_count_1_io_out ? io_r_694_b : _GEN_1533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1535 = 10'h2b7 == r_count_1_io_out ? io_r_695_b : _GEN_1534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1536 = 10'h2b8 == r_count_1_io_out ? io_r_696_b : _GEN_1535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1537 = 10'h2b9 == r_count_1_io_out ? io_r_697_b : _GEN_1536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1538 = 10'h2ba == r_count_1_io_out ? io_r_698_b : _GEN_1537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1539 = 10'h2bb == r_count_1_io_out ? io_r_699_b : _GEN_1538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1540 = 10'h2bc == r_count_1_io_out ? io_r_700_b : _GEN_1539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1541 = 10'h2bd == r_count_1_io_out ? io_r_701_b : _GEN_1540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1542 = 10'h2be == r_count_1_io_out ? io_r_702_b : _GEN_1541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1543 = 10'h2bf == r_count_1_io_out ? io_r_703_b : _GEN_1542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1544 = 10'h2c0 == r_count_1_io_out ? io_r_704_b : _GEN_1543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1545 = 10'h2c1 == r_count_1_io_out ? io_r_705_b : _GEN_1544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1546 = 10'h2c2 == r_count_1_io_out ? io_r_706_b : _GEN_1545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1547 = 10'h2c3 == r_count_1_io_out ? io_r_707_b : _GEN_1546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1548 = 10'h2c4 == r_count_1_io_out ? io_r_708_b : _GEN_1547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1549 = 10'h2c5 == r_count_1_io_out ? io_r_709_b : _GEN_1548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1550 = 10'h2c6 == r_count_1_io_out ? io_r_710_b : _GEN_1549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1551 = 10'h2c7 == r_count_1_io_out ? io_r_711_b : _GEN_1550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1552 = 10'h2c8 == r_count_1_io_out ? io_r_712_b : _GEN_1551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1553 = 10'h2c9 == r_count_1_io_out ? io_r_713_b : _GEN_1552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1554 = 10'h2ca == r_count_1_io_out ? io_r_714_b : _GEN_1553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1555 = 10'h2cb == r_count_1_io_out ? io_r_715_b : _GEN_1554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1556 = 10'h2cc == r_count_1_io_out ? io_r_716_b : _GEN_1555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1557 = 10'h2cd == r_count_1_io_out ? io_r_717_b : _GEN_1556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1558 = 10'h2ce == r_count_1_io_out ? io_r_718_b : _GEN_1557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1559 = 10'h2cf == r_count_1_io_out ? io_r_719_b : _GEN_1558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1560 = 10'h2d0 == r_count_1_io_out ? io_r_720_b : _GEN_1559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1561 = 10'h2d1 == r_count_1_io_out ? io_r_721_b : _GEN_1560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1562 = 10'h2d2 == r_count_1_io_out ? io_r_722_b : _GEN_1561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1563 = 10'h2d3 == r_count_1_io_out ? io_r_723_b : _GEN_1562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1564 = 10'h2d4 == r_count_1_io_out ? io_r_724_b : _GEN_1563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1565 = 10'h2d5 == r_count_1_io_out ? io_r_725_b : _GEN_1564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1566 = 10'h2d6 == r_count_1_io_out ? io_r_726_b : _GEN_1565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1567 = 10'h2d7 == r_count_1_io_out ? io_r_727_b : _GEN_1566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1568 = 10'h2d8 == r_count_1_io_out ? io_r_728_b : _GEN_1567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1569 = 10'h2d9 == r_count_1_io_out ? io_r_729_b : _GEN_1568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1570 = 10'h2da == r_count_1_io_out ? io_r_730_b : _GEN_1569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1571 = 10'h2db == r_count_1_io_out ? io_r_731_b : _GEN_1570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1572 = 10'h2dc == r_count_1_io_out ? io_r_732_b : _GEN_1571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1573 = 10'h2dd == r_count_1_io_out ? io_r_733_b : _GEN_1572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1574 = 10'h2de == r_count_1_io_out ? io_r_734_b : _GEN_1573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1575 = 10'h2df == r_count_1_io_out ? io_r_735_b : _GEN_1574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1576 = 10'h2e0 == r_count_1_io_out ? io_r_736_b : _GEN_1575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1577 = 10'h2e1 == r_count_1_io_out ? io_r_737_b : _GEN_1576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1578 = 10'h2e2 == r_count_1_io_out ? io_r_738_b : _GEN_1577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1579 = 10'h2e3 == r_count_1_io_out ? io_r_739_b : _GEN_1578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1580 = 10'h2e4 == r_count_1_io_out ? io_r_740_b : _GEN_1579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1581 = 10'h2e5 == r_count_1_io_out ? io_r_741_b : _GEN_1580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1582 = 10'h2e6 == r_count_1_io_out ? io_r_742_b : _GEN_1581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1583 = 10'h2e7 == r_count_1_io_out ? io_r_743_b : _GEN_1582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1584 = 10'h2e8 == r_count_1_io_out ? io_r_744_b : _GEN_1583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1585 = 10'h2e9 == r_count_1_io_out ? io_r_745_b : _GEN_1584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1586 = 10'h2ea == r_count_1_io_out ? io_r_746_b : _GEN_1585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1587 = 10'h2eb == r_count_1_io_out ? io_r_747_b : _GEN_1586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1588 = 10'h2ec == r_count_1_io_out ? io_r_748_b : _GEN_1587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1591 = 10'h1 == r_count_2_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1592 = 10'h2 == r_count_2_io_out ? io_r_2_b : _GEN_1591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1593 = 10'h3 == r_count_2_io_out ? io_r_3_b : _GEN_1592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1594 = 10'h4 == r_count_2_io_out ? io_r_4_b : _GEN_1593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1595 = 10'h5 == r_count_2_io_out ? io_r_5_b : _GEN_1594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1596 = 10'h6 == r_count_2_io_out ? io_r_6_b : _GEN_1595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1597 = 10'h7 == r_count_2_io_out ? io_r_7_b : _GEN_1596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1598 = 10'h8 == r_count_2_io_out ? io_r_8_b : _GEN_1597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1599 = 10'h9 == r_count_2_io_out ? io_r_9_b : _GEN_1598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1600 = 10'ha == r_count_2_io_out ? io_r_10_b : _GEN_1599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1601 = 10'hb == r_count_2_io_out ? io_r_11_b : _GEN_1600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1602 = 10'hc == r_count_2_io_out ? io_r_12_b : _GEN_1601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1603 = 10'hd == r_count_2_io_out ? io_r_13_b : _GEN_1602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1604 = 10'he == r_count_2_io_out ? io_r_14_b : _GEN_1603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1605 = 10'hf == r_count_2_io_out ? io_r_15_b : _GEN_1604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1606 = 10'h10 == r_count_2_io_out ? io_r_16_b : _GEN_1605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1607 = 10'h11 == r_count_2_io_out ? io_r_17_b : _GEN_1606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1608 = 10'h12 == r_count_2_io_out ? io_r_18_b : _GEN_1607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1609 = 10'h13 == r_count_2_io_out ? io_r_19_b : _GEN_1608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1610 = 10'h14 == r_count_2_io_out ? io_r_20_b : _GEN_1609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1611 = 10'h15 == r_count_2_io_out ? io_r_21_b : _GEN_1610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1612 = 10'h16 == r_count_2_io_out ? io_r_22_b : _GEN_1611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1613 = 10'h17 == r_count_2_io_out ? io_r_23_b : _GEN_1612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1614 = 10'h18 == r_count_2_io_out ? io_r_24_b : _GEN_1613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1615 = 10'h19 == r_count_2_io_out ? io_r_25_b : _GEN_1614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1616 = 10'h1a == r_count_2_io_out ? io_r_26_b : _GEN_1615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1617 = 10'h1b == r_count_2_io_out ? io_r_27_b : _GEN_1616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1618 = 10'h1c == r_count_2_io_out ? io_r_28_b : _GEN_1617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1619 = 10'h1d == r_count_2_io_out ? io_r_29_b : _GEN_1618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1620 = 10'h1e == r_count_2_io_out ? io_r_30_b : _GEN_1619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1621 = 10'h1f == r_count_2_io_out ? io_r_31_b : _GEN_1620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1622 = 10'h20 == r_count_2_io_out ? io_r_32_b : _GEN_1621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1623 = 10'h21 == r_count_2_io_out ? io_r_33_b : _GEN_1622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1624 = 10'h22 == r_count_2_io_out ? io_r_34_b : _GEN_1623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1625 = 10'h23 == r_count_2_io_out ? io_r_35_b : _GEN_1624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1626 = 10'h24 == r_count_2_io_out ? io_r_36_b : _GEN_1625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1627 = 10'h25 == r_count_2_io_out ? io_r_37_b : _GEN_1626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1628 = 10'h26 == r_count_2_io_out ? io_r_38_b : _GEN_1627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1629 = 10'h27 == r_count_2_io_out ? io_r_39_b : _GEN_1628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1630 = 10'h28 == r_count_2_io_out ? io_r_40_b : _GEN_1629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1631 = 10'h29 == r_count_2_io_out ? io_r_41_b : _GEN_1630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1632 = 10'h2a == r_count_2_io_out ? io_r_42_b : _GEN_1631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1633 = 10'h2b == r_count_2_io_out ? io_r_43_b : _GEN_1632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1634 = 10'h2c == r_count_2_io_out ? io_r_44_b : _GEN_1633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1635 = 10'h2d == r_count_2_io_out ? io_r_45_b : _GEN_1634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1636 = 10'h2e == r_count_2_io_out ? io_r_46_b : _GEN_1635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1637 = 10'h2f == r_count_2_io_out ? io_r_47_b : _GEN_1636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1638 = 10'h30 == r_count_2_io_out ? io_r_48_b : _GEN_1637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1639 = 10'h31 == r_count_2_io_out ? io_r_49_b : _GEN_1638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1640 = 10'h32 == r_count_2_io_out ? io_r_50_b : _GEN_1639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1641 = 10'h33 == r_count_2_io_out ? io_r_51_b : _GEN_1640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1642 = 10'h34 == r_count_2_io_out ? io_r_52_b : _GEN_1641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1643 = 10'h35 == r_count_2_io_out ? io_r_53_b : _GEN_1642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1644 = 10'h36 == r_count_2_io_out ? io_r_54_b : _GEN_1643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1645 = 10'h37 == r_count_2_io_out ? io_r_55_b : _GEN_1644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1646 = 10'h38 == r_count_2_io_out ? io_r_56_b : _GEN_1645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1647 = 10'h39 == r_count_2_io_out ? io_r_57_b : _GEN_1646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1648 = 10'h3a == r_count_2_io_out ? io_r_58_b : _GEN_1647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1649 = 10'h3b == r_count_2_io_out ? io_r_59_b : _GEN_1648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1650 = 10'h3c == r_count_2_io_out ? io_r_60_b : _GEN_1649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1651 = 10'h3d == r_count_2_io_out ? io_r_61_b : _GEN_1650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1652 = 10'h3e == r_count_2_io_out ? io_r_62_b : _GEN_1651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1653 = 10'h3f == r_count_2_io_out ? io_r_63_b : _GEN_1652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1654 = 10'h40 == r_count_2_io_out ? io_r_64_b : _GEN_1653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1655 = 10'h41 == r_count_2_io_out ? io_r_65_b : _GEN_1654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1656 = 10'h42 == r_count_2_io_out ? io_r_66_b : _GEN_1655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1657 = 10'h43 == r_count_2_io_out ? io_r_67_b : _GEN_1656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1658 = 10'h44 == r_count_2_io_out ? io_r_68_b : _GEN_1657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1659 = 10'h45 == r_count_2_io_out ? io_r_69_b : _GEN_1658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1660 = 10'h46 == r_count_2_io_out ? io_r_70_b : _GEN_1659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1661 = 10'h47 == r_count_2_io_out ? io_r_71_b : _GEN_1660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1662 = 10'h48 == r_count_2_io_out ? io_r_72_b : _GEN_1661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1663 = 10'h49 == r_count_2_io_out ? io_r_73_b : _GEN_1662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1664 = 10'h4a == r_count_2_io_out ? io_r_74_b : _GEN_1663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1665 = 10'h4b == r_count_2_io_out ? io_r_75_b : _GEN_1664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1666 = 10'h4c == r_count_2_io_out ? io_r_76_b : _GEN_1665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1667 = 10'h4d == r_count_2_io_out ? io_r_77_b : _GEN_1666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1668 = 10'h4e == r_count_2_io_out ? io_r_78_b : _GEN_1667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1669 = 10'h4f == r_count_2_io_out ? io_r_79_b : _GEN_1668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1670 = 10'h50 == r_count_2_io_out ? io_r_80_b : _GEN_1669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1671 = 10'h51 == r_count_2_io_out ? io_r_81_b : _GEN_1670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1672 = 10'h52 == r_count_2_io_out ? io_r_82_b : _GEN_1671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1673 = 10'h53 == r_count_2_io_out ? io_r_83_b : _GEN_1672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1674 = 10'h54 == r_count_2_io_out ? io_r_84_b : _GEN_1673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1675 = 10'h55 == r_count_2_io_out ? io_r_85_b : _GEN_1674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1676 = 10'h56 == r_count_2_io_out ? io_r_86_b : _GEN_1675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1677 = 10'h57 == r_count_2_io_out ? io_r_87_b : _GEN_1676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1678 = 10'h58 == r_count_2_io_out ? io_r_88_b : _GEN_1677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1679 = 10'h59 == r_count_2_io_out ? io_r_89_b : _GEN_1678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1680 = 10'h5a == r_count_2_io_out ? io_r_90_b : _GEN_1679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1681 = 10'h5b == r_count_2_io_out ? io_r_91_b : _GEN_1680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1682 = 10'h5c == r_count_2_io_out ? io_r_92_b : _GEN_1681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1683 = 10'h5d == r_count_2_io_out ? io_r_93_b : _GEN_1682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1684 = 10'h5e == r_count_2_io_out ? io_r_94_b : _GEN_1683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1685 = 10'h5f == r_count_2_io_out ? io_r_95_b : _GEN_1684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1686 = 10'h60 == r_count_2_io_out ? io_r_96_b : _GEN_1685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1687 = 10'h61 == r_count_2_io_out ? io_r_97_b : _GEN_1686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1688 = 10'h62 == r_count_2_io_out ? io_r_98_b : _GEN_1687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1689 = 10'h63 == r_count_2_io_out ? io_r_99_b : _GEN_1688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1690 = 10'h64 == r_count_2_io_out ? io_r_100_b : _GEN_1689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1691 = 10'h65 == r_count_2_io_out ? io_r_101_b : _GEN_1690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1692 = 10'h66 == r_count_2_io_out ? io_r_102_b : _GEN_1691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1693 = 10'h67 == r_count_2_io_out ? io_r_103_b : _GEN_1692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1694 = 10'h68 == r_count_2_io_out ? io_r_104_b : _GEN_1693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1695 = 10'h69 == r_count_2_io_out ? io_r_105_b : _GEN_1694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1696 = 10'h6a == r_count_2_io_out ? io_r_106_b : _GEN_1695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1697 = 10'h6b == r_count_2_io_out ? io_r_107_b : _GEN_1696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1698 = 10'h6c == r_count_2_io_out ? io_r_108_b : _GEN_1697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1699 = 10'h6d == r_count_2_io_out ? io_r_109_b : _GEN_1698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1700 = 10'h6e == r_count_2_io_out ? io_r_110_b : _GEN_1699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1701 = 10'h6f == r_count_2_io_out ? io_r_111_b : _GEN_1700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1702 = 10'h70 == r_count_2_io_out ? io_r_112_b : _GEN_1701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1703 = 10'h71 == r_count_2_io_out ? io_r_113_b : _GEN_1702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1704 = 10'h72 == r_count_2_io_out ? io_r_114_b : _GEN_1703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1705 = 10'h73 == r_count_2_io_out ? io_r_115_b : _GEN_1704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1706 = 10'h74 == r_count_2_io_out ? io_r_116_b : _GEN_1705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1707 = 10'h75 == r_count_2_io_out ? io_r_117_b : _GEN_1706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1708 = 10'h76 == r_count_2_io_out ? io_r_118_b : _GEN_1707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1709 = 10'h77 == r_count_2_io_out ? io_r_119_b : _GEN_1708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1710 = 10'h78 == r_count_2_io_out ? io_r_120_b : _GEN_1709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1711 = 10'h79 == r_count_2_io_out ? io_r_121_b : _GEN_1710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1712 = 10'h7a == r_count_2_io_out ? io_r_122_b : _GEN_1711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1713 = 10'h7b == r_count_2_io_out ? io_r_123_b : _GEN_1712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1714 = 10'h7c == r_count_2_io_out ? io_r_124_b : _GEN_1713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1715 = 10'h7d == r_count_2_io_out ? io_r_125_b : _GEN_1714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1716 = 10'h7e == r_count_2_io_out ? io_r_126_b : _GEN_1715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1717 = 10'h7f == r_count_2_io_out ? io_r_127_b : _GEN_1716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1718 = 10'h80 == r_count_2_io_out ? io_r_128_b : _GEN_1717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1719 = 10'h81 == r_count_2_io_out ? io_r_129_b : _GEN_1718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1720 = 10'h82 == r_count_2_io_out ? io_r_130_b : _GEN_1719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1721 = 10'h83 == r_count_2_io_out ? io_r_131_b : _GEN_1720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1722 = 10'h84 == r_count_2_io_out ? io_r_132_b : _GEN_1721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1723 = 10'h85 == r_count_2_io_out ? io_r_133_b : _GEN_1722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1724 = 10'h86 == r_count_2_io_out ? io_r_134_b : _GEN_1723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1725 = 10'h87 == r_count_2_io_out ? io_r_135_b : _GEN_1724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1726 = 10'h88 == r_count_2_io_out ? io_r_136_b : _GEN_1725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1727 = 10'h89 == r_count_2_io_out ? io_r_137_b : _GEN_1726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1728 = 10'h8a == r_count_2_io_out ? io_r_138_b : _GEN_1727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1729 = 10'h8b == r_count_2_io_out ? io_r_139_b : _GEN_1728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1730 = 10'h8c == r_count_2_io_out ? io_r_140_b : _GEN_1729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1731 = 10'h8d == r_count_2_io_out ? io_r_141_b : _GEN_1730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1732 = 10'h8e == r_count_2_io_out ? io_r_142_b : _GEN_1731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1733 = 10'h8f == r_count_2_io_out ? io_r_143_b : _GEN_1732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1734 = 10'h90 == r_count_2_io_out ? io_r_144_b : _GEN_1733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1735 = 10'h91 == r_count_2_io_out ? io_r_145_b : _GEN_1734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1736 = 10'h92 == r_count_2_io_out ? io_r_146_b : _GEN_1735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1737 = 10'h93 == r_count_2_io_out ? io_r_147_b : _GEN_1736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1738 = 10'h94 == r_count_2_io_out ? io_r_148_b : _GEN_1737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1739 = 10'h95 == r_count_2_io_out ? io_r_149_b : _GEN_1738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1740 = 10'h96 == r_count_2_io_out ? io_r_150_b : _GEN_1739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1741 = 10'h97 == r_count_2_io_out ? io_r_151_b : _GEN_1740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1742 = 10'h98 == r_count_2_io_out ? io_r_152_b : _GEN_1741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1743 = 10'h99 == r_count_2_io_out ? io_r_153_b : _GEN_1742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1744 = 10'h9a == r_count_2_io_out ? io_r_154_b : _GEN_1743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1745 = 10'h9b == r_count_2_io_out ? io_r_155_b : _GEN_1744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1746 = 10'h9c == r_count_2_io_out ? io_r_156_b : _GEN_1745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1747 = 10'h9d == r_count_2_io_out ? io_r_157_b : _GEN_1746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1748 = 10'h9e == r_count_2_io_out ? io_r_158_b : _GEN_1747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1749 = 10'h9f == r_count_2_io_out ? io_r_159_b : _GEN_1748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1750 = 10'ha0 == r_count_2_io_out ? io_r_160_b : _GEN_1749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1751 = 10'ha1 == r_count_2_io_out ? io_r_161_b : _GEN_1750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1752 = 10'ha2 == r_count_2_io_out ? io_r_162_b : _GEN_1751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1753 = 10'ha3 == r_count_2_io_out ? io_r_163_b : _GEN_1752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1754 = 10'ha4 == r_count_2_io_out ? io_r_164_b : _GEN_1753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1755 = 10'ha5 == r_count_2_io_out ? io_r_165_b : _GEN_1754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1756 = 10'ha6 == r_count_2_io_out ? io_r_166_b : _GEN_1755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1757 = 10'ha7 == r_count_2_io_out ? io_r_167_b : _GEN_1756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1758 = 10'ha8 == r_count_2_io_out ? io_r_168_b : _GEN_1757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1759 = 10'ha9 == r_count_2_io_out ? io_r_169_b : _GEN_1758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1760 = 10'haa == r_count_2_io_out ? io_r_170_b : _GEN_1759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1761 = 10'hab == r_count_2_io_out ? io_r_171_b : _GEN_1760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1762 = 10'hac == r_count_2_io_out ? io_r_172_b : _GEN_1761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1763 = 10'had == r_count_2_io_out ? io_r_173_b : _GEN_1762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1764 = 10'hae == r_count_2_io_out ? io_r_174_b : _GEN_1763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1765 = 10'haf == r_count_2_io_out ? io_r_175_b : _GEN_1764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1766 = 10'hb0 == r_count_2_io_out ? io_r_176_b : _GEN_1765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1767 = 10'hb1 == r_count_2_io_out ? io_r_177_b : _GEN_1766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1768 = 10'hb2 == r_count_2_io_out ? io_r_178_b : _GEN_1767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1769 = 10'hb3 == r_count_2_io_out ? io_r_179_b : _GEN_1768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1770 = 10'hb4 == r_count_2_io_out ? io_r_180_b : _GEN_1769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1771 = 10'hb5 == r_count_2_io_out ? io_r_181_b : _GEN_1770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1772 = 10'hb6 == r_count_2_io_out ? io_r_182_b : _GEN_1771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1773 = 10'hb7 == r_count_2_io_out ? io_r_183_b : _GEN_1772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1774 = 10'hb8 == r_count_2_io_out ? io_r_184_b : _GEN_1773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1775 = 10'hb9 == r_count_2_io_out ? io_r_185_b : _GEN_1774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1776 = 10'hba == r_count_2_io_out ? io_r_186_b : _GEN_1775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1777 = 10'hbb == r_count_2_io_out ? io_r_187_b : _GEN_1776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1778 = 10'hbc == r_count_2_io_out ? io_r_188_b : _GEN_1777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1779 = 10'hbd == r_count_2_io_out ? io_r_189_b : _GEN_1778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1780 = 10'hbe == r_count_2_io_out ? io_r_190_b : _GEN_1779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1781 = 10'hbf == r_count_2_io_out ? io_r_191_b : _GEN_1780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1782 = 10'hc0 == r_count_2_io_out ? io_r_192_b : _GEN_1781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1783 = 10'hc1 == r_count_2_io_out ? io_r_193_b : _GEN_1782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1784 = 10'hc2 == r_count_2_io_out ? io_r_194_b : _GEN_1783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1785 = 10'hc3 == r_count_2_io_out ? io_r_195_b : _GEN_1784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1786 = 10'hc4 == r_count_2_io_out ? io_r_196_b : _GEN_1785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1787 = 10'hc5 == r_count_2_io_out ? io_r_197_b : _GEN_1786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1788 = 10'hc6 == r_count_2_io_out ? io_r_198_b : _GEN_1787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1789 = 10'hc7 == r_count_2_io_out ? io_r_199_b : _GEN_1788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1790 = 10'hc8 == r_count_2_io_out ? io_r_200_b : _GEN_1789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1791 = 10'hc9 == r_count_2_io_out ? io_r_201_b : _GEN_1790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1792 = 10'hca == r_count_2_io_out ? io_r_202_b : _GEN_1791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1793 = 10'hcb == r_count_2_io_out ? io_r_203_b : _GEN_1792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1794 = 10'hcc == r_count_2_io_out ? io_r_204_b : _GEN_1793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1795 = 10'hcd == r_count_2_io_out ? io_r_205_b : _GEN_1794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1796 = 10'hce == r_count_2_io_out ? io_r_206_b : _GEN_1795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1797 = 10'hcf == r_count_2_io_out ? io_r_207_b : _GEN_1796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1798 = 10'hd0 == r_count_2_io_out ? io_r_208_b : _GEN_1797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1799 = 10'hd1 == r_count_2_io_out ? io_r_209_b : _GEN_1798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1800 = 10'hd2 == r_count_2_io_out ? io_r_210_b : _GEN_1799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1801 = 10'hd3 == r_count_2_io_out ? io_r_211_b : _GEN_1800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1802 = 10'hd4 == r_count_2_io_out ? io_r_212_b : _GEN_1801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1803 = 10'hd5 == r_count_2_io_out ? io_r_213_b : _GEN_1802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1804 = 10'hd6 == r_count_2_io_out ? io_r_214_b : _GEN_1803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1805 = 10'hd7 == r_count_2_io_out ? io_r_215_b : _GEN_1804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1806 = 10'hd8 == r_count_2_io_out ? io_r_216_b : _GEN_1805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1807 = 10'hd9 == r_count_2_io_out ? io_r_217_b : _GEN_1806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1808 = 10'hda == r_count_2_io_out ? io_r_218_b : _GEN_1807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1809 = 10'hdb == r_count_2_io_out ? io_r_219_b : _GEN_1808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1810 = 10'hdc == r_count_2_io_out ? io_r_220_b : _GEN_1809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1811 = 10'hdd == r_count_2_io_out ? io_r_221_b : _GEN_1810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1812 = 10'hde == r_count_2_io_out ? io_r_222_b : _GEN_1811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1813 = 10'hdf == r_count_2_io_out ? io_r_223_b : _GEN_1812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1814 = 10'he0 == r_count_2_io_out ? io_r_224_b : _GEN_1813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1815 = 10'he1 == r_count_2_io_out ? io_r_225_b : _GEN_1814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1816 = 10'he2 == r_count_2_io_out ? io_r_226_b : _GEN_1815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1817 = 10'he3 == r_count_2_io_out ? io_r_227_b : _GEN_1816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1818 = 10'he4 == r_count_2_io_out ? io_r_228_b : _GEN_1817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1819 = 10'he5 == r_count_2_io_out ? io_r_229_b : _GEN_1818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1820 = 10'he6 == r_count_2_io_out ? io_r_230_b : _GEN_1819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1821 = 10'he7 == r_count_2_io_out ? io_r_231_b : _GEN_1820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1822 = 10'he8 == r_count_2_io_out ? io_r_232_b : _GEN_1821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1823 = 10'he9 == r_count_2_io_out ? io_r_233_b : _GEN_1822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1824 = 10'hea == r_count_2_io_out ? io_r_234_b : _GEN_1823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1825 = 10'heb == r_count_2_io_out ? io_r_235_b : _GEN_1824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1826 = 10'hec == r_count_2_io_out ? io_r_236_b : _GEN_1825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1827 = 10'hed == r_count_2_io_out ? io_r_237_b : _GEN_1826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1828 = 10'hee == r_count_2_io_out ? io_r_238_b : _GEN_1827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1829 = 10'hef == r_count_2_io_out ? io_r_239_b : _GEN_1828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1830 = 10'hf0 == r_count_2_io_out ? io_r_240_b : _GEN_1829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1831 = 10'hf1 == r_count_2_io_out ? io_r_241_b : _GEN_1830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1832 = 10'hf2 == r_count_2_io_out ? io_r_242_b : _GEN_1831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1833 = 10'hf3 == r_count_2_io_out ? io_r_243_b : _GEN_1832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1834 = 10'hf4 == r_count_2_io_out ? io_r_244_b : _GEN_1833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1835 = 10'hf5 == r_count_2_io_out ? io_r_245_b : _GEN_1834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1836 = 10'hf6 == r_count_2_io_out ? io_r_246_b : _GEN_1835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1837 = 10'hf7 == r_count_2_io_out ? io_r_247_b : _GEN_1836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1838 = 10'hf8 == r_count_2_io_out ? io_r_248_b : _GEN_1837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1839 = 10'hf9 == r_count_2_io_out ? io_r_249_b : _GEN_1838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1840 = 10'hfa == r_count_2_io_out ? io_r_250_b : _GEN_1839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1841 = 10'hfb == r_count_2_io_out ? io_r_251_b : _GEN_1840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1842 = 10'hfc == r_count_2_io_out ? io_r_252_b : _GEN_1841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1843 = 10'hfd == r_count_2_io_out ? io_r_253_b : _GEN_1842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1844 = 10'hfe == r_count_2_io_out ? io_r_254_b : _GEN_1843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1845 = 10'hff == r_count_2_io_out ? io_r_255_b : _GEN_1844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1846 = 10'h100 == r_count_2_io_out ? io_r_256_b : _GEN_1845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1847 = 10'h101 == r_count_2_io_out ? io_r_257_b : _GEN_1846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1848 = 10'h102 == r_count_2_io_out ? io_r_258_b : _GEN_1847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1849 = 10'h103 == r_count_2_io_out ? io_r_259_b : _GEN_1848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1850 = 10'h104 == r_count_2_io_out ? io_r_260_b : _GEN_1849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1851 = 10'h105 == r_count_2_io_out ? io_r_261_b : _GEN_1850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1852 = 10'h106 == r_count_2_io_out ? io_r_262_b : _GEN_1851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1853 = 10'h107 == r_count_2_io_out ? io_r_263_b : _GEN_1852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1854 = 10'h108 == r_count_2_io_out ? io_r_264_b : _GEN_1853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1855 = 10'h109 == r_count_2_io_out ? io_r_265_b : _GEN_1854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1856 = 10'h10a == r_count_2_io_out ? io_r_266_b : _GEN_1855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1857 = 10'h10b == r_count_2_io_out ? io_r_267_b : _GEN_1856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1858 = 10'h10c == r_count_2_io_out ? io_r_268_b : _GEN_1857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1859 = 10'h10d == r_count_2_io_out ? io_r_269_b : _GEN_1858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1860 = 10'h10e == r_count_2_io_out ? io_r_270_b : _GEN_1859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1861 = 10'h10f == r_count_2_io_out ? io_r_271_b : _GEN_1860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1862 = 10'h110 == r_count_2_io_out ? io_r_272_b : _GEN_1861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1863 = 10'h111 == r_count_2_io_out ? io_r_273_b : _GEN_1862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1864 = 10'h112 == r_count_2_io_out ? io_r_274_b : _GEN_1863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1865 = 10'h113 == r_count_2_io_out ? io_r_275_b : _GEN_1864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1866 = 10'h114 == r_count_2_io_out ? io_r_276_b : _GEN_1865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1867 = 10'h115 == r_count_2_io_out ? io_r_277_b : _GEN_1866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1868 = 10'h116 == r_count_2_io_out ? io_r_278_b : _GEN_1867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1869 = 10'h117 == r_count_2_io_out ? io_r_279_b : _GEN_1868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1870 = 10'h118 == r_count_2_io_out ? io_r_280_b : _GEN_1869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1871 = 10'h119 == r_count_2_io_out ? io_r_281_b : _GEN_1870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1872 = 10'h11a == r_count_2_io_out ? io_r_282_b : _GEN_1871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1873 = 10'h11b == r_count_2_io_out ? io_r_283_b : _GEN_1872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1874 = 10'h11c == r_count_2_io_out ? io_r_284_b : _GEN_1873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1875 = 10'h11d == r_count_2_io_out ? io_r_285_b : _GEN_1874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1876 = 10'h11e == r_count_2_io_out ? io_r_286_b : _GEN_1875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1877 = 10'h11f == r_count_2_io_out ? io_r_287_b : _GEN_1876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1878 = 10'h120 == r_count_2_io_out ? io_r_288_b : _GEN_1877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1879 = 10'h121 == r_count_2_io_out ? io_r_289_b : _GEN_1878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1880 = 10'h122 == r_count_2_io_out ? io_r_290_b : _GEN_1879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1881 = 10'h123 == r_count_2_io_out ? io_r_291_b : _GEN_1880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1882 = 10'h124 == r_count_2_io_out ? io_r_292_b : _GEN_1881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1883 = 10'h125 == r_count_2_io_out ? io_r_293_b : _GEN_1882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1884 = 10'h126 == r_count_2_io_out ? io_r_294_b : _GEN_1883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1885 = 10'h127 == r_count_2_io_out ? io_r_295_b : _GEN_1884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1886 = 10'h128 == r_count_2_io_out ? io_r_296_b : _GEN_1885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1887 = 10'h129 == r_count_2_io_out ? io_r_297_b : _GEN_1886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1888 = 10'h12a == r_count_2_io_out ? io_r_298_b : _GEN_1887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1889 = 10'h12b == r_count_2_io_out ? io_r_299_b : _GEN_1888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1890 = 10'h12c == r_count_2_io_out ? io_r_300_b : _GEN_1889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1891 = 10'h12d == r_count_2_io_out ? io_r_301_b : _GEN_1890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1892 = 10'h12e == r_count_2_io_out ? io_r_302_b : _GEN_1891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1893 = 10'h12f == r_count_2_io_out ? io_r_303_b : _GEN_1892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1894 = 10'h130 == r_count_2_io_out ? io_r_304_b : _GEN_1893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1895 = 10'h131 == r_count_2_io_out ? io_r_305_b : _GEN_1894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1896 = 10'h132 == r_count_2_io_out ? io_r_306_b : _GEN_1895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1897 = 10'h133 == r_count_2_io_out ? io_r_307_b : _GEN_1896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1898 = 10'h134 == r_count_2_io_out ? io_r_308_b : _GEN_1897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1899 = 10'h135 == r_count_2_io_out ? io_r_309_b : _GEN_1898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1900 = 10'h136 == r_count_2_io_out ? io_r_310_b : _GEN_1899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1901 = 10'h137 == r_count_2_io_out ? io_r_311_b : _GEN_1900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1902 = 10'h138 == r_count_2_io_out ? io_r_312_b : _GEN_1901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1903 = 10'h139 == r_count_2_io_out ? io_r_313_b : _GEN_1902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1904 = 10'h13a == r_count_2_io_out ? io_r_314_b : _GEN_1903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1905 = 10'h13b == r_count_2_io_out ? io_r_315_b : _GEN_1904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1906 = 10'h13c == r_count_2_io_out ? io_r_316_b : _GEN_1905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1907 = 10'h13d == r_count_2_io_out ? io_r_317_b : _GEN_1906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1908 = 10'h13e == r_count_2_io_out ? io_r_318_b : _GEN_1907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1909 = 10'h13f == r_count_2_io_out ? io_r_319_b : _GEN_1908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1910 = 10'h140 == r_count_2_io_out ? io_r_320_b : _GEN_1909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1911 = 10'h141 == r_count_2_io_out ? io_r_321_b : _GEN_1910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1912 = 10'h142 == r_count_2_io_out ? io_r_322_b : _GEN_1911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1913 = 10'h143 == r_count_2_io_out ? io_r_323_b : _GEN_1912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1914 = 10'h144 == r_count_2_io_out ? io_r_324_b : _GEN_1913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1915 = 10'h145 == r_count_2_io_out ? io_r_325_b : _GEN_1914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1916 = 10'h146 == r_count_2_io_out ? io_r_326_b : _GEN_1915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1917 = 10'h147 == r_count_2_io_out ? io_r_327_b : _GEN_1916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1918 = 10'h148 == r_count_2_io_out ? io_r_328_b : _GEN_1917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1919 = 10'h149 == r_count_2_io_out ? io_r_329_b : _GEN_1918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1920 = 10'h14a == r_count_2_io_out ? io_r_330_b : _GEN_1919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1921 = 10'h14b == r_count_2_io_out ? io_r_331_b : _GEN_1920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1922 = 10'h14c == r_count_2_io_out ? io_r_332_b : _GEN_1921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1923 = 10'h14d == r_count_2_io_out ? io_r_333_b : _GEN_1922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1924 = 10'h14e == r_count_2_io_out ? io_r_334_b : _GEN_1923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1925 = 10'h14f == r_count_2_io_out ? io_r_335_b : _GEN_1924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1926 = 10'h150 == r_count_2_io_out ? io_r_336_b : _GEN_1925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1927 = 10'h151 == r_count_2_io_out ? io_r_337_b : _GEN_1926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1928 = 10'h152 == r_count_2_io_out ? io_r_338_b : _GEN_1927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1929 = 10'h153 == r_count_2_io_out ? io_r_339_b : _GEN_1928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1930 = 10'h154 == r_count_2_io_out ? io_r_340_b : _GEN_1929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1931 = 10'h155 == r_count_2_io_out ? io_r_341_b : _GEN_1930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1932 = 10'h156 == r_count_2_io_out ? io_r_342_b : _GEN_1931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1933 = 10'h157 == r_count_2_io_out ? io_r_343_b : _GEN_1932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1934 = 10'h158 == r_count_2_io_out ? io_r_344_b : _GEN_1933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1935 = 10'h159 == r_count_2_io_out ? io_r_345_b : _GEN_1934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1936 = 10'h15a == r_count_2_io_out ? io_r_346_b : _GEN_1935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1937 = 10'h15b == r_count_2_io_out ? io_r_347_b : _GEN_1936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1938 = 10'h15c == r_count_2_io_out ? io_r_348_b : _GEN_1937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1939 = 10'h15d == r_count_2_io_out ? io_r_349_b : _GEN_1938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1940 = 10'h15e == r_count_2_io_out ? io_r_350_b : _GEN_1939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1941 = 10'h15f == r_count_2_io_out ? io_r_351_b : _GEN_1940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1942 = 10'h160 == r_count_2_io_out ? io_r_352_b : _GEN_1941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1943 = 10'h161 == r_count_2_io_out ? io_r_353_b : _GEN_1942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1944 = 10'h162 == r_count_2_io_out ? io_r_354_b : _GEN_1943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1945 = 10'h163 == r_count_2_io_out ? io_r_355_b : _GEN_1944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1946 = 10'h164 == r_count_2_io_out ? io_r_356_b : _GEN_1945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1947 = 10'h165 == r_count_2_io_out ? io_r_357_b : _GEN_1946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1948 = 10'h166 == r_count_2_io_out ? io_r_358_b : _GEN_1947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1949 = 10'h167 == r_count_2_io_out ? io_r_359_b : _GEN_1948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1950 = 10'h168 == r_count_2_io_out ? io_r_360_b : _GEN_1949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1951 = 10'h169 == r_count_2_io_out ? io_r_361_b : _GEN_1950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1952 = 10'h16a == r_count_2_io_out ? io_r_362_b : _GEN_1951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1953 = 10'h16b == r_count_2_io_out ? io_r_363_b : _GEN_1952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1954 = 10'h16c == r_count_2_io_out ? io_r_364_b : _GEN_1953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1955 = 10'h16d == r_count_2_io_out ? io_r_365_b : _GEN_1954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1956 = 10'h16e == r_count_2_io_out ? io_r_366_b : _GEN_1955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1957 = 10'h16f == r_count_2_io_out ? io_r_367_b : _GEN_1956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1958 = 10'h170 == r_count_2_io_out ? io_r_368_b : _GEN_1957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1959 = 10'h171 == r_count_2_io_out ? io_r_369_b : _GEN_1958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1960 = 10'h172 == r_count_2_io_out ? io_r_370_b : _GEN_1959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1961 = 10'h173 == r_count_2_io_out ? io_r_371_b : _GEN_1960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1962 = 10'h174 == r_count_2_io_out ? io_r_372_b : _GEN_1961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1963 = 10'h175 == r_count_2_io_out ? io_r_373_b : _GEN_1962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1964 = 10'h176 == r_count_2_io_out ? io_r_374_b : _GEN_1963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1965 = 10'h177 == r_count_2_io_out ? io_r_375_b : _GEN_1964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1966 = 10'h178 == r_count_2_io_out ? io_r_376_b : _GEN_1965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1967 = 10'h179 == r_count_2_io_out ? io_r_377_b : _GEN_1966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1968 = 10'h17a == r_count_2_io_out ? io_r_378_b : _GEN_1967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1969 = 10'h17b == r_count_2_io_out ? io_r_379_b : _GEN_1968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1970 = 10'h17c == r_count_2_io_out ? io_r_380_b : _GEN_1969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1971 = 10'h17d == r_count_2_io_out ? io_r_381_b : _GEN_1970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1972 = 10'h17e == r_count_2_io_out ? io_r_382_b : _GEN_1971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1973 = 10'h17f == r_count_2_io_out ? io_r_383_b : _GEN_1972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1974 = 10'h180 == r_count_2_io_out ? io_r_384_b : _GEN_1973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1975 = 10'h181 == r_count_2_io_out ? io_r_385_b : _GEN_1974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1976 = 10'h182 == r_count_2_io_out ? io_r_386_b : _GEN_1975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1977 = 10'h183 == r_count_2_io_out ? io_r_387_b : _GEN_1976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1978 = 10'h184 == r_count_2_io_out ? io_r_388_b : _GEN_1977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1979 = 10'h185 == r_count_2_io_out ? io_r_389_b : _GEN_1978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1980 = 10'h186 == r_count_2_io_out ? io_r_390_b : _GEN_1979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1981 = 10'h187 == r_count_2_io_out ? io_r_391_b : _GEN_1980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1982 = 10'h188 == r_count_2_io_out ? io_r_392_b : _GEN_1981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1983 = 10'h189 == r_count_2_io_out ? io_r_393_b : _GEN_1982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1984 = 10'h18a == r_count_2_io_out ? io_r_394_b : _GEN_1983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1985 = 10'h18b == r_count_2_io_out ? io_r_395_b : _GEN_1984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1986 = 10'h18c == r_count_2_io_out ? io_r_396_b : _GEN_1985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1987 = 10'h18d == r_count_2_io_out ? io_r_397_b : _GEN_1986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1988 = 10'h18e == r_count_2_io_out ? io_r_398_b : _GEN_1987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1989 = 10'h18f == r_count_2_io_out ? io_r_399_b : _GEN_1988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1990 = 10'h190 == r_count_2_io_out ? io_r_400_b : _GEN_1989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1991 = 10'h191 == r_count_2_io_out ? io_r_401_b : _GEN_1990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1992 = 10'h192 == r_count_2_io_out ? io_r_402_b : _GEN_1991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1993 = 10'h193 == r_count_2_io_out ? io_r_403_b : _GEN_1992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1994 = 10'h194 == r_count_2_io_out ? io_r_404_b : _GEN_1993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1995 = 10'h195 == r_count_2_io_out ? io_r_405_b : _GEN_1994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1996 = 10'h196 == r_count_2_io_out ? io_r_406_b : _GEN_1995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1997 = 10'h197 == r_count_2_io_out ? io_r_407_b : _GEN_1996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1998 = 10'h198 == r_count_2_io_out ? io_r_408_b : _GEN_1997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1999 = 10'h199 == r_count_2_io_out ? io_r_409_b : _GEN_1998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2000 = 10'h19a == r_count_2_io_out ? io_r_410_b : _GEN_1999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2001 = 10'h19b == r_count_2_io_out ? io_r_411_b : _GEN_2000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2002 = 10'h19c == r_count_2_io_out ? io_r_412_b : _GEN_2001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2003 = 10'h19d == r_count_2_io_out ? io_r_413_b : _GEN_2002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2004 = 10'h19e == r_count_2_io_out ? io_r_414_b : _GEN_2003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2005 = 10'h19f == r_count_2_io_out ? io_r_415_b : _GEN_2004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2006 = 10'h1a0 == r_count_2_io_out ? io_r_416_b : _GEN_2005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2007 = 10'h1a1 == r_count_2_io_out ? io_r_417_b : _GEN_2006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2008 = 10'h1a2 == r_count_2_io_out ? io_r_418_b : _GEN_2007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2009 = 10'h1a3 == r_count_2_io_out ? io_r_419_b : _GEN_2008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2010 = 10'h1a4 == r_count_2_io_out ? io_r_420_b : _GEN_2009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2011 = 10'h1a5 == r_count_2_io_out ? io_r_421_b : _GEN_2010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2012 = 10'h1a6 == r_count_2_io_out ? io_r_422_b : _GEN_2011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2013 = 10'h1a7 == r_count_2_io_out ? io_r_423_b : _GEN_2012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2014 = 10'h1a8 == r_count_2_io_out ? io_r_424_b : _GEN_2013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2015 = 10'h1a9 == r_count_2_io_out ? io_r_425_b : _GEN_2014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2016 = 10'h1aa == r_count_2_io_out ? io_r_426_b : _GEN_2015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2017 = 10'h1ab == r_count_2_io_out ? io_r_427_b : _GEN_2016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2018 = 10'h1ac == r_count_2_io_out ? io_r_428_b : _GEN_2017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2019 = 10'h1ad == r_count_2_io_out ? io_r_429_b : _GEN_2018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2020 = 10'h1ae == r_count_2_io_out ? io_r_430_b : _GEN_2019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2021 = 10'h1af == r_count_2_io_out ? io_r_431_b : _GEN_2020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2022 = 10'h1b0 == r_count_2_io_out ? io_r_432_b : _GEN_2021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2023 = 10'h1b1 == r_count_2_io_out ? io_r_433_b : _GEN_2022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2024 = 10'h1b2 == r_count_2_io_out ? io_r_434_b : _GEN_2023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2025 = 10'h1b3 == r_count_2_io_out ? io_r_435_b : _GEN_2024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2026 = 10'h1b4 == r_count_2_io_out ? io_r_436_b : _GEN_2025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2027 = 10'h1b5 == r_count_2_io_out ? io_r_437_b : _GEN_2026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2028 = 10'h1b6 == r_count_2_io_out ? io_r_438_b : _GEN_2027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2029 = 10'h1b7 == r_count_2_io_out ? io_r_439_b : _GEN_2028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2030 = 10'h1b8 == r_count_2_io_out ? io_r_440_b : _GEN_2029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2031 = 10'h1b9 == r_count_2_io_out ? io_r_441_b : _GEN_2030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2032 = 10'h1ba == r_count_2_io_out ? io_r_442_b : _GEN_2031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2033 = 10'h1bb == r_count_2_io_out ? io_r_443_b : _GEN_2032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2034 = 10'h1bc == r_count_2_io_out ? io_r_444_b : _GEN_2033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2035 = 10'h1bd == r_count_2_io_out ? io_r_445_b : _GEN_2034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2036 = 10'h1be == r_count_2_io_out ? io_r_446_b : _GEN_2035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2037 = 10'h1bf == r_count_2_io_out ? io_r_447_b : _GEN_2036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2038 = 10'h1c0 == r_count_2_io_out ? io_r_448_b : _GEN_2037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2039 = 10'h1c1 == r_count_2_io_out ? io_r_449_b : _GEN_2038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2040 = 10'h1c2 == r_count_2_io_out ? io_r_450_b : _GEN_2039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2041 = 10'h1c3 == r_count_2_io_out ? io_r_451_b : _GEN_2040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2042 = 10'h1c4 == r_count_2_io_out ? io_r_452_b : _GEN_2041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2043 = 10'h1c5 == r_count_2_io_out ? io_r_453_b : _GEN_2042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2044 = 10'h1c6 == r_count_2_io_out ? io_r_454_b : _GEN_2043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2045 = 10'h1c7 == r_count_2_io_out ? io_r_455_b : _GEN_2044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2046 = 10'h1c8 == r_count_2_io_out ? io_r_456_b : _GEN_2045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2047 = 10'h1c9 == r_count_2_io_out ? io_r_457_b : _GEN_2046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2048 = 10'h1ca == r_count_2_io_out ? io_r_458_b : _GEN_2047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2049 = 10'h1cb == r_count_2_io_out ? io_r_459_b : _GEN_2048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2050 = 10'h1cc == r_count_2_io_out ? io_r_460_b : _GEN_2049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2051 = 10'h1cd == r_count_2_io_out ? io_r_461_b : _GEN_2050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2052 = 10'h1ce == r_count_2_io_out ? io_r_462_b : _GEN_2051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2053 = 10'h1cf == r_count_2_io_out ? io_r_463_b : _GEN_2052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2054 = 10'h1d0 == r_count_2_io_out ? io_r_464_b : _GEN_2053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2055 = 10'h1d1 == r_count_2_io_out ? io_r_465_b : _GEN_2054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2056 = 10'h1d2 == r_count_2_io_out ? io_r_466_b : _GEN_2055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2057 = 10'h1d3 == r_count_2_io_out ? io_r_467_b : _GEN_2056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2058 = 10'h1d4 == r_count_2_io_out ? io_r_468_b : _GEN_2057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2059 = 10'h1d5 == r_count_2_io_out ? io_r_469_b : _GEN_2058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2060 = 10'h1d6 == r_count_2_io_out ? io_r_470_b : _GEN_2059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2061 = 10'h1d7 == r_count_2_io_out ? io_r_471_b : _GEN_2060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2062 = 10'h1d8 == r_count_2_io_out ? io_r_472_b : _GEN_2061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2063 = 10'h1d9 == r_count_2_io_out ? io_r_473_b : _GEN_2062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2064 = 10'h1da == r_count_2_io_out ? io_r_474_b : _GEN_2063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2065 = 10'h1db == r_count_2_io_out ? io_r_475_b : _GEN_2064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2066 = 10'h1dc == r_count_2_io_out ? io_r_476_b : _GEN_2065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2067 = 10'h1dd == r_count_2_io_out ? io_r_477_b : _GEN_2066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2068 = 10'h1de == r_count_2_io_out ? io_r_478_b : _GEN_2067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2069 = 10'h1df == r_count_2_io_out ? io_r_479_b : _GEN_2068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2070 = 10'h1e0 == r_count_2_io_out ? io_r_480_b : _GEN_2069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2071 = 10'h1e1 == r_count_2_io_out ? io_r_481_b : _GEN_2070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2072 = 10'h1e2 == r_count_2_io_out ? io_r_482_b : _GEN_2071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2073 = 10'h1e3 == r_count_2_io_out ? io_r_483_b : _GEN_2072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2074 = 10'h1e4 == r_count_2_io_out ? io_r_484_b : _GEN_2073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2075 = 10'h1e5 == r_count_2_io_out ? io_r_485_b : _GEN_2074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2076 = 10'h1e6 == r_count_2_io_out ? io_r_486_b : _GEN_2075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2077 = 10'h1e7 == r_count_2_io_out ? io_r_487_b : _GEN_2076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2078 = 10'h1e8 == r_count_2_io_out ? io_r_488_b : _GEN_2077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2079 = 10'h1e9 == r_count_2_io_out ? io_r_489_b : _GEN_2078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2080 = 10'h1ea == r_count_2_io_out ? io_r_490_b : _GEN_2079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2081 = 10'h1eb == r_count_2_io_out ? io_r_491_b : _GEN_2080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2082 = 10'h1ec == r_count_2_io_out ? io_r_492_b : _GEN_2081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2083 = 10'h1ed == r_count_2_io_out ? io_r_493_b : _GEN_2082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2084 = 10'h1ee == r_count_2_io_out ? io_r_494_b : _GEN_2083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2085 = 10'h1ef == r_count_2_io_out ? io_r_495_b : _GEN_2084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2086 = 10'h1f0 == r_count_2_io_out ? io_r_496_b : _GEN_2085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2087 = 10'h1f1 == r_count_2_io_out ? io_r_497_b : _GEN_2086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2088 = 10'h1f2 == r_count_2_io_out ? io_r_498_b : _GEN_2087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2089 = 10'h1f3 == r_count_2_io_out ? io_r_499_b : _GEN_2088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2090 = 10'h1f4 == r_count_2_io_out ? io_r_500_b : _GEN_2089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2091 = 10'h1f5 == r_count_2_io_out ? io_r_501_b : _GEN_2090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2092 = 10'h1f6 == r_count_2_io_out ? io_r_502_b : _GEN_2091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2093 = 10'h1f7 == r_count_2_io_out ? io_r_503_b : _GEN_2092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2094 = 10'h1f8 == r_count_2_io_out ? io_r_504_b : _GEN_2093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2095 = 10'h1f9 == r_count_2_io_out ? io_r_505_b : _GEN_2094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2096 = 10'h1fa == r_count_2_io_out ? io_r_506_b : _GEN_2095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2097 = 10'h1fb == r_count_2_io_out ? io_r_507_b : _GEN_2096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2098 = 10'h1fc == r_count_2_io_out ? io_r_508_b : _GEN_2097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2099 = 10'h1fd == r_count_2_io_out ? io_r_509_b : _GEN_2098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2100 = 10'h1fe == r_count_2_io_out ? io_r_510_b : _GEN_2099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2101 = 10'h1ff == r_count_2_io_out ? io_r_511_b : _GEN_2100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2102 = 10'h200 == r_count_2_io_out ? io_r_512_b : _GEN_2101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2103 = 10'h201 == r_count_2_io_out ? io_r_513_b : _GEN_2102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2104 = 10'h202 == r_count_2_io_out ? io_r_514_b : _GEN_2103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2105 = 10'h203 == r_count_2_io_out ? io_r_515_b : _GEN_2104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2106 = 10'h204 == r_count_2_io_out ? io_r_516_b : _GEN_2105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2107 = 10'h205 == r_count_2_io_out ? io_r_517_b : _GEN_2106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2108 = 10'h206 == r_count_2_io_out ? io_r_518_b : _GEN_2107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2109 = 10'h207 == r_count_2_io_out ? io_r_519_b : _GEN_2108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2110 = 10'h208 == r_count_2_io_out ? io_r_520_b : _GEN_2109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2111 = 10'h209 == r_count_2_io_out ? io_r_521_b : _GEN_2110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2112 = 10'h20a == r_count_2_io_out ? io_r_522_b : _GEN_2111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2113 = 10'h20b == r_count_2_io_out ? io_r_523_b : _GEN_2112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2114 = 10'h20c == r_count_2_io_out ? io_r_524_b : _GEN_2113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2115 = 10'h20d == r_count_2_io_out ? io_r_525_b : _GEN_2114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2116 = 10'h20e == r_count_2_io_out ? io_r_526_b : _GEN_2115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2117 = 10'h20f == r_count_2_io_out ? io_r_527_b : _GEN_2116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2118 = 10'h210 == r_count_2_io_out ? io_r_528_b : _GEN_2117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2119 = 10'h211 == r_count_2_io_out ? io_r_529_b : _GEN_2118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2120 = 10'h212 == r_count_2_io_out ? io_r_530_b : _GEN_2119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2121 = 10'h213 == r_count_2_io_out ? io_r_531_b : _GEN_2120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2122 = 10'h214 == r_count_2_io_out ? io_r_532_b : _GEN_2121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2123 = 10'h215 == r_count_2_io_out ? io_r_533_b : _GEN_2122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2124 = 10'h216 == r_count_2_io_out ? io_r_534_b : _GEN_2123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2125 = 10'h217 == r_count_2_io_out ? io_r_535_b : _GEN_2124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2126 = 10'h218 == r_count_2_io_out ? io_r_536_b : _GEN_2125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2127 = 10'h219 == r_count_2_io_out ? io_r_537_b : _GEN_2126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2128 = 10'h21a == r_count_2_io_out ? io_r_538_b : _GEN_2127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2129 = 10'h21b == r_count_2_io_out ? io_r_539_b : _GEN_2128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2130 = 10'h21c == r_count_2_io_out ? io_r_540_b : _GEN_2129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2131 = 10'h21d == r_count_2_io_out ? io_r_541_b : _GEN_2130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2132 = 10'h21e == r_count_2_io_out ? io_r_542_b : _GEN_2131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2133 = 10'h21f == r_count_2_io_out ? io_r_543_b : _GEN_2132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2134 = 10'h220 == r_count_2_io_out ? io_r_544_b : _GEN_2133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2135 = 10'h221 == r_count_2_io_out ? io_r_545_b : _GEN_2134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2136 = 10'h222 == r_count_2_io_out ? io_r_546_b : _GEN_2135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2137 = 10'h223 == r_count_2_io_out ? io_r_547_b : _GEN_2136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2138 = 10'h224 == r_count_2_io_out ? io_r_548_b : _GEN_2137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2139 = 10'h225 == r_count_2_io_out ? io_r_549_b : _GEN_2138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2140 = 10'h226 == r_count_2_io_out ? io_r_550_b : _GEN_2139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2141 = 10'h227 == r_count_2_io_out ? io_r_551_b : _GEN_2140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2142 = 10'h228 == r_count_2_io_out ? io_r_552_b : _GEN_2141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2143 = 10'h229 == r_count_2_io_out ? io_r_553_b : _GEN_2142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2144 = 10'h22a == r_count_2_io_out ? io_r_554_b : _GEN_2143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2145 = 10'h22b == r_count_2_io_out ? io_r_555_b : _GEN_2144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2146 = 10'h22c == r_count_2_io_out ? io_r_556_b : _GEN_2145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2147 = 10'h22d == r_count_2_io_out ? io_r_557_b : _GEN_2146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2148 = 10'h22e == r_count_2_io_out ? io_r_558_b : _GEN_2147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2149 = 10'h22f == r_count_2_io_out ? io_r_559_b : _GEN_2148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2150 = 10'h230 == r_count_2_io_out ? io_r_560_b : _GEN_2149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2151 = 10'h231 == r_count_2_io_out ? io_r_561_b : _GEN_2150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2152 = 10'h232 == r_count_2_io_out ? io_r_562_b : _GEN_2151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2153 = 10'h233 == r_count_2_io_out ? io_r_563_b : _GEN_2152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2154 = 10'h234 == r_count_2_io_out ? io_r_564_b : _GEN_2153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2155 = 10'h235 == r_count_2_io_out ? io_r_565_b : _GEN_2154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2156 = 10'h236 == r_count_2_io_out ? io_r_566_b : _GEN_2155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2157 = 10'h237 == r_count_2_io_out ? io_r_567_b : _GEN_2156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2158 = 10'h238 == r_count_2_io_out ? io_r_568_b : _GEN_2157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2159 = 10'h239 == r_count_2_io_out ? io_r_569_b : _GEN_2158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2160 = 10'h23a == r_count_2_io_out ? io_r_570_b : _GEN_2159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2161 = 10'h23b == r_count_2_io_out ? io_r_571_b : _GEN_2160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2162 = 10'h23c == r_count_2_io_out ? io_r_572_b : _GEN_2161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2163 = 10'h23d == r_count_2_io_out ? io_r_573_b : _GEN_2162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2164 = 10'h23e == r_count_2_io_out ? io_r_574_b : _GEN_2163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2165 = 10'h23f == r_count_2_io_out ? io_r_575_b : _GEN_2164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2166 = 10'h240 == r_count_2_io_out ? io_r_576_b : _GEN_2165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2167 = 10'h241 == r_count_2_io_out ? io_r_577_b : _GEN_2166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2168 = 10'h242 == r_count_2_io_out ? io_r_578_b : _GEN_2167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2169 = 10'h243 == r_count_2_io_out ? io_r_579_b : _GEN_2168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2170 = 10'h244 == r_count_2_io_out ? io_r_580_b : _GEN_2169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2171 = 10'h245 == r_count_2_io_out ? io_r_581_b : _GEN_2170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2172 = 10'h246 == r_count_2_io_out ? io_r_582_b : _GEN_2171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2173 = 10'h247 == r_count_2_io_out ? io_r_583_b : _GEN_2172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2174 = 10'h248 == r_count_2_io_out ? io_r_584_b : _GEN_2173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2175 = 10'h249 == r_count_2_io_out ? io_r_585_b : _GEN_2174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2176 = 10'h24a == r_count_2_io_out ? io_r_586_b : _GEN_2175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2177 = 10'h24b == r_count_2_io_out ? io_r_587_b : _GEN_2176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2178 = 10'h24c == r_count_2_io_out ? io_r_588_b : _GEN_2177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2179 = 10'h24d == r_count_2_io_out ? io_r_589_b : _GEN_2178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2180 = 10'h24e == r_count_2_io_out ? io_r_590_b : _GEN_2179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2181 = 10'h24f == r_count_2_io_out ? io_r_591_b : _GEN_2180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2182 = 10'h250 == r_count_2_io_out ? io_r_592_b : _GEN_2181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2183 = 10'h251 == r_count_2_io_out ? io_r_593_b : _GEN_2182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2184 = 10'h252 == r_count_2_io_out ? io_r_594_b : _GEN_2183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2185 = 10'h253 == r_count_2_io_out ? io_r_595_b : _GEN_2184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2186 = 10'h254 == r_count_2_io_out ? io_r_596_b : _GEN_2185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2187 = 10'h255 == r_count_2_io_out ? io_r_597_b : _GEN_2186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2188 = 10'h256 == r_count_2_io_out ? io_r_598_b : _GEN_2187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2189 = 10'h257 == r_count_2_io_out ? io_r_599_b : _GEN_2188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2190 = 10'h258 == r_count_2_io_out ? io_r_600_b : _GEN_2189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2191 = 10'h259 == r_count_2_io_out ? io_r_601_b : _GEN_2190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2192 = 10'h25a == r_count_2_io_out ? io_r_602_b : _GEN_2191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2193 = 10'h25b == r_count_2_io_out ? io_r_603_b : _GEN_2192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2194 = 10'h25c == r_count_2_io_out ? io_r_604_b : _GEN_2193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2195 = 10'h25d == r_count_2_io_out ? io_r_605_b : _GEN_2194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2196 = 10'h25e == r_count_2_io_out ? io_r_606_b : _GEN_2195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2197 = 10'h25f == r_count_2_io_out ? io_r_607_b : _GEN_2196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2198 = 10'h260 == r_count_2_io_out ? io_r_608_b : _GEN_2197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2199 = 10'h261 == r_count_2_io_out ? io_r_609_b : _GEN_2198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2200 = 10'h262 == r_count_2_io_out ? io_r_610_b : _GEN_2199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2201 = 10'h263 == r_count_2_io_out ? io_r_611_b : _GEN_2200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2202 = 10'h264 == r_count_2_io_out ? io_r_612_b : _GEN_2201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2203 = 10'h265 == r_count_2_io_out ? io_r_613_b : _GEN_2202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2204 = 10'h266 == r_count_2_io_out ? io_r_614_b : _GEN_2203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2205 = 10'h267 == r_count_2_io_out ? io_r_615_b : _GEN_2204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2206 = 10'h268 == r_count_2_io_out ? io_r_616_b : _GEN_2205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2207 = 10'h269 == r_count_2_io_out ? io_r_617_b : _GEN_2206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2208 = 10'h26a == r_count_2_io_out ? io_r_618_b : _GEN_2207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2209 = 10'h26b == r_count_2_io_out ? io_r_619_b : _GEN_2208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2210 = 10'h26c == r_count_2_io_out ? io_r_620_b : _GEN_2209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2211 = 10'h26d == r_count_2_io_out ? io_r_621_b : _GEN_2210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2212 = 10'h26e == r_count_2_io_out ? io_r_622_b : _GEN_2211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2213 = 10'h26f == r_count_2_io_out ? io_r_623_b : _GEN_2212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2214 = 10'h270 == r_count_2_io_out ? io_r_624_b : _GEN_2213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2215 = 10'h271 == r_count_2_io_out ? io_r_625_b : _GEN_2214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2216 = 10'h272 == r_count_2_io_out ? io_r_626_b : _GEN_2215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2217 = 10'h273 == r_count_2_io_out ? io_r_627_b : _GEN_2216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2218 = 10'h274 == r_count_2_io_out ? io_r_628_b : _GEN_2217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2219 = 10'h275 == r_count_2_io_out ? io_r_629_b : _GEN_2218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2220 = 10'h276 == r_count_2_io_out ? io_r_630_b : _GEN_2219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2221 = 10'h277 == r_count_2_io_out ? io_r_631_b : _GEN_2220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2222 = 10'h278 == r_count_2_io_out ? io_r_632_b : _GEN_2221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2223 = 10'h279 == r_count_2_io_out ? io_r_633_b : _GEN_2222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2224 = 10'h27a == r_count_2_io_out ? io_r_634_b : _GEN_2223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2225 = 10'h27b == r_count_2_io_out ? io_r_635_b : _GEN_2224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2226 = 10'h27c == r_count_2_io_out ? io_r_636_b : _GEN_2225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2227 = 10'h27d == r_count_2_io_out ? io_r_637_b : _GEN_2226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2228 = 10'h27e == r_count_2_io_out ? io_r_638_b : _GEN_2227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2229 = 10'h27f == r_count_2_io_out ? io_r_639_b : _GEN_2228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2230 = 10'h280 == r_count_2_io_out ? io_r_640_b : _GEN_2229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2231 = 10'h281 == r_count_2_io_out ? io_r_641_b : _GEN_2230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2232 = 10'h282 == r_count_2_io_out ? io_r_642_b : _GEN_2231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2233 = 10'h283 == r_count_2_io_out ? io_r_643_b : _GEN_2232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2234 = 10'h284 == r_count_2_io_out ? io_r_644_b : _GEN_2233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2235 = 10'h285 == r_count_2_io_out ? io_r_645_b : _GEN_2234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2236 = 10'h286 == r_count_2_io_out ? io_r_646_b : _GEN_2235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2237 = 10'h287 == r_count_2_io_out ? io_r_647_b : _GEN_2236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2238 = 10'h288 == r_count_2_io_out ? io_r_648_b : _GEN_2237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2239 = 10'h289 == r_count_2_io_out ? io_r_649_b : _GEN_2238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2240 = 10'h28a == r_count_2_io_out ? io_r_650_b : _GEN_2239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2241 = 10'h28b == r_count_2_io_out ? io_r_651_b : _GEN_2240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2242 = 10'h28c == r_count_2_io_out ? io_r_652_b : _GEN_2241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2243 = 10'h28d == r_count_2_io_out ? io_r_653_b : _GEN_2242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2244 = 10'h28e == r_count_2_io_out ? io_r_654_b : _GEN_2243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2245 = 10'h28f == r_count_2_io_out ? io_r_655_b : _GEN_2244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2246 = 10'h290 == r_count_2_io_out ? io_r_656_b : _GEN_2245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2247 = 10'h291 == r_count_2_io_out ? io_r_657_b : _GEN_2246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2248 = 10'h292 == r_count_2_io_out ? io_r_658_b : _GEN_2247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2249 = 10'h293 == r_count_2_io_out ? io_r_659_b : _GEN_2248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2250 = 10'h294 == r_count_2_io_out ? io_r_660_b : _GEN_2249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2251 = 10'h295 == r_count_2_io_out ? io_r_661_b : _GEN_2250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2252 = 10'h296 == r_count_2_io_out ? io_r_662_b : _GEN_2251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2253 = 10'h297 == r_count_2_io_out ? io_r_663_b : _GEN_2252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2254 = 10'h298 == r_count_2_io_out ? io_r_664_b : _GEN_2253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2255 = 10'h299 == r_count_2_io_out ? io_r_665_b : _GEN_2254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2256 = 10'h29a == r_count_2_io_out ? io_r_666_b : _GEN_2255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2257 = 10'h29b == r_count_2_io_out ? io_r_667_b : _GEN_2256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2258 = 10'h29c == r_count_2_io_out ? io_r_668_b : _GEN_2257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2259 = 10'h29d == r_count_2_io_out ? io_r_669_b : _GEN_2258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2260 = 10'h29e == r_count_2_io_out ? io_r_670_b : _GEN_2259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2261 = 10'h29f == r_count_2_io_out ? io_r_671_b : _GEN_2260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2262 = 10'h2a0 == r_count_2_io_out ? io_r_672_b : _GEN_2261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2263 = 10'h2a1 == r_count_2_io_out ? io_r_673_b : _GEN_2262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2264 = 10'h2a2 == r_count_2_io_out ? io_r_674_b : _GEN_2263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2265 = 10'h2a3 == r_count_2_io_out ? io_r_675_b : _GEN_2264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2266 = 10'h2a4 == r_count_2_io_out ? io_r_676_b : _GEN_2265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2267 = 10'h2a5 == r_count_2_io_out ? io_r_677_b : _GEN_2266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2268 = 10'h2a6 == r_count_2_io_out ? io_r_678_b : _GEN_2267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2269 = 10'h2a7 == r_count_2_io_out ? io_r_679_b : _GEN_2268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2270 = 10'h2a8 == r_count_2_io_out ? io_r_680_b : _GEN_2269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2271 = 10'h2a9 == r_count_2_io_out ? io_r_681_b : _GEN_2270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2272 = 10'h2aa == r_count_2_io_out ? io_r_682_b : _GEN_2271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2273 = 10'h2ab == r_count_2_io_out ? io_r_683_b : _GEN_2272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2274 = 10'h2ac == r_count_2_io_out ? io_r_684_b : _GEN_2273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2275 = 10'h2ad == r_count_2_io_out ? io_r_685_b : _GEN_2274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2276 = 10'h2ae == r_count_2_io_out ? io_r_686_b : _GEN_2275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2277 = 10'h2af == r_count_2_io_out ? io_r_687_b : _GEN_2276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2278 = 10'h2b0 == r_count_2_io_out ? io_r_688_b : _GEN_2277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2279 = 10'h2b1 == r_count_2_io_out ? io_r_689_b : _GEN_2278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2280 = 10'h2b2 == r_count_2_io_out ? io_r_690_b : _GEN_2279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2281 = 10'h2b3 == r_count_2_io_out ? io_r_691_b : _GEN_2280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2282 = 10'h2b4 == r_count_2_io_out ? io_r_692_b : _GEN_2281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2283 = 10'h2b5 == r_count_2_io_out ? io_r_693_b : _GEN_2282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2284 = 10'h2b6 == r_count_2_io_out ? io_r_694_b : _GEN_2283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2285 = 10'h2b7 == r_count_2_io_out ? io_r_695_b : _GEN_2284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2286 = 10'h2b8 == r_count_2_io_out ? io_r_696_b : _GEN_2285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2287 = 10'h2b9 == r_count_2_io_out ? io_r_697_b : _GEN_2286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2288 = 10'h2ba == r_count_2_io_out ? io_r_698_b : _GEN_2287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2289 = 10'h2bb == r_count_2_io_out ? io_r_699_b : _GEN_2288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2290 = 10'h2bc == r_count_2_io_out ? io_r_700_b : _GEN_2289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2291 = 10'h2bd == r_count_2_io_out ? io_r_701_b : _GEN_2290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2292 = 10'h2be == r_count_2_io_out ? io_r_702_b : _GEN_2291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2293 = 10'h2bf == r_count_2_io_out ? io_r_703_b : _GEN_2292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2294 = 10'h2c0 == r_count_2_io_out ? io_r_704_b : _GEN_2293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2295 = 10'h2c1 == r_count_2_io_out ? io_r_705_b : _GEN_2294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2296 = 10'h2c2 == r_count_2_io_out ? io_r_706_b : _GEN_2295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2297 = 10'h2c3 == r_count_2_io_out ? io_r_707_b : _GEN_2296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2298 = 10'h2c4 == r_count_2_io_out ? io_r_708_b : _GEN_2297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2299 = 10'h2c5 == r_count_2_io_out ? io_r_709_b : _GEN_2298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2300 = 10'h2c6 == r_count_2_io_out ? io_r_710_b : _GEN_2299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2301 = 10'h2c7 == r_count_2_io_out ? io_r_711_b : _GEN_2300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2302 = 10'h2c8 == r_count_2_io_out ? io_r_712_b : _GEN_2301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2303 = 10'h2c9 == r_count_2_io_out ? io_r_713_b : _GEN_2302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2304 = 10'h2ca == r_count_2_io_out ? io_r_714_b : _GEN_2303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2305 = 10'h2cb == r_count_2_io_out ? io_r_715_b : _GEN_2304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2306 = 10'h2cc == r_count_2_io_out ? io_r_716_b : _GEN_2305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2307 = 10'h2cd == r_count_2_io_out ? io_r_717_b : _GEN_2306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2308 = 10'h2ce == r_count_2_io_out ? io_r_718_b : _GEN_2307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2309 = 10'h2cf == r_count_2_io_out ? io_r_719_b : _GEN_2308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2310 = 10'h2d0 == r_count_2_io_out ? io_r_720_b : _GEN_2309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2311 = 10'h2d1 == r_count_2_io_out ? io_r_721_b : _GEN_2310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2312 = 10'h2d2 == r_count_2_io_out ? io_r_722_b : _GEN_2311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2313 = 10'h2d3 == r_count_2_io_out ? io_r_723_b : _GEN_2312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2314 = 10'h2d4 == r_count_2_io_out ? io_r_724_b : _GEN_2313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2315 = 10'h2d5 == r_count_2_io_out ? io_r_725_b : _GEN_2314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2316 = 10'h2d6 == r_count_2_io_out ? io_r_726_b : _GEN_2315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2317 = 10'h2d7 == r_count_2_io_out ? io_r_727_b : _GEN_2316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2318 = 10'h2d8 == r_count_2_io_out ? io_r_728_b : _GEN_2317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2319 = 10'h2d9 == r_count_2_io_out ? io_r_729_b : _GEN_2318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2320 = 10'h2da == r_count_2_io_out ? io_r_730_b : _GEN_2319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2321 = 10'h2db == r_count_2_io_out ? io_r_731_b : _GEN_2320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2322 = 10'h2dc == r_count_2_io_out ? io_r_732_b : _GEN_2321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2323 = 10'h2dd == r_count_2_io_out ? io_r_733_b : _GEN_2322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2324 = 10'h2de == r_count_2_io_out ? io_r_734_b : _GEN_2323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2325 = 10'h2df == r_count_2_io_out ? io_r_735_b : _GEN_2324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2326 = 10'h2e0 == r_count_2_io_out ? io_r_736_b : _GEN_2325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2327 = 10'h2e1 == r_count_2_io_out ? io_r_737_b : _GEN_2326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2328 = 10'h2e2 == r_count_2_io_out ? io_r_738_b : _GEN_2327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2329 = 10'h2e3 == r_count_2_io_out ? io_r_739_b : _GEN_2328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2330 = 10'h2e4 == r_count_2_io_out ? io_r_740_b : _GEN_2329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2331 = 10'h2e5 == r_count_2_io_out ? io_r_741_b : _GEN_2330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2332 = 10'h2e6 == r_count_2_io_out ? io_r_742_b : _GEN_2331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2333 = 10'h2e7 == r_count_2_io_out ? io_r_743_b : _GEN_2332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2334 = 10'h2e8 == r_count_2_io_out ? io_r_744_b : _GEN_2333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2335 = 10'h2e9 == r_count_2_io_out ? io_r_745_b : _GEN_2334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2336 = 10'h2ea == r_count_2_io_out ? io_r_746_b : _GEN_2335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2337 = 10'h2eb == r_count_2_io_out ? io_r_747_b : _GEN_2336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2338 = 10'h2ec == r_count_2_io_out ? io_r_748_b : _GEN_2337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2341 = 10'h1 == r_count_3_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2342 = 10'h2 == r_count_3_io_out ? io_r_2_b : _GEN_2341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2343 = 10'h3 == r_count_3_io_out ? io_r_3_b : _GEN_2342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2344 = 10'h4 == r_count_3_io_out ? io_r_4_b : _GEN_2343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2345 = 10'h5 == r_count_3_io_out ? io_r_5_b : _GEN_2344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2346 = 10'h6 == r_count_3_io_out ? io_r_6_b : _GEN_2345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2347 = 10'h7 == r_count_3_io_out ? io_r_7_b : _GEN_2346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2348 = 10'h8 == r_count_3_io_out ? io_r_8_b : _GEN_2347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2349 = 10'h9 == r_count_3_io_out ? io_r_9_b : _GEN_2348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2350 = 10'ha == r_count_3_io_out ? io_r_10_b : _GEN_2349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2351 = 10'hb == r_count_3_io_out ? io_r_11_b : _GEN_2350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2352 = 10'hc == r_count_3_io_out ? io_r_12_b : _GEN_2351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2353 = 10'hd == r_count_3_io_out ? io_r_13_b : _GEN_2352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2354 = 10'he == r_count_3_io_out ? io_r_14_b : _GEN_2353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2355 = 10'hf == r_count_3_io_out ? io_r_15_b : _GEN_2354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2356 = 10'h10 == r_count_3_io_out ? io_r_16_b : _GEN_2355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2357 = 10'h11 == r_count_3_io_out ? io_r_17_b : _GEN_2356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2358 = 10'h12 == r_count_3_io_out ? io_r_18_b : _GEN_2357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2359 = 10'h13 == r_count_3_io_out ? io_r_19_b : _GEN_2358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2360 = 10'h14 == r_count_3_io_out ? io_r_20_b : _GEN_2359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2361 = 10'h15 == r_count_3_io_out ? io_r_21_b : _GEN_2360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2362 = 10'h16 == r_count_3_io_out ? io_r_22_b : _GEN_2361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2363 = 10'h17 == r_count_3_io_out ? io_r_23_b : _GEN_2362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2364 = 10'h18 == r_count_3_io_out ? io_r_24_b : _GEN_2363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2365 = 10'h19 == r_count_3_io_out ? io_r_25_b : _GEN_2364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2366 = 10'h1a == r_count_3_io_out ? io_r_26_b : _GEN_2365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2367 = 10'h1b == r_count_3_io_out ? io_r_27_b : _GEN_2366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2368 = 10'h1c == r_count_3_io_out ? io_r_28_b : _GEN_2367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2369 = 10'h1d == r_count_3_io_out ? io_r_29_b : _GEN_2368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2370 = 10'h1e == r_count_3_io_out ? io_r_30_b : _GEN_2369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2371 = 10'h1f == r_count_3_io_out ? io_r_31_b : _GEN_2370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2372 = 10'h20 == r_count_3_io_out ? io_r_32_b : _GEN_2371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2373 = 10'h21 == r_count_3_io_out ? io_r_33_b : _GEN_2372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2374 = 10'h22 == r_count_3_io_out ? io_r_34_b : _GEN_2373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2375 = 10'h23 == r_count_3_io_out ? io_r_35_b : _GEN_2374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2376 = 10'h24 == r_count_3_io_out ? io_r_36_b : _GEN_2375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2377 = 10'h25 == r_count_3_io_out ? io_r_37_b : _GEN_2376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2378 = 10'h26 == r_count_3_io_out ? io_r_38_b : _GEN_2377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2379 = 10'h27 == r_count_3_io_out ? io_r_39_b : _GEN_2378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2380 = 10'h28 == r_count_3_io_out ? io_r_40_b : _GEN_2379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2381 = 10'h29 == r_count_3_io_out ? io_r_41_b : _GEN_2380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2382 = 10'h2a == r_count_3_io_out ? io_r_42_b : _GEN_2381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2383 = 10'h2b == r_count_3_io_out ? io_r_43_b : _GEN_2382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2384 = 10'h2c == r_count_3_io_out ? io_r_44_b : _GEN_2383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2385 = 10'h2d == r_count_3_io_out ? io_r_45_b : _GEN_2384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2386 = 10'h2e == r_count_3_io_out ? io_r_46_b : _GEN_2385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2387 = 10'h2f == r_count_3_io_out ? io_r_47_b : _GEN_2386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2388 = 10'h30 == r_count_3_io_out ? io_r_48_b : _GEN_2387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2389 = 10'h31 == r_count_3_io_out ? io_r_49_b : _GEN_2388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2390 = 10'h32 == r_count_3_io_out ? io_r_50_b : _GEN_2389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2391 = 10'h33 == r_count_3_io_out ? io_r_51_b : _GEN_2390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2392 = 10'h34 == r_count_3_io_out ? io_r_52_b : _GEN_2391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2393 = 10'h35 == r_count_3_io_out ? io_r_53_b : _GEN_2392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2394 = 10'h36 == r_count_3_io_out ? io_r_54_b : _GEN_2393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2395 = 10'h37 == r_count_3_io_out ? io_r_55_b : _GEN_2394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2396 = 10'h38 == r_count_3_io_out ? io_r_56_b : _GEN_2395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2397 = 10'h39 == r_count_3_io_out ? io_r_57_b : _GEN_2396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2398 = 10'h3a == r_count_3_io_out ? io_r_58_b : _GEN_2397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2399 = 10'h3b == r_count_3_io_out ? io_r_59_b : _GEN_2398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2400 = 10'h3c == r_count_3_io_out ? io_r_60_b : _GEN_2399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2401 = 10'h3d == r_count_3_io_out ? io_r_61_b : _GEN_2400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2402 = 10'h3e == r_count_3_io_out ? io_r_62_b : _GEN_2401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2403 = 10'h3f == r_count_3_io_out ? io_r_63_b : _GEN_2402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2404 = 10'h40 == r_count_3_io_out ? io_r_64_b : _GEN_2403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2405 = 10'h41 == r_count_3_io_out ? io_r_65_b : _GEN_2404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2406 = 10'h42 == r_count_3_io_out ? io_r_66_b : _GEN_2405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2407 = 10'h43 == r_count_3_io_out ? io_r_67_b : _GEN_2406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2408 = 10'h44 == r_count_3_io_out ? io_r_68_b : _GEN_2407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2409 = 10'h45 == r_count_3_io_out ? io_r_69_b : _GEN_2408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2410 = 10'h46 == r_count_3_io_out ? io_r_70_b : _GEN_2409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2411 = 10'h47 == r_count_3_io_out ? io_r_71_b : _GEN_2410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2412 = 10'h48 == r_count_3_io_out ? io_r_72_b : _GEN_2411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2413 = 10'h49 == r_count_3_io_out ? io_r_73_b : _GEN_2412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2414 = 10'h4a == r_count_3_io_out ? io_r_74_b : _GEN_2413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2415 = 10'h4b == r_count_3_io_out ? io_r_75_b : _GEN_2414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2416 = 10'h4c == r_count_3_io_out ? io_r_76_b : _GEN_2415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2417 = 10'h4d == r_count_3_io_out ? io_r_77_b : _GEN_2416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2418 = 10'h4e == r_count_3_io_out ? io_r_78_b : _GEN_2417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2419 = 10'h4f == r_count_3_io_out ? io_r_79_b : _GEN_2418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2420 = 10'h50 == r_count_3_io_out ? io_r_80_b : _GEN_2419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2421 = 10'h51 == r_count_3_io_out ? io_r_81_b : _GEN_2420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2422 = 10'h52 == r_count_3_io_out ? io_r_82_b : _GEN_2421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2423 = 10'h53 == r_count_3_io_out ? io_r_83_b : _GEN_2422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2424 = 10'h54 == r_count_3_io_out ? io_r_84_b : _GEN_2423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2425 = 10'h55 == r_count_3_io_out ? io_r_85_b : _GEN_2424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2426 = 10'h56 == r_count_3_io_out ? io_r_86_b : _GEN_2425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2427 = 10'h57 == r_count_3_io_out ? io_r_87_b : _GEN_2426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2428 = 10'h58 == r_count_3_io_out ? io_r_88_b : _GEN_2427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2429 = 10'h59 == r_count_3_io_out ? io_r_89_b : _GEN_2428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2430 = 10'h5a == r_count_3_io_out ? io_r_90_b : _GEN_2429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2431 = 10'h5b == r_count_3_io_out ? io_r_91_b : _GEN_2430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2432 = 10'h5c == r_count_3_io_out ? io_r_92_b : _GEN_2431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2433 = 10'h5d == r_count_3_io_out ? io_r_93_b : _GEN_2432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2434 = 10'h5e == r_count_3_io_out ? io_r_94_b : _GEN_2433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2435 = 10'h5f == r_count_3_io_out ? io_r_95_b : _GEN_2434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2436 = 10'h60 == r_count_3_io_out ? io_r_96_b : _GEN_2435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2437 = 10'h61 == r_count_3_io_out ? io_r_97_b : _GEN_2436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2438 = 10'h62 == r_count_3_io_out ? io_r_98_b : _GEN_2437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2439 = 10'h63 == r_count_3_io_out ? io_r_99_b : _GEN_2438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2440 = 10'h64 == r_count_3_io_out ? io_r_100_b : _GEN_2439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2441 = 10'h65 == r_count_3_io_out ? io_r_101_b : _GEN_2440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2442 = 10'h66 == r_count_3_io_out ? io_r_102_b : _GEN_2441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2443 = 10'h67 == r_count_3_io_out ? io_r_103_b : _GEN_2442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2444 = 10'h68 == r_count_3_io_out ? io_r_104_b : _GEN_2443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2445 = 10'h69 == r_count_3_io_out ? io_r_105_b : _GEN_2444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2446 = 10'h6a == r_count_3_io_out ? io_r_106_b : _GEN_2445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2447 = 10'h6b == r_count_3_io_out ? io_r_107_b : _GEN_2446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2448 = 10'h6c == r_count_3_io_out ? io_r_108_b : _GEN_2447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2449 = 10'h6d == r_count_3_io_out ? io_r_109_b : _GEN_2448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2450 = 10'h6e == r_count_3_io_out ? io_r_110_b : _GEN_2449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2451 = 10'h6f == r_count_3_io_out ? io_r_111_b : _GEN_2450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2452 = 10'h70 == r_count_3_io_out ? io_r_112_b : _GEN_2451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2453 = 10'h71 == r_count_3_io_out ? io_r_113_b : _GEN_2452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2454 = 10'h72 == r_count_3_io_out ? io_r_114_b : _GEN_2453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2455 = 10'h73 == r_count_3_io_out ? io_r_115_b : _GEN_2454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2456 = 10'h74 == r_count_3_io_out ? io_r_116_b : _GEN_2455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2457 = 10'h75 == r_count_3_io_out ? io_r_117_b : _GEN_2456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2458 = 10'h76 == r_count_3_io_out ? io_r_118_b : _GEN_2457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2459 = 10'h77 == r_count_3_io_out ? io_r_119_b : _GEN_2458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2460 = 10'h78 == r_count_3_io_out ? io_r_120_b : _GEN_2459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2461 = 10'h79 == r_count_3_io_out ? io_r_121_b : _GEN_2460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2462 = 10'h7a == r_count_3_io_out ? io_r_122_b : _GEN_2461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2463 = 10'h7b == r_count_3_io_out ? io_r_123_b : _GEN_2462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2464 = 10'h7c == r_count_3_io_out ? io_r_124_b : _GEN_2463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2465 = 10'h7d == r_count_3_io_out ? io_r_125_b : _GEN_2464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2466 = 10'h7e == r_count_3_io_out ? io_r_126_b : _GEN_2465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2467 = 10'h7f == r_count_3_io_out ? io_r_127_b : _GEN_2466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2468 = 10'h80 == r_count_3_io_out ? io_r_128_b : _GEN_2467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2469 = 10'h81 == r_count_3_io_out ? io_r_129_b : _GEN_2468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2470 = 10'h82 == r_count_3_io_out ? io_r_130_b : _GEN_2469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2471 = 10'h83 == r_count_3_io_out ? io_r_131_b : _GEN_2470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2472 = 10'h84 == r_count_3_io_out ? io_r_132_b : _GEN_2471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2473 = 10'h85 == r_count_3_io_out ? io_r_133_b : _GEN_2472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2474 = 10'h86 == r_count_3_io_out ? io_r_134_b : _GEN_2473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2475 = 10'h87 == r_count_3_io_out ? io_r_135_b : _GEN_2474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2476 = 10'h88 == r_count_3_io_out ? io_r_136_b : _GEN_2475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2477 = 10'h89 == r_count_3_io_out ? io_r_137_b : _GEN_2476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2478 = 10'h8a == r_count_3_io_out ? io_r_138_b : _GEN_2477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2479 = 10'h8b == r_count_3_io_out ? io_r_139_b : _GEN_2478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2480 = 10'h8c == r_count_3_io_out ? io_r_140_b : _GEN_2479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2481 = 10'h8d == r_count_3_io_out ? io_r_141_b : _GEN_2480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2482 = 10'h8e == r_count_3_io_out ? io_r_142_b : _GEN_2481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2483 = 10'h8f == r_count_3_io_out ? io_r_143_b : _GEN_2482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2484 = 10'h90 == r_count_3_io_out ? io_r_144_b : _GEN_2483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2485 = 10'h91 == r_count_3_io_out ? io_r_145_b : _GEN_2484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2486 = 10'h92 == r_count_3_io_out ? io_r_146_b : _GEN_2485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2487 = 10'h93 == r_count_3_io_out ? io_r_147_b : _GEN_2486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2488 = 10'h94 == r_count_3_io_out ? io_r_148_b : _GEN_2487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2489 = 10'h95 == r_count_3_io_out ? io_r_149_b : _GEN_2488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2490 = 10'h96 == r_count_3_io_out ? io_r_150_b : _GEN_2489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2491 = 10'h97 == r_count_3_io_out ? io_r_151_b : _GEN_2490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2492 = 10'h98 == r_count_3_io_out ? io_r_152_b : _GEN_2491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2493 = 10'h99 == r_count_3_io_out ? io_r_153_b : _GEN_2492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2494 = 10'h9a == r_count_3_io_out ? io_r_154_b : _GEN_2493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2495 = 10'h9b == r_count_3_io_out ? io_r_155_b : _GEN_2494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2496 = 10'h9c == r_count_3_io_out ? io_r_156_b : _GEN_2495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2497 = 10'h9d == r_count_3_io_out ? io_r_157_b : _GEN_2496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2498 = 10'h9e == r_count_3_io_out ? io_r_158_b : _GEN_2497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2499 = 10'h9f == r_count_3_io_out ? io_r_159_b : _GEN_2498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2500 = 10'ha0 == r_count_3_io_out ? io_r_160_b : _GEN_2499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2501 = 10'ha1 == r_count_3_io_out ? io_r_161_b : _GEN_2500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2502 = 10'ha2 == r_count_3_io_out ? io_r_162_b : _GEN_2501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2503 = 10'ha3 == r_count_3_io_out ? io_r_163_b : _GEN_2502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2504 = 10'ha4 == r_count_3_io_out ? io_r_164_b : _GEN_2503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2505 = 10'ha5 == r_count_3_io_out ? io_r_165_b : _GEN_2504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2506 = 10'ha6 == r_count_3_io_out ? io_r_166_b : _GEN_2505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2507 = 10'ha7 == r_count_3_io_out ? io_r_167_b : _GEN_2506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2508 = 10'ha8 == r_count_3_io_out ? io_r_168_b : _GEN_2507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2509 = 10'ha9 == r_count_3_io_out ? io_r_169_b : _GEN_2508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2510 = 10'haa == r_count_3_io_out ? io_r_170_b : _GEN_2509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2511 = 10'hab == r_count_3_io_out ? io_r_171_b : _GEN_2510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2512 = 10'hac == r_count_3_io_out ? io_r_172_b : _GEN_2511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2513 = 10'had == r_count_3_io_out ? io_r_173_b : _GEN_2512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2514 = 10'hae == r_count_3_io_out ? io_r_174_b : _GEN_2513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2515 = 10'haf == r_count_3_io_out ? io_r_175_b : _GEN_2514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2516 = 10'hb0 == r_count_3_io_out ? io_r_176_b : _GEN_2515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2517 = 10'hb1 == r_count_3_io_out ? io_r_177_b : _GEN_2516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2518 = 10'hb2 == r_count_3_io_out ? io_r_178_b : _GEN_2517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2519 = 10'hb3 == r_count_3_io_out ? io_r_179_b : _GEN_2518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2520 = 10'hb4 == r_count_3_io_out ? io_r_180_b : _GEN_2519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2521 = 10'hb5 == r_count_3_io_out ? io_r_181_b : _GEN_2520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2522 = 10'hb6 == r_count_3_io_out ? io_r_182_b : _GEN_2521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2523 = 10'hb7 == r_count_3_io_out ? io_r_183_b : _GEN_2522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2524 = 10'hb8 == r_count_3_io_out ? io_r_184_b : _GEN_2523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2525 = 10'hb9 == r_count_3_io_out ? io_r_185_b : _GEN_2524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2526 = 10'hba == r_count_3_io_out ? io_r_186_b : _GEN_2525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2527 = 10'hbb == r_count_3_io_out ? io_r_187_b : _GEN_2526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2528 = 10'hbc == r_count_3_io_out ? io_r_188_b : _GEN_2527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2529 = 10'hbd == r_count_3_io_out ? io_r_189_b : _GEN_2528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2530 = 10'hbe == r_count_3_io_out ? io_r_190_b : _GEN_2529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2531 = 10'hbf == r_count_3_io_out ? io_r_191_b : _GEN_2530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2532 = 10'hc0 == r_count_3_io_out ? io_r_192_b : _GEN_2531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2533 = 10'hc1 == r_count_3_io_out ? io_r_193_b : _GEN_2532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2534 = 10'hc2 == r_count_3_io_out ? io_r_194_b : _GEN_2533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2535 = 10'hc3 == r_count_3_io_out ? io_r_195_b : _GEN_2534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2536 = 10'hc4 == r_count_3_io_out ? io_r_196_b : _GEN_2535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2537 = 10'hc5 == r_count_3_io_out ? io_r_197_b : _GEN_2536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2538 = 10'hc6 == r_count_3_io_out ? io_r_198_b : _GEN_2537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2539 = 10'hc7 == r_count_3_io_out ? io_r_199_b : _GEN_2538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2540 = 10'hc8 == r_count_3_io_out ? io_r_200_b : _GEN_2539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2541 = 10'hc9 == r_count_3_io_out ? io_r_201_b : _GEN_2540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2542 = 10'hca == r_count_3_io_out ? io_r_202_b : _GEN_2541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2543 = 10'hcb == r_count_3_io_out ? io_r_203_b : _GEN_2542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2544 = 10'hcc == r_count_3_io_out ? io_r_204_b : _GEN_2543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2545 = 10'hcd == r_count_3_io_out ? io_r_205_b : _GEN_2544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2546 = 10'hce == r_count_3_io_out ? io_r_206_b : _GEN_2545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2547 = 10'hcf == r_count_3_io_out ? io_r_207_b : _GEN_2546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2548 = 10'hd0 == r_count_3_io_out ? io_r_208_b : _GEN_2547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2549 = 10'hd1 == r_count_3_io_out ? io_r_209_b : _GEN_2548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2550 = 10'hd2 == r_count_3_io_out ? io_r_210_b : _GEN_2549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2551 = 10'hd3 == r_count_3_io_out ? io_r_211_b : _GEN_2550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2552 = 10'hd4 == r_count_3_io_out ? io_r_212_b : _GEN_2551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2553 = 10'hd5 == r_count_3_io_out ? io_r_213_b : _GEN_2552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2554 = 10'hd6 == r_count_3_io_out ? io_r_214_b : _GEN_2553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2555 = 10'hd7 == r_count_3_io_out ? io_r_215_b : _GEN_2554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2556 = 10'hd8 == r_count_3_io_out ? io_r_216_b : _GEN_2555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2557 = 10'hd9 == r_count_3_io_out ? io_r_217_b : _GEN_2556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2558 = 10'hda == r_count_3_io_out ? io_r_218_b : _GEN_2557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2559 = 10'hdb == r_count_3_io_out ? io_r_219_b : _GEN_2558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2560 = 10'hdc == r_count_3_io_out ? io_r_220_b : _GEN_2559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2561 = 10'hdd == r_count_3_io_out ? io_r_221_b : _GEN_2560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2562 = 10'hde == r_count_3_io_out ? io_r_222_b : _GEN_2561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2563 = 10'hdf == r_count_3_io_out ? io_r_223_b : _GEN_2562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2564 = 10'he0 == r_count_3_io_out ? io_r_224_b : _GEN_2563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2565 = 10'he1 == r_count_3_io_out ? io_r_225_b : _GEN_2564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2566 = 10'he2 == r_count_3_io_out ? io_r_226_b : _GEN_2565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2567 = 10'he3 == r_count_3_io_out ? io_r_227_b : _GEN_2566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2568 = 10'he4 == r_count_3_io_out ? io_r_228_b : _GEN_2567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2569 = 10'he5 == r_count_3_io_out ? io_r_229_b : _GEN_2568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2570 = 10'he6 == r_count_3_io_out ? io_r_230_b : _GEN_2569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2571 = 10'he7 == r_count_3_io_out ? io_r_231_b : _GEN_2570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2572 = 10'he8 == r_count_3_io_out ? io_r_232_b : _GEN_2571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2573 = 10'he9 == r_count_3_io_out ? io_r_233_b : _GEN_2572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2574 = 10'hea == r_count_3_io_out ? io_r_234_b : _GEN_2573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2575 = 10'heb == r_count_3_io_out ? io_r_235_b : _GEN_2574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2576 = 10'hec == r_count_3_io_out ? io_r_236_b : _GEN_2575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2577 = 10'hed == r_count_3_io_out ? io_r_237_b : _GEN_2576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2578 = 10'hee == r_count_3_io_out ? io_r_238_b : _GEN_2577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2579 = 10'hef == r_count_3_io_out ? io_r_239_b : _GEN_2578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2580 = 10'hf0 == r_count_3_io_out ? io_r_240_b : _GEN_2579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2581 = 10'hf1 == r_count_3_io_out ? io_r_241_b : _GEN_2580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2582 = 10'hf2 == r_count_3_io_out ? io_r_242_b : _GEN_2581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2583 = 10'hf3 == r_count_3_io_out ? io_r_243_b : _GEN_2582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2584 = 10'hf4 == r_count_3_io_out ? io_r_244_b : _GEN_2583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2585 = 10'hf5 == r_count_3_io_out ? io_r_245_b : _GEN_2584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2586 = 10'hf6 == r_count_3_io_out ? io_r_246_b : _GEN_2585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2587 = 10'hf7 == r_count_3_io_out ? io_r_247_b : _GEN_2586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2588 = 10'hf8 == r_count_3_io_out ? io_r_248_b : _GEN_2587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2589 = 10'hf9 == r_count_3_io_out ? io_r_249_b : _GEN_2588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2590 = 10'hfa == r_count_3_io_out ? io_r_250_b : _GEN_2589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2591 = 10'hfb == r_count_3_io_out ? io_r_251_b : _GEN_2590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2592 = 10'hfc == r_count_3_io_out ? io_r_252_b : _GEN_2591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2593 = 10'hfd == r_count_3_io_out ? io_r_253_b : _GEN_2592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2594 = 10'hfe == r_count_3_io_out ? io_r_254_b : _GEN_2593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2595 = 10'hff == r_count_3_io_out ? io_r_255_b : _GEN_2594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2596 = 10'h100 == r_count_3_io_out ? io_r_256_b : _GEN_2595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2597 = 10'h101 == r_count_3_io_out ? io_r_257_b : _GEN_2596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2598 = 10'h102 == r_count_3_io_out ? io_r_258_b : _GEN_2597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2599 = 10'h103 == r_count_3_io_out ? io_r_259_b : _GEN_2598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2600 = 10'h104 == r_count_3_io_out ? io_r_260_b : _GEN_2599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2601 = 10'h105 == r_count_3_io_out ? io_r_261_b : _GEN_2600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2602 = 10'h106 == r_count_3_io_out ? io_r_262_b : _GEN_2601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2603 = 10'h107 == r_count_3_io_out ? io_r_263_b : _GEN_2602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2604 = 10'h108 == r_count_3_io_out ? io_r_264_b : _GEN_2603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2605 = 10'h109 == r_count_3_io_out ? io_r_265_b : _GEN_2604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2606 = 10'h10a == r_count_3_io_out ? io_r_266_b : _GEN_2605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2607 = 10'h10b == r_count_3_io_out ? io_r_267_b : _GEN_2606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2608 = 10'h10c == r_count_3_io_out ? io_r_268_b : _GEN_2607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2609 = 10'h10d == r_count_3_io_out ? io_r_269_b : _GEN_2608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2610 = 10'h10e == r_count_3_io_out ? io_r_270_b : _GEN_2609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2611 = 10'h10f == r_count_3_io_out ? io_r_271_b : _GEN_2610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2612 = 10'h110 == r_count_3_io_out ? io_r_272_b : _GEN_2611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2613 = 10'h111 == r_count_3_io_out ? io_r_273_b : _GEN_2612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2614 = 10'h112 == r_count_3_io_out ? io_r_274_b : _GEN_2613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2615 = 10'h113 == r_count_3_io_out ? io_r_275_b : _GEN_2614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2616 = 10'h114 == r_count_3_io_out ? io_r_276_b : _GEN_2615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2617 = 10'h115 == r_count_3_io_out ? io_r_277_b : _GEN_2616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2618 = 10'h116 == r_count_3_io_out ? io_r_278_b : _GEN_2617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2619 = 10'h117 == r_count_3_io_out ? io_r_279_b : _GEN_2618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2620 = 10'h118 == r_count_3_io_out ? io_r_280_b : _GEN_2619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2621 = 10'h119 == r_count_3_io_out ? io_r_281_b : _GEN_2620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2622 = 10'h11a == r_count_3_io_out ? io_r_282_b : _GEN_2621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2623 = 10'h11b == r_count_3_io_out ? io_r_283_b : _GEN_2622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2624 = 10'h11c == r_count_3_io_out ? io_r_284_b : _GEN_2623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2625 = 10'h11d == r_count_3_io_out ? io_r_285_b : _GEN_2624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2626 = 10'h11e == r_count_3_io_out ? io_r_286_b : _GEN_2625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2627 = 10'h11f == r_count_3_io_out ? io_r_287_b : _GEN_2626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2628 = 10'h120 == r_count_3_io_out ? io_r_288_b : _GEN_2627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2629 = 10'h121 == r_count_3_io_out ? io_r_289_b : _GEN_2628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2630 = 10'h122 == r_count_3_io_out ? io_r_290_b : _GEN_2629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2631 = 10'h123 == r_count_3_io_out ? io_r_291_b : _GEN_2630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2632 = 10'h124 == r_count_3_io_out ? io_r_292_b : _GEN_2631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2633 = 10'h125 == r_count_3_io_out ? io_r_293_b : _GEN_2632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2634 = 10'h126 == r_count_3_io_out ? io_r_294_b : _GEN_2633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2635 = 10'h127 == r_count_3_io_out ? io_r_295_b : _GEN_2634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2636 = 10'h128 == r_count_3_io_out ? io_r_296_b : _GEN_2635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2637 = 10'h129 == r_count_3_io_out ? io_r_297_b : _GEN_2636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2638 = 10'h12a == r_count_3_io_out ? io_r_298_b : _GEN_2637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2639 = 10'h12b == r_count_3_io_out ? io_r_299_b : _GEN_2638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2640 = 10'h12c == r_count_3_io_out ? io_r_300_b : _GEN_2639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2641 = 10'h12d == r_count_3_io_out ? io_r_301_b : _GEN_2640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2642 = 10'h12e == r_count_3_io_out ? io_r_302_b : _GEN_2641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2643 = 10'h12f == r_count_3_io_out ? io_r_303_b : _GEN_2642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2644 = 10'h130 == r_count_3_io_out ? io_r_304_b : _GEN_2643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2645 = 10'h131 == r_count_3_io_out ? io_r_305_b : _GEN_2644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2646 = 10'h132 == r_count_3_io_out ? io_r_306_b : _GEN_2645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2647 = 10'h133 == r_count_3_io_out ? io_r_307_b : _GEN_2646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2648 = 10'h134 == r_count_3_io_out ? io_r_308_b : _GEN_2647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2649 = 10'h135 == r_count_3_io_out ? io_r_309_b : _GEN_2648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2650 = 10'h136 == r_count_3_io_out ? io_r_310_b : _GEN_2649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2651 = 10'h137 == r_count_3_io_out ? io_r_311_b : _GEN_2650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2652 = 10'h138 == r_count_3_io_out ? io_r_312_b : _GEN_2651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2653 = 10'h139 == r_count_3_io_out ? io_r_313_b : _GEN_2652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2654 = 10'h13a == r_count_3_io_out ? io_r_314_b : _GEN_2653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2655 = 10'h13b == r_count_3_io_out ? io_r_315_b : _GEN_2654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2656 = 10'h13c == r_count_3_io_out ? io_r_316_b : _GEN_2655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2657 = 10'h13d == r_count_3_io_out ? io_r_317_b : _GEN_2656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2658 = 10'h13e == r_count_3_io_out ? io_r_318_b : _GEN_2657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2659 = 10'h13f == r_count_3_io_out ? io_r_319_b : _GEN_2658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2660 = 10'h140 == r_count_3_io_out ? io_r_320_b : _GEN_2659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2661 = 10'h141 == r_count_3_io_out ? io_r_321_b : _GEN_2660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2662 = 10'h142 == r_count_3_io_out ? io_r_322_b : _GEN_2661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2663 = 10'h143 == r_count_3_io_out ? io_r_323_b : _GEN_2662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2664 = 10'h144 == r_count_3_io_out ? io_r_324_b : _GEN_2663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2665 = 10'h145 == r_count_3_io_out ? io_r_325_b : _GEN_2664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2666 = 10'h146 == r_count_3_io_out ? io_r_326_b : _GEN_2665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2667 = 10'h147 == r_count_3_io_out ? io_r_327_b : _GEN_2666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2668 = 10'h148 == r_count_3_io_out ? io_r_328_b : _GEN_2667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2669 = 10'h149 == r_count_3_io_out ? io_r_329_b : _GEN_2668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2670 = 10'h14a == r_count_3_io_out ? io_r_330_b : _GEN_2669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2671 = 10'h14b == r_count_3_io_out ? io_r_331_b : _GEN_2670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2672 = 10'h14c == r_count_3_io_out ? io_r_332_b : _GEN_2671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2673 = 10'h14d == r_count_3_io_out ? io_r_333_b : _GEN_2672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2674 = 10'h14e == r_count_3_io_out ? io_r_334_b : _GEN_2673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2675 = 10'h14f == r_count_3_io_out ? io_r_335_b : _GEN_2674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2676 = 10'h150 == r_count_3_io_out ? io_r_336_b : _GEN_2675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2677 = 10'h151 == r_count_3_io_out ? io_r_337_b : _GEN_2676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2678 = 10'h152 == r_count_3_io_out ? io_r_338_b : _GEN_2677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2679 = 10'h153 == r_count_3_io_out ? io_r_339_b : _GEN_2678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2680 = 10'h154 == r_count_3_io_out ? io_r_340_b : _GEN_2679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2681 = 10'h155 == r_count_3_io_out ? io_r_341_b : _GEN_2680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2682 = 10'h156 == r_count_3_io_out ? io_r_342_b : _GEN_2681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2683 = 10'h157 == r_count_3_io_out ? io_r_343_b : _GEN_2682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2684 = 10'h158 == r_count_3_io_out ? io_r_344_b : _GEN_2683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2685 = 10'h159 == r_count_3_io_out ? io_r_345_b : _GEN_2684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2686 = 10'h15a == r_count_3_io_out ? io_r_346_b : _GEN_2685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2687 = 10'h15b == r_count_3_io_out ? io_r_347_b : _GEN_2686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2688 = 10'h15c == r_count_3_io_out ? io_r_348_b : _GEN_2687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2689 = 10'h15d == r_count_3_io_out ? io_r_349_b : _GEN_2688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2690 = 10'h15e == r_count_3_io_out ? io_r_350_b : _GEN_2689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2691 = 10'h15f == r_count_3_io_out ? io_r_351_b : _GEN_2690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2692 = 10'h160 == r_count_3_io_out ? io_r_352_b : _GEN_2691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2693 = 10'h161 == r_count_3_io_out ? io_r_353_b : _GEN_2692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2694 = 10'h162 == r_count_3_io_out ? io_r_354_b : _GEN_2693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2695 = 10'h163 == r_count_3_io_out ? io_r_355_b : _GEN_2694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2696 = 10'h164 == r_count_3_io_out ? io_r_356_b : _GEN_2695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2697 = 10'h165 == r_count_3_io_out ? io_r_357_b : _GEN_2696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2698 = 10'h166 == r_count_3_io_out ? io_r_358_b : _GEN_2697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2699 = 10'h167 == r_count_3_io_out ? io_r_359_b : _GEN_2698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2700 = 10'h168 == r_count_3_io_out ? io_r_360_b : _GEN_2699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2701 = 10'h169 == r_count_3_io_out ? io_r_361_b : _GEN_2700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2702 = 10'h16a == r_count_3_io_out ? io_r_362_b : _GEN_2701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2703 = 10'h16b == r_count_3_io_out ? io_r_363_b : _GEN_2702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2704 = 10'h16c == r_count_3_io_out ? io_r_364_b : _GEN_2703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2705 = 10'h16d == r_count_3_io_out ? io_r_365_b : _GEN_2704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2706 = 10'h16e == r_count_3_io_out ? io_r_366_b : _GEN_2705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2707 = 10'h16f == r_count_3_io_out ? io_r_367_b : _GEN_2706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2708 = 10'h170 == r_count_3_io_out ? io_r_368_b : _GEN_2707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2709 = 10'h171 == r_count_3_io_out ? io_r_369_b : _GEN_2708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2710 = 10'h172 == r_count_3_io_out ? io_r_370_b : _GEN_2709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2711 = 10'h173 == r_count_3_io_out ? io_r_371_b : _GEN_2710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2712 = 10'h174 == r_count_3_io_out ? io_r_372_b : _GEN_2711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2713 = 10'h175 == r_count_3_io_out ? io_r_373_b : _GEN_2712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2714 = 10'h176 == r_count_3_io_out ? io_r_374_b : _GEN_2713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2715 = 10'h177 == r_count_3_io_out ? io_r_375_b : _GEN_2714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2716 = 10'h178 == r_count_3_io_out ? io_r_376_b : _GEN_2715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2717 = 10'h179 == r_count_3_io_out ? io_r_377_b : _GEN_2716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2718 = 10'h17a == r_count_3_io_out ? io_r_378_b : _GEN_2717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2719 = 10'h17b == r_count_3_io_out ? io_r_379_b : _GEN_2718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2720 = 10'h17c == r_count_3_io_out ? io_r_380_b : _GEN_2719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2721 = 10'h17d == r_count_3_io_out ? io_r_381_b : _GEN_2720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2722 = 10'h17e == r_count_3_io_out ? io_r_382_b : _GEN_2721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2723 = 10'h17f == r_count_3_io_out ? io_r_383_b : _GEN_2722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2724 = 10'h180 == r_count_3_io_out ? io_r_384_b : _GEN_2723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2725 = 10'h181 == r_count_3_io_out ? io_r_385_b : _GEN_2724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2726 = 10'h182 == r_count_3_io_out ? io_r_386_b : _GEN_2725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2727 = 10'h183 == r_count_3_io_out ? io_r_387_b : _GEN_2726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2728 = 10'h184 == r_count_3_io_out ? io_r_388_b : _GEN_2727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2729 = 10'h185 == r_count_3_io_out ? io_r_389_b : _GEN_2728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2730 = 10'h186 == r_count_3_io_out ? io_r_390_b : _GEN_2729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2731 = 10'h187 == r_count_3_io_out ? io_r_391_b : _GEN_2730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2732 = 10'h188 == r_count_3_io_out ? io_r_392_b : _GEN_2731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2733 = 10'h189 == r_count_3_io_out ? io_r_393_b : _GEN_2732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2734 = 10'h18a == r_count_3_io_out ? io_r_394_b : _GEN_2733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2735 = 10'h18b == r_count_3_io_out ? io_r_395_b : _GEN_2734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2736 = 10'h18c == r_count_3_io_out ? io_r_396_b : _GEN_2735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2737 = 10'h18d == r_count_3_io_out ? io_r_397_b : _GEN_2736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2738 = 10'h18e == r_count_3_io_out ? io_r_398_b : _GEN_2737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2739 = 10'h18f == r_count_3_io_out ? io_r_399_b : _GEN_2738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2740 = 10'h190 == r_count_3_io_out ? io_r_400_b : _GEN_2739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2741 = 10'h191 == r_count_3_io_out ? io_r_401_b : _GEN_2740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2742 = 10'h192 == r_count_3_io_out ? io_r_402_b : _GEN_2741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2743 = 10'h193 == r_count_3_io_out ? io_r_403_b : _GEN_2742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2744 = 10'h194 == r_count_3_io_out ? io_r_404_b : _GEN_2743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2745 = 10'h195 == r_count_3_io_out ? io_r_405_b : _GEN_2744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2746 = 10'h196 == r_count_3_io_out ? io_r_406_b : _GEN_2745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2747 = 10'h197 == r_count_3_io_out ? io_r_407_b : _GEN_2746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2748 = 10'h198 == r_count_3_io_out ? io_r_408_b : _GEN_2747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2749 = 10'h199 == r_count_3_io_out ? io_r_409_b : _GEN_2748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2750 = 10'h19a == r_count_3_io_out ? io_r_410_b : _GEN_2749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2751 = 10'h19b == r_count_3_io_out ? io_r_411_b : _GEN_2750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2752 = 10'h19c == r_count_3_io_out ? io_r_412_b : _GEN_2751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2753 = 10'h19d == r_count_3_io_out ? io_r_413_b : _GEN_2752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2754 = 10'h19e == r_count_3_io_out ? io_r_414_b : _GEN_2753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2755 = 10'h19f == r_count_3_io_out ? io_r_415_b : _GEN_2754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2756 = 10'h1a0 == r_count_3_io_out ? io_r_416_b : _GEN_2755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2757 = 10'h1a1 == r_count_3_io_out ? io_r_417_b : _GEN_2756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2758 = 10'h1a2 == r_count_3_io_out ? io_r_418_b : _GEN_2757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2759 = 10'h1a3 == r_count_3_io_out ? io_r_419_b : _GEN_2758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2760 = 10'h1a4 == r_count_3_io_out ? io_r_420_b : _GEN_2759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2761 = 10'h1a5 == r_count_3_io_out ? io_r_421_b : _GEN_2760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2762 = 10'h1a6 == r_count_3_io_out ? io_r_422_b : _GEN_2761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2763 = 10'h1a7 == r_count_3_io_out ? io_r_423_b : _GEN_2762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2764 = 10'h1a8 == r_count_3_io_out ? io_r_424_b : _GEN_2763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2765 = 10'h1a9 == r_count_3_io_out ? io_r_425_b : _GEN_2764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2766 = 10'h1aa == r_count_3_io_out ? io_r_426_b : _GEN_2765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2767 = 10'h1ab == r_count_3_io_out ? io_r_427_b : _GEN_2766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2768 = 10'h1ac == r_count_3_io_out ? io_r_428_b : _GEN_2767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2769 = 10'h1ad == r_count_3_io_out ? io_r_429_b : _GEN_2768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2770 = 10'h1ae == r_count_3_io_out ? io_r_430_b : _GEN_2769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2771 = 10'h1af == r_count_3_io_out ? io_r_431_b : _GEN_2770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2772 = 10'h1b0 == r_count_3_io_out ? io_r_432_b : _GEN_2771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2773 = 10'h1b1 == r_count_3_io_out ? io_r_433_b : _GEN_2772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2774 = 10'h1b2 == r_count_3_io_out ? io_r_434_b : _GEN_2773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2775 = 10'h1b3 == r_count_3_io_out ? io_r_435_b : _GEN_2774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2776 = 10'h1b4 == r_count_3_io_out ? io_r_436_b : _GEN_2775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2777 = 10'h1b5 == r_count_3_io_out ? io_r_437_b : _GEN_2776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2778 = 10'h1b6 == r_count_3_io_out ? io_r_438_b : _GEN_2777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2779 = 10'h1b7 == r_count_3_io_out ? io_r_439_b : _GEN_2778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2780 = 10'h1b8 == r_count_3_io_out ? io_r_440_b : _GEN_2779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2781 = 10'h1b9 == r_count_3_io_out ? io_r_441_b : _GEN_2780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2782 = 10'h1ba == r_count_3_io_out ? io_r_442_b : _GEN_2781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2783 = 10'h1bb == r_count_3_io_out ? io_r_443_b : _GEN_2782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2784 = 10'h1bc == r_count_3_io_out ? io_r_444_b : _GEN_2783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2785 = 10'h1bd == r_count_3_io_out ? io_r_445_b : _GEN_2784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2786 = 10'h1be == r_count_3_io_out ? io_r_446_b : _GEN_2785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2787 = 10'h1bf == r_count_3_io_out ? io_r_447_b : _GEN_2786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2788 = 10'h1c0 == r_count_3_io_out ? io_r_448_b : _GEN_2787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2789 = 10'h1c1 == r_count_3_io_out ? io_r_449_b : _GEN_2788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2790 = 10'h1c2 == r_count_3_io_out ? io_r_450_b : _GEN_2789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2791 = 10'h1c3 == r_count_3_io_out ? io_r_451_b : _GEN_2790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2792 = 10'h1c4 == r_count_3_io_out ? io_r_452_b : _GEN_2791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2793 = 10'h1c5 == r_count_3_io_out ? io_r_453_b : _GEN_2792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2794 = 10'h1c6 == r_count_3_io_out ? io_r_454_b : _GEN_2793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2795 = 10'h1c7 == r_count_3_io_out ? io_r_455_b : _GEN_2794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2796 = 10'h1c8 == r_count_3_io_out ? io_r_456_b : _GEN_2795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2797 = 10'h1c9 == r_count_3_io_out ? io_r_457_b : _GEN_2796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2798 = 10'h1ca == r_count_3_io_out ? io_r_458_b : _GEN_2797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2799 = 10'h1cb == r_count_3_io_out ? io_r_459_b : _GEN_2798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2800 = 10'h1cc == r_count_3_io_out ? io_r_460_b : _GEN_2799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2801 = 10'h1cd == r_count_3_io_out ? io_r_461_b : _GEN_2800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2802 = 10'h1ce == r_count_3_io_out ? io_r_462_b : _GEN_2801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2803 = 10'h1cf == r_count_3_io_out ? io_r_463_b : _GEN_2802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2804 = 10'h1d0 == r_count_3_io_out ? io_r_464_b : _GEN_2803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2805 = 10'h1d1 == r_count_3_io_out ? io_r_465_b : _GEN_2804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2806 = 10'h1d2 == r_count_3_io_out ? io_r_466_b : _GEN_2805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2807 = 10'h1d3 == r_count_3_io_out ? io_r_467_b : _GEN_2806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2808 = 10'h1d4 == r_count_3_io_out ? io_r_468_b : _GEN_2807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2809 = 10'h1d5 == r_count_3_io_out ? io_r_469_b : _GEN_2808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2810 = 10'h1d6 == r_count_3_io_out ? io_r_470_b : _GEN_2809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2811 = 10'h1d7 == r_count_3_io_out ? io_r_471_b : _GEN_2810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2812 = 10'h1d8 == r_count_3_io_out ? io_r_472_b : _GEN_2811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2813 = 10'h1d9 == r_count_3_io_out ? io_r_473_b : _GEN_2812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2814 = 10'h1da == r_count_3_io_out ? io_r_474_b : _GEN_2813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2815 = 10'h1db == r_count_3_io_out ? io_r_475_b : _GEN_2814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2816 = 10'h1dc == r_count_3_io_out ? io_r_476_b : _GEN_2815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2817 = 10'h1dd == r_count_3_io_out ? io_r_477_b : _GEN_2816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2818 = 10'h1de == r_count_3_io_out ? io_r_478_b : _GEN_2817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2819 = 10'h1df == r_count_3_io_out ? io_r_479_b : _GEN_2818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2820 = 10'h1e0 == r_count_3_io_out ? io_r_480_b : _GEN_2819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2821 = 10'h1e1 == r_count_3_io_out ? io_r_481_b : _GEN_2820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2822 = 10'h1e2 == r_count_3_io_out ? io_r_482_b : _GEN_2821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2823 = 10'h1e3 == r_count_3_io_out ? io_r_483_b : _GEN_2822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2824 = 10'h1e4 == r_count_3_io_out ? io_r_484_b : _GEN_2823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2825 = 10'h1e5 == r_count_3_io_out ? io_r_485_b : _GEN_2824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2826 = 10'h1e6 == r_count_3_io_out ? io_r_486_b : _GEN_2825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2827 = 10'h1e7 == r_count_3_io_out ? io_r_487_b : _GEN_2826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2828 = 10'h1e8 == r_count_3_io_out ? io_r_488_b : _GEN_2827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2829 = 10'h1e9 == r_count_3_io_out ? io_r_489_b : _GEN_2828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2830 = 10'h1ea == r_count_3_io_out ? io_r_490_b : _GEN_2829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2831 = 10'h1eb == r_count_3_io_out ? io_r_491_b : _GEN_2830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2832 = 10'h1ec == r_count_3_io_out ? io_r_492_b : _GEN_2831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2833 = 10'h1ed == r_count_3_io_out ? io_r_493_b : _GEN_2832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2834 = 10'h1ee == r_count_3_io_out ? io_r_494_b : _GEN_2833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2835 = 10'h1ef == r_count_3_io_out ? io_r_495_b : _GEN_2834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2836 = 10'h1f0 == r_count_3_io_out ? io_r_496_b : _GEN_2835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2837 = 10'h1f1 == r_count_3_io_out ? io_r_497_b : _GEN_2836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2838 = 10'h1f2 == r_count_3_io_out ? io_r_498_b : _GEN_2837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2839 = 10'h1f3 == r_count_3_io_out ? io_r_499_b : _GEN_2838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2840 = 10'h1f4 == r_count_3_io_out ? io_r_500_b : _GEN_2839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2841 = 10'h1f5 == r_count_3_io_out ? io_r_501_b : _GEN_2840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2842 = 10'h1f6 == r_count_3_io_out ? io_r_502_b : _GEN_2841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2843 = 10'h1f7 == r_count_3_io_out ? io_r_503_b : _GEN_2842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2844 = 10'h1f8 == r_count_3_io_out ? io_r_504_b : _GEN_2843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2845 = 10'h1f9 == r_count_3_io_out ? io_r_505_b : _GEN_2844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2846 = 10'h1fa == r_count_3_io_out ? io_r_506_b : _GEN_2845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2847 = 10'h1fb == r_count_3_io_out ? io_r_507_b : _GEN_2846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2848 = 10'h1fc == r_count_3_io_out ? io_r_508_b : _GEN_2847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2849 = 10'h1fd == r_count_3_io_out ? io_r_509_b : _GEN_2848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2850 = 10'h1fe == r_count_3_io_out ? io_r_510_b : _GEN_2849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2851 = 10'h1ff == r_count_3_io_out ? io_r_511_b : _GEN_2850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2852 = 10'h200 == r_count_3_io_out ? io_r_512_b : _GEN_2851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2853 = 10'h201 == r_count_3_io_out ? io_r_513_b : _GEN_2852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2854 = 10'h202 == r_count_3_io_out ? io_r_514_b : _GEN_2853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2855 = 10'h203 == r_count_3_io_out ? io_r_515_b : _GEN_2854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2856 = 10'h204 == r_count_3_io_out ? io_r_516_b : _GEN_2855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2857 = 10'h205 == r_count_3_io_out ? io_r_517_b : _GEN_2856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2858 = 10'h206 == r_count_3_io_out ? io_r_518_b : _GEN_2857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2859 = 10'h207 == r_count_3_io_out ? io_r_519_b : _GEN_2858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2860 = 10'h208 == r_count_3_io_out ? io_r_520_b : _GEN_2859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2861 = 10'h209 == r_count_3_io_out ? io_r_521_b : _GEN_2860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2862 = 10'h20a == r_count_3_io_out ? io_r_522_b : _GEN_2861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2863 = 10'h20b == r_count_3_io_out ? io_r_523_b : _GEN_2862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2864 = 10'h20c == r_count_3_io_out ? io_r_524_b : _GEN_2863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2865 = 10'h20d == r_count_3_io_out ? io_r_525_b : _GEN_2864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2866 = 10'h20e == r_count_3_io_out ? io_r_526_b : _GEN_2865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2867 = 10'h20f == r_count_3_io_out ? io_r_527_b : _GEN_2866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2868 = 10'h210 == r_count_3_io_out ? io_r_528_b : _GEN_2867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2869 = 10'h211 == r_count_3_io_out ? io_r_529_b : _GEN_2868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2870 = 10'h212 == r_count_3_io_out ? io_r_530_b : _GEN_2869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2871 = 10'h213 == r_count_3_io_out ? io_r_531_b : _GEN_2870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2872 = 10'h214 == r_count_3_io_out ? io_r_532_b : _GEN_2871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2873 = 10'h215 == r_count_3_io_out ? io_r_533_b : _GEN_2872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2874 = 10'h216 == r_count_3_io_out ? io_r_534_b : _GEN_2873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2875 = 10'h217 == r_count_3_io_out ? io_r_535_b : _GEN_2874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2876 = 10'h218 == r_count_3_io_out ? io_r_536_b : _GEN_2875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2877 = 10'h219 == r_count_3_io_out ? io_r_537_b : _GEN_2876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2878 = 10'h21a == r_count_3_io_out ? io_r_538_b : _GEN_2877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2879 = 10'h21b == r_count_3_io_out ? io_r_539_b : _GEN_2878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2880 = 10'h21c == r_count_3_io_out ? io_r_540_b : _GEN_2879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2881 = 10'h21d == r_count_3_io_out ? io_r_541_b : _GEN_2880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2882 = 10'h21e == r_count_3_io_out ? io_r_542_b : _GEN_2881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2883 = 10'h21f == r_count_3_io_out ? io_r_543_b : _GEN_2882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2884 = 10'h220 == r_count_3_io_out ? io_r_544_b : _GEN_2883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2885 = 10'h221 == r_count_3_io_out ? io_r_545_b : _GEN_2884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2886 = 10'h222 == r_count_3_io_out ? io_r_546_b : _GEN_2885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2887 = 10'h223 == r_count_3_io_out ? io_r_547_b : _GEN_2886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2888 = 10'h224 == r_count_3_io_out ? io_r_548_b : _GEN_2887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2889 = 10'h225 == r_count_3_io_out ? io_r_549_b : _GEN_2888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2890 = 10'h226 == r_count_3_io_out ? io_r_550_b : _GEN_2889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2891 = 10'h227 == r_count_3_io_out ? io_r_551_b : _GEN_2890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2892 = 10'h228 == r_count_3_io_out ? io_r_552_b : _GEN_2891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2893 = 10'h229 == r_count_3_io_out ? io_r_553_b : _GEN_2892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2894 = 10'h22a == r_count_3_io_out ? io_r_554_b : _GEN_2893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2895 = 10'h22b == r_count_3_io_out ? io_r_555_b : _GEN_2894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2896 = 10'h22c == r_count_3_io_out ? io_r_556_b : _GEN_2895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2897 = 10'h22d == r_count_3_io_out ? io_r_557_b : _GEN_2896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2898 = 10'h22e == r_count_3_io_out ? io_r_558_b : _GEN_2897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2899 = 10'h22f == r_count_3_io_out ? io_r_559_b : _GEN_2898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2900 = 10'h230 == r_count_3_io_out ? io_r_560_b : _GEN_2899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2901 = 10'h231 == r_count_3_io_out ? io_r_561_b : _GEN_2900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2902 = 10'h232 == r_count_3_io_out ? io_r_562_b : _GEN_2901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2903 = 10'h233 == r_count_3_io_out ? io_r_563_b : _GEN_2902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2904 = 10'h234 == r_count_3_io_out ? io_r_564_b : _GEN_2903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2905 = 10'h235 == r_count_3_io_out ? io_r_565_b : _GEN_2904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2906 = 10'h236 == r_count_3_io_out ? io_r_566_b : _GEN_2905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2907 = 10'h237 == r_count_3_io_out ? io_r_567_b : _GEN_2906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2908 = 10'h238 == r_count_3_io_out ? io_r_568_b : _GEN_2907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2909 = 10'h239 == r_count_3_io_out ? io_r_569_b : _GEN_2908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2910 = 10'h23a == r_count_3_io_out ? io_r_570_b : _GEN_2909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2911 = 10'h23b == r_count_3_io_out ? io_r_571_b : _GEN_2910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2912 = 10'h23c == r_count_3_io_out ? io_r_572_b : _GEN_2911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2913 = 10'h23d == r_count_3_io_out ? io_r_573_b : _GEN_2912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2914 = 10'h23e == r_count_3_io_out ? io_r_574_b : _GEN_2913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2915 = 10'h23f == r_count_3_io_out ? io_r_575_b : _GEN_2914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2916 = 10'h240 == r_count_3_io_out ? io_r_576_b : _GEN_2915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2917 = 10'h241 == r_count_3_io_out ? io_r_577_b : _GEN_2916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2918 = 10'h242 == r_count_3_io_out ? io_r_578_b : _GEN_2917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2919 = 10'h243 == r_count_3_io_out ? io_r_579_b : _GEN_2918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2920 = 10'h244 == r_count_3_io_out ? io_r_580_b : _GEN_2919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2921 = 10'h245 == r_count_3_io_out ? io_r_581_b : _GEN_2920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2922 = 10'h246 == r_count_3_io_out ? io_r_582_b : _GEN_2921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2923 = 10'h247 == r_count_3_io_out ? io_r_583_b : _GEN_2922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2924 = 10'h248 == r_count_3_io_out ? io_r_584_b : _GEN_2923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2925 = 10'h249 == r_count_3_io_out ? io_r_585_b : _GEN_2924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2926 = 10'h24a == r_count_3_io_out ? io_r_586_b : _GEN_2925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2927 = 10'h24b == r_count_3_io_out ? io_r_587_b : _GEN_2926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2928 = 10'h24c == r_count_3_io_out ? io_r_588_b : _GEN_2927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2929 = 10'h24d == r_count_3_io_out ? io_r_589_b : _GEN_2928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2930 = 10'h24e == r_count_3_io_out ? io_r_590_b : _GEN_2929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2931 = 10'h24f == r_count_3_io_out ? io_r_591_b : _GEN_2930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2932 = 10'h250 == r_count_3_io_out ? io_r_592_b : _GEN_2931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2933 = 10'h251 == r_count_3_io_out ? io_r_593_b : _GEN_2932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2934 = 10'h252 == r_count_3_io_out ? io_r_594_b : _GEN_2933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2935 = 10'h253 == r_count_3_io_out ? io_r_595_b : _GEN_2934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2936 = 10'h254 == r_count_3_io_out ? io_r_596_b : _GEN_2935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2937 = 10'h255 == r_count_3_io_out ? io_r_597_b : _GEN_2936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2938 = 10'h256 == r_count_3_io_out ? io_r_598_b : _GEN_2937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2939 = 10'h257 == r_count_3_io_out ? io_r_599_b : _GEN_2938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2940 = 10'h258 == r_count_3_io_out ? io_r_600_b : _GEN_2939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2941 = 10'h259 == r_count_3_io_out ? io_r_601_b : _GEN_2940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2942 = 10'h25a == r_count_3_io_out ? io_r_602_b : _GEN_2941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2943 = 10'h25b == r_count_3_io_out ? io_r_603_b : _GEN_2942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2944 = 10'h25c == r_count_3_io_out ? io_r_604_b : _GEN_2943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2945 = 10'h25d == r_count_3_io_out ? io_r_605_b : _GEN_2944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2946 = 10'h25e == r_count_3_io_out ? io_r_606_b : _GEN_2945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2947 = 10'h25f == r_count_3_io_out ? io_r_607_b : _GEN_2946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2948 = 10'h260 == r_count_3_io_out ? io_r_608_b : _GEN_2947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2949 = 10'h261 == r_count_3_io_out ? io_r_609_b : _GEN_2948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2950 = 10'h262 == r_count_3_io_out ? io_r_610_b : _GEN_2949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2951 = 10'h263 == r_count_3_io_out ? io_r_611_b : _GEN_2950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2952 = 10'h264 == r_count_3_io_out ? io_r_612_b : _GEN_2951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2953 = 10'h265 == r_count_3_io_out ? io_r_613_b : _GEN_2952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2954 = 10'h266 == r_count_3_io_out ? io_r_614_b : _GEN_2953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2955 = 10'h267 == r_count_3_io_out ? io_r_615_b : _GEN_2954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2956 = 10'h268 == r_count_3_io_out ? io_r_616_b : _GEN_2955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2957 = 10'h269 == r_count_3_io_out ? io_r_617_b : _GEN_2956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2958 = 10'h26a == r_count_3_io_out ? io_r_618_b : _GEN_2957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2959 = 10'h26b == r_count_3_io_out ? io_r_619_b : _GEN_2958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2960 = 10'h26c == r_count_3_io_out ? io_r_620_b : _GEN_2959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2961 = 10'h26d == r_count_3_io_out ? io_r_621_b : _GEN_2960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2962 = 10'h26e == r_count_3_io_out ? io_r_622_b : _GEN_2961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2963 = 10'h26f == r_count_3_io_out ? io_r_623_b : _GEN_2962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2964 = 10'h270 == r_count_3_io_out ? io_r_624_b : _GEN_2963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2965 = 10'h271 == r_count_3_io_out ? io_r_625_b : _GEN_2964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2966 = 10'h272 == r_count_3_io_out ? io_r_626_b : _GEN_2965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2967 = 10'h273 == r_count_3_io_out ? io_r_627_b : _GEN_2966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2968 = 10'h274 == r_count_3_io_out ? io_r_628_b : _GEN_2967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2969 = 10'h275 == r_count_3_io_out ? io_r_629_b : _GEN_2968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2970 = 10'h276 == r_count_3_io_out ? io_r_630_b : _GEN_2969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2971 = 10'h277 == r_count_3_io_out ? io_r_631_b : _GEN_2970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2972 = 10'h278 == r_count_3_io_out ? io_r_632_b : _GEN_2971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2973 = 10'h279 == r_count_3_io_out ? io_r_633_b : _GEN_2972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2974 = 10'h27a == r_count_3_io_out ? io_r_634_b : _GEN_2973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2975 = 10'h27b == r_count_3_io_out ? io_r_635_b : _GEN_2974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2976 = 10'h27c == r_count_3_io_out ? io_r_636_b : _GEN_2975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2977 = 10'h27d == r_count_3_io_out ? io_r_637_b : _GEN_2976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2978 = 10'h27e == r_count_3_io_out ? io_r_638_b : _GEN_2977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2979 = 10'h27f == r_count_3_io_out ? io_r_639_b : _GEN_2978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2980 = 10'h280 == r_count_3_io_out ? io_r_640_b : _GEN_2979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2981 = 10'h281 == r_count_3_io_out ? io_r_641_b : _GEN_2980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2982 = 10'h282 == r_count_3_io_out ? io_r_642_b : _GEN_2981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2983 = 10'h283 == r_count_3_io_out ? io_r_643_b : _GEN_2982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2984 = 10'h284 == r_count_3_io_out ? io_r_644_b : _GEN_2983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2985 = 10'h285 == r_count_3_io_out ? io_r_645_b : _GEN_2984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2986 = 10'h286 == r_count_3_io_out ? io_r_646_b : _GEN_2985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2987 = 10'h287 == r_count_3_io_out ? io_r_647_b : _GEN_2986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2988 = 10'h288 == r_count_3_io_out ? io_r_648_b : _GEN_2987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2989 = 10'h289 == r_count_3_io_out ? io_r_649_b : _GEN_2988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2990 = 10'h28a == r_count_3_io_out ? io_r_650_b : _GEN_2989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2991 = 10'h28b == r_count_3_io_out ? io_r_651_b : _GEN_2990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2992 = 10'h28c == r_count_3_io_out ? io_r_652_b : _GEN_2991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2993 = 10'h28d == r_count_3_io_out ? io_r_653_b : _GEN_2992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2994 = 10'h28e == r_count_3_io_out ? io_r_654_b : _GEN_2993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2995 = 10'h28f == r_count_3_io_out ? io_r_655_b : _GEN_2994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2996 = 10'h290 == r_count_3_io_out ? io_r_656_b : _GEN_2995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2997 = 10'h291 == r_count_3_io_out ? io_r_657_b : _GEN_2996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2998 = 10'h292 == r_count_3_io_out ? io_r_658_b : _GEN_2997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2999 = 10'h293 == r_count_3_io_out ? io_r_659_b : _GEN_2998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3000 = 10'h294 == r_count_3_io_out ? io_r_660_b : _GEN_2999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3001 = 10'h295 == r_count_3_io_out ? io_r_661_b : _GEN_3000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3002 = 10'h296 == r_count_3_io_out ? io_r_662_b : _GEN_3001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3003 = 10'h297 == r_count_3_io_out ? io_r_663_b : _GEN_3002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3004 = 10'h298 == r_count_3_io_out ? io_r_664_b : _GEN_3003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3005 = 10'h299 == r_count_3_io_out ? io_r_665_b : _GEN_3004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3006 = 10'h29a == r_count_3_io_out ? io_r_666_b : _GEN_3005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3007 = 10'h29b == r_count_3_io_out ? io_r_667_b : _GEN_3006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3008 = 10'h29c == r_count_3_io_out ? io_r_668_b : _GEN_3007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3009 = 10'h29d == r_count_3_io_out ? io_r_669_b : _GEN_3008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3010 = 10'h29e == r_count_3_io_out ? io_r_670_b : _GEN_3009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3011 = 10'h29f == r_count_3_io_out ? io_r_671_b : _GEN_3010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3012 = 10'h2a0 == r_count_3_io_out ? io_r_672_b : _GEN_3011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3013 = 10'h2a1 == r_count_3_io_out ? io_r_673_b : _GEN_3012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3014 = 10'h2a2 == r_count_3_io_out ? io_r_674_b : _GEN_3013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3015 = 10'h2a3 == r_count_3_io_out ? io_r_675_b : _GEN_3014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3016 = 10'h2a4 == r_count_3_io_out ? io_r_676_b : _GEN_3015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3017 = 10'h2a5 == r_count_3_io_out ? io_r_677_b : _GEN_3016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3018 = 10'h2a6 == r_count_3_io_out ? io_r_678_b : _GEN_3017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3019 = 10'h2a7 == r_count_3_io_out ? io_r_679_b : _GEN_3018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3020 = 10'h2a8 == r_count_3_io_out ? io_r_680_b : _GEN_3019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3021 = 10'h2a9 == r_count_3_io_out ? io_r_681_b : _GEN_3020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3022 = 10'h2aa == r_count_3_io_out ? io_r_682_b : _GEN_3021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3023 = 10'h2ab == r_count_3_io_out ? io_r_683_b : _GEN_3022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3024 = 10'h2ac == r_count_3_io_out ? io_r_684_b : _GEN_3023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3025 = 10'h2ad == r_count_3_io_out ? io_r_685_b : _GEN_3024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3026 = 10'h2ae == r_count_3_io_out ? io_r_686_b : _GEN_3025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3027 = 10'h2af == r_count_3_io_out ? io_r_687_b : _GEN_3026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3028 = 10'h2b0 == r_count_3_io_out ? io_r_688_b : _GEN_3027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3029 = 10'h2b1 == r_count_3_io_out ? io_r_689_b : _GEN_3028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3030 = 10'h2b2 == r_count_3_io_out ? io_r_690_b : _GEN_3029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3031 = 10'h2b3 == r_count_3_io_out ? io_r_691_b : _GEN_3030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3032 = 10'h2b4 == r_count_3_io_out ? io_r_692_b : _GEN_3031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3033 = 10'h2b5 == r_count_3_io_out ? io_r_693_b : _GEN_3032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3034 = 10'h2b6 == r_count_3_io_out ? io_r_694_b : _GEN_3033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3035 = 10'h2b7 == r_count_3_io_out ? io_r_695_b : _GEN_3034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3036 = 10'h2b8 == r_count_3_io_out ? io_r_696_b : _GEN_3035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3037 = 10'h2b9 == r_count_3_io_out ? io_r_697_b : _GEN_3036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3038 = 10'h2ba == r_count_3_io_out ? io_r_698_b : _GEN_3037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3039 = 10'h2bb == r_count_3_io_out ? io_r_699_b : _GEN_3038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3040 = 10'h2bc == r_count_3_io_out ? io_r_700_b : _GEN_3039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3041 = 10'h2bd == r_count_3_io_out ? io_r_701_b : _GEN_3040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3042 = 10'h2be == r_count_3_io_out ? io_r_702_b : _GEN_3041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3043 = 10'h2bf == r_count_3_io_out ? io_r_703_b : _GEN_3042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3044 = 10'h2c0 == r_count_3_io_out ? io_r_704_b : _GEN_3043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3045 = 10'h2c1 == r_count_3_io_out ? io_r_705_b : _GEN_3044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3046 = 10'h2c2 == r_count_3_io_out ? io_r_706_b : _GEN_3045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3047 = 10'h2c3 == r_count_3_io_out ? io_r_707_b : _GEN_3046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3048 = 10'h2c4 == r_count_3_io_out ? io_r_708_b : _GEN_3047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3049 = 10'h2c5 == r_count_3_io_out ? io_r_709_b : _GEN_3048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3050 = 10'h2c6 == r_count_3_io_out ? io_r_710_b : _GEN_3049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3051 = 10'h2c7 == r_count_3_io_out ? io_r_711_b : _GEN_3050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3052 = 10'h2c8 == r_count_3_io_out ? io_r_712_b : _GEN_3051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3053 = 10'h2c9 == r_count_3_io_out ? io_r_713_b : _GEN_3052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3054 = 10'h2ca == r_count_3_io_out ? io_r_714_b : _GEN_3053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3055 = 10'h2cb == r_count_3_io_out ? io_r_715_b : _GEN_3054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3056 = 10'h2cc == r_count_3_io_out ? io_r_716_b : _GEN_3055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3057 = 10'h2cd == r_count_3_io_out ? io_r_717_b : _GEN_3056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3058 = 10'h2ce == r_count_3_io_out ? io_r_718_b : _GEN_3057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3059 = 10'h2cf == r_count_3_io_out ? io_r_719_b : _GEN_3058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3060 = 10'h2d0 == r_count_3_io_out ? io_r_720_b : _GEN_3059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3061 = 10'h2d1 == r_count_3_io_out ? io_r_721_b : _GEN_3060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3062 = 10'h2d2 == r_count_3_io_out ? io_r_722_b : _GEN_3061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3063 = 10'h2d3 == r_count_3_io_out ? io_r_723_b : _GEN_3062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3064 = 10'h2d4 == r_count_3_io_out ? io_r_724_b : _GEN_3063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3065 = 10'h2d5 == r_count_3_io_out ? io_r_725_b : _GEN_3064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3066 = 10'h2d6 == r_count_3_io_out ? io_r_726_b : _GEN_3065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3067 = 10'h2d7 == r_count_3_io_out ? io_r_727_b : _GEN_3066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3068 = 10'h2d8 == r_count_3_io_out ? io_r_728_b : _GEN_3067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3069 = 10'h2d9 == r_count_3_io_out ? io_r_729_b : _GEN_3068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3070 = 10'h2da == r_count_3_io_out ? io_r_730_b : _GEN_3069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3071 = 10'h2db == r_count_3_io_out ? io_r_731_b : _GEN_3070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3072 = 10'h2dc == r_count_3_io_out ? io_r_732_b : _GEN_3071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3073 = 10'h2dd == r_count_3_io_out ? io_r_733_b : _GEN_3072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3074 = 10'h2de == r_count_3_io_out ? io_r_734_b : _GEN_3073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3075 = 10'h2df == r_count_3_io_out ? io_r_735_b : _GEN_3074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3076 = 10'h2e0 == r_count_3_io_out ? io_r_736_b : _GEN_3075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3077 = 10'h2e1 == r_count_3_io_out ? io_r_737_b : _GEN_3076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3078 = 10'h2e2 == r_count_3_io_out ? io_r_738_b : _GEN_3077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3079 = 10'h2e3 == r_count_3_io_out ? io_r_739_b : _GEN_3078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3080 = 10'h2e4 == r_count_3_io_out ? io_r_740_b : _GEN_3079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3081 = 10'h2e5 == r_count_3_io_out ? io_r_741_b : _GEN_3080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3082 = 10'h2e6 == r_count_3_io_out ? io_r_742_b : _GEN_3081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3083 = 10'h2e7 == r_count_3_io_out ? io_r_743_b : _GEN_3082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3084 = 10'h2e8 == r_count_3_io_out ? io_r_744_b : _GEN_3083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3085 = 10'h2e9 == r_count_3_io_out ? io_r_745_b : _GEN_3084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3086 = 10'h2ea == r_count_3_io_out ? io_r_746_b : _GEN_3085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3087 = 10'h2eb == r_count_3_io_out ? io_r_747_b : _GEN_3086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3088 = 10'h2ec == r_count_3_io_out ? io_r_748_b : _GEN_3087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3091 = 10'h1 == r_count_4_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3092 = 10'h2 == r_count_4_io_out ? io_r_2_b : _GEN_3091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3093 = 10'h3 == r_count_4_io_out ? io_r_3_b : _GEN_3092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3094 = 10'h4 == r_count_4_io_out ? io_r_4_b : _GEN_3093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3095 = 10'h5 == r_count_4_io_out ? io_r_5_b : _GEN_3094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3096 = 10'h6 == r_count_4_io_out ? io_r_6_b : _GEN_3095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3097 = 10'h7 == r_count_4_io_out ? io_r_7_b : _GEN_3096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3098 = 10'h8 == r_count_4_io_out ? io_r_8_b : _GEN_3097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3099 = 10'h9 == r_count_4_io_out ? io_r_9_b : _GEN_3098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3100 = 10'ha == r_count_4_io_out ? io_r_10_b : _GEN_3099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3101 = 10'hb == r_count_4_io_out ? io_r_11_b : _GEN_3100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3102 = 10'hc == r_count_4_io_out ? io_r_12_b : _GEN_3101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3103 = 10'hd == r_count_4_io_out ? io_r_13_b : _GEN_3102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3104 = 10'he == r_count_4_io_out ? io_r_14_b : _GEN_3103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3105 = 10'hf == r_count_4_io_out ? io_r_15_b : _GEN_3104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3106 = 10'h10 == r_count_4_io_out ? io_r_16_b : _GEN_3105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3107 = 10'h11 == r_count_4_io_out ? io_r_17_b : _GEN_3106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3108 = 10'h12 == r_count_4_io_out ? io_r_18_b : _GEN_3107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3109 = 10'h13 == r_count_4_io_out ? io_r_19_b : _GEN_3108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3110 = 10'h14 == r_count_4_io_out ? io_r_20_b : _GEN_3109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3111 = 10'h15 == r_count_4_io_out ? io_r_21_b : _GEN_3110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3112 = 10'h16 == r_count_4_io_out ? io_r_22_b : _GEN_3111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3113 = 10'h17 == r_count_4_io_out ? io_r_23_b : _GEN_3112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3114 = 10'h18 == r_count_4_io_out ? io_r_24_b : _GEN_3113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3115 = 10'h19 == r_count_4_io_out ? io_r_25_b : _GEN_3114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3116 = 10'h1a == r_count_4_io_out ? io_r_26_b : _GEN_3115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3117 = 10'h1b == r_count_4_io_out ? io_r_27_b : _GEN_3116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3118 = 10'h1c == r_count_4_io_out ? io_r_28_b : _GEN_3117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3119 = 10'h1d == r_count_4_io_out ? io_r_29_b : _GEN_3118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3120 = 10'h1e == r_count_4_io_out ? io_r_30_b : _GEN_3119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3121 = 10'h1f == r_count_4_io_out ? io_r_31_b : _GEN_3120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3122 = 10'h20 == r_count_4_io_out ? io_r_32_b : _GEN_3121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3123 = 10'h21 == r_count_4_io_out ? io_r_33_b : _GEN_3122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3124 = 10'h22 == r_count_4_io_out ? io_r_34_b : _GEN_3123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3125 = 10'h23 == r_count_4_io_out ? io_r_35_b : _GEN_3124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3126 = 10'h24 == r_count_4_io_out ? io_r_36_b : _GEN_3125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3127 = 10'h25 == r_count_4_io_out ? io_r_37_b : _GEN_3126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3128 = 10'h26 == r_count_4_io_out ? io_r_38_b : _GEN_3127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3129 = 10'h27 == r_count_4_io_out ? io_r_39_b : _GEN_3128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3130 = 10'h28 == r_count_4_io_out ? io_r_40_b : _GEN_3129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3131 = 10'h29 == r_count_4_io_out ? io_r_41_b : _GEN_3130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3132 = 10'h2a == r_count_4_io_out ? io_r_42_b : _GEN_3131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3133 = 10'h2b == r_count_4_io_out ? io_r_43_b : _GEN_3132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3134 = 10'h2c == r_count_4_io_out ? io_r_44_b : _GEN_3133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3135 = 10'h2d == r_count_4_io_out ? io_r_45_b : _GEN_3134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3136 = 10'h2e == r_count_4_io_out ? io_r_46_b : _GEN_3135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3137 = 10'h2f == r_count_4_io_out ? io_r_47_b : _GEN_3136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3138 = 10'h30 == r_count_4_io_out ? io_r_48_b : _GEN_3137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3139 = 10'h31 == r_count_4_io_out ? io_r_49_b : _GEN_3138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3140 = 10'h32 == r_count_4_io_out ? io_r_50_b : _GEN_3139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3141 = 10'h33 == r_count_4_io_out ? io_r_51_b : _GEN_3140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3142 = 10'h34 == r_count_4_io_out ? io_r_52_b : _GEN_3141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3143 = 10'h35 == r_count_4_io_out ? io_r_53_b : _GEN_3142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3144 = 10'h36 == r_count_4_io_out ? io_r_54_b : _GEN_3143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3145 = 10'h37 == r_count_4_io_out ? io_r_55_b : _GEN_3144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3146 = 10'h38 == r_count_4_io_out ? io_r_56_b : _GEN_3145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3147 = 10'h39 == r_count_4_io_out ? io_r_57_b : _GEN_3146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3148 = 10'h3a == r_count_4_io_out ? io_r_58_b : _GEN_3147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3149 = 10'h3b == r_count_4_io_out ? io_r_59_b : _GEN_3148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3150 = 10'h3c == r_count_4_io_out ? io_r_60_b : _GEN_3149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3151 = 10'h3d == r_count_4_io_out ? io_r_61_b : _GEN_3150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3152 = 10'h3e == r_count_4_io_out ? io_r_62_b : _GEN_3151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3153 = 10'h3f == r_count_4_io_out ? io_r_63_b : _GEN_3152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3154 = 10'h40 == r_count_4_io_out ? io_r_64_b : _GEN_3153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3155 = 10'h41 == r_count_4_io_out ? io_r_65_b : _GEN_3154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3156 = 10'h42 == r_count_4_io_out ? io_r_66_b : _GEN_3155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3157 = 10'h43 == r_count_4_io_out ? io_r_67_b : _GEN_3156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3158 = 10'h44 == r_count_4_io_out ? io_r_68_b : _GEN_3157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3159 = 10'h45 == r_count_4_io_out ? io_r_69_b : _GEN_3158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3160 = 10'h46 == r_count_4_io_out ? io_r_70_b : _GEN_3159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3161 = 10'h47 == r_count_4_io_out ? io_r_71_b : _GEN_3160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3162 = 10'h48 == r_count_4_io_out ? io_r_72_b : _GEN_3161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3163 = 10'h49 == r_count_4_io_out ? io_r_73_b : _GEN_3162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3164 = 10'h4a == r_count_4_io_out ? io_r_74_b : _GEN_3163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3165 = 10'h4b == r_count_4_io_out ? io_r_75_b : _GEN_3164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3166 = 10'h4c == r_count_4_io_out ? io_r_76_b : _GEN_3165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3167 = 10'h4d == r_count_4_io_out ? io_r_77_b : _GEN_3166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3168 = 10'h4e == r_count_4_io_out ? io_r_78_b : _GEN_3167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3169 = 10'h4f == r_count_4_io_out ? io_r_79_b : _GEN_3168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3170 = 10'h50 == r_count_4_io_out ? io_r_80_b : _GEN_3169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3171 = 10'h51 == r_count_4_io_out ? io_r_81_b : _GEN_3170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3172 = 10'h52 == r_count_4_io_out ? io_r_82_b : _GEN_3171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3173 = 10'h53 == r_count_4_io_out ? io_r_83_b : _GEN_3172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3174 = 10'h54 == r_count_4_io_out ? io_r_84_b : _GEN_3173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3175 = 10'h55 == r_count_4_io_out ? io_r_85_b : _GEN_3174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3176 = 10'h56 == r_count_4_io_out ? io_r_86_b : _GEN_3175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3177 = 10'h57 == r_count_4_io_out ? io_r_87_b : _GEN_3176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3178 = 10'h58 == r_count_4_io_out ? io_r_88_b : _GEN_3177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3179 = 10'h59 == r_count_4_io_out ? io_r_89_b : _GEN_3178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3180 = 10'h5a == r_count_4_io_out ? io_r_90_b : _GEN_3179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3181 = 10'h5b == r_count_4_io_out ? io_r_91_b : _GEN_3180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3182 = 10'h5c == r_count_4_io_out ? io_r_92_b : _GEN_3181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3183 = 10'h5d == r_count_4_io_out ? io_r_93_b : _GEN_3182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3184 = 10'h5e == r_count_4_io_out ? io_r_94_b : _GEN_3183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3185 = 10'h5f == r_count_4_io_out ? io_r_95_b : _GEN_3184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3186 = 10'h60 == r_count_4_io_out ? io_r_96_b : _GEN_3185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3187 = 10'h61 == r_count_4_io_out ? io_r_97_b : _GEN_3186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3188 = 10'h62 == r_count_4_io_out ? io_r_98_b : _GEN_3187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3189 = 10'h63 == r_count_4_io_out ? io_r_99_b : _GEN_3188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3190 = 10'h64 == r_count_4_io_out ? io_r_100_b : _GEN_3189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3191 = 10'h65 == r_count_4_io_out ? io_r_101_b : _GEN_3190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3192 = 10'h66 == r_count_4_io_out ? io_r_102_b : _GEN_3191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3193 = 10'h67 == r_count_4_io_out ? io_r_103_b : _GEN_3192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3194 = 10'h68 == r_count_4_io_out ? io_r_104_b : _GEN_3193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3195 = 10'h69 == r_count_4_io_out ? io_r_105_b : _GEN_3194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3196 = 10'h6a == r_count_4_io_out ? io_r_106_b : _GEN_3195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3197 = 10'h6b == r_count_4_io_out ? io_r_107_b : _GEN_3196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3198 = 10'h6c == r_count_4_io_out ? io_r_108_b : _GEN_3197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3199 = 10'h6d == r_count_4_io_out ? io_r_109_b : _GEN_3198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3200 = 10'h6e == r_count_4_io_out ? io_r_110_b : _GEN_3199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3201 = 10'h6f == r_count_4_io_out ? io_r_111_b : _GEN_3200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3202 = 10'h70 == r_count_4_io_out ? io_r_112_b : _GEN_3201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3203 = 10'h71 == r_count_4_io_out ? io_r_113_b : _GEN_3202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3204 = 10'h72 == r_count_4_io_out ? io_r_114_b : _GEN_3203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3205 = 10'h73 == r_count_4_io_out ? io_r_115_b : _GEN_3204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3206 = 10'h74 == r_count_4_io_out ? io_r_116_b : _GEN_3205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3207 = 10'h75 == r_count_4_io_out ? io_r_117_b : _GEN_3206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3208 = 10'h76 == r_count_4_io_out ? io_r_118_b : _GEN_3207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3209 = 10'h77 == r_count_4_io_out ? io_r_119_b : _GEN_3208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3210 = 10'h78 == r_count_4_io_out ? io_r_120_b : _GEN_3209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3211 = 10'h79 == r_count_4_io_out ? io_r_121_b : _GEN_3210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3212 = 10'h7a == r_count_4_io_out ? io_r_122_b : _GEN_3211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3213 = 10'h7b == r_count_4_io_out ? io_r_123_b : _GEN_3212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3214 = 10'h7c == r_count_4_io_out ? io_r_124_b : _GEN_3213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3215 = 10'h7d == r_count_4_io_out ? io_r_125_b : _GEN_3214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3216 = 10'h7e == r_count_4_io_out ? io_r_126_b : _GEN_3215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3217 = 10'h7f == r_count_4_io_out ? io_r_127_b : _GEN_3216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3218 = 10'h80 == r_count_4_io_out ? io_r_128_b : _GEN_3217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3219 = 10'h81 == r_count_4_io_out ? io_r_129_b : _GEN_3218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3220 = 10'h82 == r_count_4_io_out ? io_r_130_b : _GEN_3219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3221 = 10'h83 == r_count_4_io_out ? io_r_131_b : _GEN_3220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3222 = 10'h84 == r_count_4_io_out ? io_r_132_b : _GEN_3221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3223 = 10'h85 == r_count_4_io_out ? io_r_133_b : _GEN_3222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3224 = 10'h86 == r_count_4_io_out ? io_r_134_b : _GEN_3223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3225 = 10'h87 == r_count_4_io_out ? io_r_135_b : _GEN_3224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3226 = 10'h88 == r_count_4_io_out ? io_r_136_b : _GEN_3225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3227 = 10'h89 == r_count_4_io_out ? io_r_137_b : _GEN_3226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3228 = 10'h8a == r_count_4_io_out ? io_r_138_b : _GEN_3227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3229 = 10'h8b == r_count_4_io_out ? io_r_139_b : _GEN_3228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3230 = 10'h8c == r_count_4_io_out ? io_r_140_b : _GEN_3229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3231 = 10'h8d == r_count_4_io_out ? io_r_141_b : _GEN_3230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3232 = 10'h8e == r_count_4_io_out ? io_r_142_b : _GEN_3231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3233 = 10'h8f == r_count_4_io_out ? io_r_143_b : _GEN_3232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3234 = 10'h90 == r_count_4_io_out ? io_r_144_b : _GEN_3233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3235 = 10'h91 == r_count_4_io_out ? io_r_145_b : _GEN_3234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3236 = 10'h92 == r_count_4_io_out ? io_r_146_b : _GEN_3235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3237 = 10'h93 == r_count_4_io_out ? io_r_147_b : _GEN_3236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3238 = 10'h94 == r_count_4_io_out ? io_r_148_b : _GEN_3237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3239 = 10'h95 == r_count_4_io_out ? io_r_149_b : _GEN_3238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3240 = 10'h96 == r_count_4_io_out ? io_r_150_b : _GEN_3239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3241 = 10'h97 == r_count_4_io_out ? io_r_151_b : _GEN_3240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3242 = 10'h98 == r_count_4_io_out ? io_r_152_b : _GEN_3241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3243 = 10'h99 == r_count_4_io_out ? io_r_153_b : _GEN_3242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3244 = 10'h9a == r_count_4_io_out ? io_r_154_b : _GEN_3243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3245 = 10'h9b == r_count_4_io_out ? io_r_155_b : _GEN_3244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3246 = 10'h9c == r_count_4_io_out ? io_r_156_b : _GEN_3245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3247 = 10'h9d == r_count_4_io_out ? io_r_157_b : _GEN_3246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3248 = 10'h9e == r_count_4_io_out ? io_r_158_b : _GEN_3247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3249 = 10'h9f == r_count_4_io_out ? io_r_159_b : _GEN_3248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3250 = 10'ha0 == r_count_4_io_out ? io_r_160_b : _GEN_3249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3251 = 10'ha1 == r_count_4_io_out ? io_r_161_b : _GEN_3250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3252 = 10'ha2 == r_count_4_io_out ? io_r_162_b : _GEN_3251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3253 = 10'ha3 == r_count_4_io_out ? io_r_163_b : _GEN_3252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3254 = 10'ha4 == r_count_4_io_out ? io_r_164_b : _GEN_3253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3255 = 10'ha5 == r_count_4_io_out ? io_r_165_b : _GEN_3254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3256 = 10'ha6 == r_count_4_io_out ? io_r_166_b : _GEN_3255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3257 = 10'ha7 == r_count_4_io_out ? io_r_167_b : _GEN_3256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3258 = 10'ha8 == r_count_4_io_out ? io_r_168_b : _GEN_3257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3259 = 10'ha9 == r_count_4_io_out ? io_r_169_b : _GEN_3258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3260 = 10'haa == r_count_4_io_out ? io_r_170_b : _GEN_3259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3261 = 10'hab == r_count_4_io_out ? io_r_171_b : _GEN_3260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3262 = 10'hac == r_count_4_io_out ? io_r_172_b : _GEN_3261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3263 = 10'had == r_count_4_io_out ? io_r_173_b : _GEN_3262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3264 = 10'hae == r_count_4_io_out ? io_r_174_b : _GEN_3263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3265 = 10'haf == r_count_4_io_out ? io_r_175_b : _GEN_3264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3266 = 10'hb0 == r_count_4_io_out ? io_r_176_b : _GEN_3265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3267 = 10'hb1 == r_count_4_io_out ? io_r_177_b : _GEN_3266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3268 = 10'hb2 == r_count_4_io_out ? io_r_178_b : _GEN_3267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3269 = 10'hb3 == r_count_4_io_out ? io_r_179_b : _GEN_3268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3270 = 10'hb4 == r_count_4_io_out ? io_r_180_b : _GEN_3269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3271 = 10'hb5 == r_count_4_io_out ? io_r_181_b : _GEN_3270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3272 = 10'hb6 == r_count_4_io_out ? io_r_182_b : _GEN_3271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3273 = 10'hb7 == r_count_4_io_out ? io_r_183_b : _GEN_3272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3274 = 10'hb8 == r_count_4_io_out ? io_r_184_b : _GEN_3273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3275 = 10'hb9 == r_count_4_io_out ? io_r_185_b : _GEN_3274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3276 = 10'hba == r_count_4_io_out ? io_r_186_b : _GEN_3275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3277 = 10'hbb == r_count_4_io_out ? io_r_187_b : _GEN_3276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3278 = 10'hbc == r_count_4_io_out ? io_r_188_b : _GEN_3277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3279 = 10'hbd == r_count_4_io_out ? io_r_189_b : _GEN_3278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3280 = 10'hbe == r_count_4_io_out ? io_r_190_b : _GEN_3279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3281 = 10'hbf == r_count_4_io_out ? io_r_191_b : _GEN_3280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3282 = 10'hc0 == r_count_4_io_out ? io_r_192_b : _GEN_3281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3283 = 10'hc1 == r_count_4_io_out ? io_r_193_b : _GEN_3282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3284 = 10'hc2 == r_count_4_io_out ? io_r_194_b : _GEN_3283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3285 = 10'hc3 == r_count_4_io_out ? io_r_195_b : _GEN_3284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3286 = 10'hc4 == r_count_4_io_out ? io_r_196_b : _GEN_3285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3287 = 10'hc5 == r_count_4_io_out ? io_r_197_b : _GEN_3286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3288 = 10'hc6 == r_count_4_io_out ? io_r_198_b : _GEN_3287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3289 = 10'hc7 == r_count_4_io_out ? io_r_199_b : _GEN_3288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3290 = 10'hc8 == r_count_4_io_out ? io_r_200_b : _GEN_3289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3291 = 10'hc9 == r_count_4_io_out ? io_r_201_b : _GEN_3290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3292 = 10'hca == r_count_4_io_out ? io_r_202_b : _GEN_3291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3293 = 10'hcb == r_count_4_io_out ? io_r_203_b : _GEN_3292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3294 = 10'hcc == r_count_4_io_out ? io_r_204_b : _GEN_3293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3295 = 10'hcd == r_count_4_io_out ? io_r_205_b : _GEN_3294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3296 = 10'hce == r_count_4_io_out ? io_r_206_b : _GEN_3295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3297 = 10'hcf == r_count_4_io_out ? io_r_207_b : _GEN_3296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3298 = 10'hd0 == r_count_4_io_out ? io_r_208_b : _GEN_3297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3299 = 10'hd1 == r_count_4_io_out ? io_r_209_b : _GEN_3298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3300 = 10'hd2 == r_count_4_io_out ? io_r_210_b : _GEN_3299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3301 = 10'hd3 == r_count_4_io_out ? io_r_211_b : _GEN_3300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3302 = 10'hd4 == r_count_4_io_out ? io_r_212_b : _GEN_3301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3303 = 10'hd5 == r_count_4_io_out ? io_r_213_b : _GEN_3302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3304 = 10'hd6 == r_count_4_io_out ? io_r_214_b : _GEN_3303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3305 = 10'hd7 == r_count_4_io_out ? io_r_215_b : _GEN_3304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3306 = 10'hd8 == r_count_4_io_out ? io_r_216_b : _GEN_3305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3307 = 10'hd9 == r_count_4_io_out ? io_r_217_b : _GEN_3306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3308 = 10'hda == r_count_4_io_out ? io_r_218_b : _GEN_3307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3309 = 10'hdb == r_count_4_io_out ? io_r_219_b : _GEN_3308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3310 = 10'hdc == r_count_4_io_out ? io_r_220_b : _GEN_3309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3311 = 10'hdd == r_count_4_io_out ? io_r_221_b : _GEN_3310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3312 = 10'hde == r_count_4_io_out ? io_r_222_b : _GEN_3311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3313 = 10'hdf == r_count_4_io_out ? io_r_223_b : _GEN_3312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3314 = 10'he0 == r_count_4_io_out ? io_r_224_b : _GEN_3313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3315 = 10'he1 == r_count_4_io_out ? io_r_225_b : _GEN_3314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3316 = 10'he2 == r_count_4_io_out ? io_r_226_b : _GEN_3315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3317 = 10'he3 == r_count_4_io_out ? io_r_227_b : _GEN_3316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3318 = 10'he4 == r_count_4_io_out ? io_r_228_b : _GEN_3317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3319 = 10'he5 == r_count_4_io_out ? io_r_229_b : _GEN_3318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3320 = 10'he6 == r_count_4_io_out ? io_r_230_b : _GEN_3319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3321 = 10'he7 == r_count_4_io_out ? io_r_231_b : _GEN_3320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3322 = 10'he8 == r_count_4_io_out ? io_r_232_b : _GEN_3321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3323 = 10'he9 == r_count_4_io_out ? io_r_233_b : _GEN_3322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3324 = 10'hea == r_count_4_io_out ? io_r_234_b : _GEN_3323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3325 = 10'heb == r_count_4_io_out ? io_r_235_b : _GEN_3324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3326 = 10'hec == r_count_4_io_out ? io_r_236_b : _GEN_3325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3327 = 10'hed == r_count_4_io_out ? io_r_237_b : _GEN_3326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3328 = 10'hee == r_count_4_io_out ? io_r_238_b : _GEN_3327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3329 = 10'hef == r_count_4_io_out ? io_r_239_b : _GEN_3328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3330 = 10'hf0 == r_count_4_io_out ? io_r_240_b : _GEN_3329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3331 = 10'hf1 == r_count_4_io_out ? io_r_241_b : _GEN_3330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3332 = 10'hf2 == r_count_4_io_out ? io_r_242_b : _GEN_3331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3333 = 10'hf3 == r_count_4_io_out ? io_r_243_b : _GEN_3332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3334 = 10'hf4 == r_count_4_io_out ? io_r_244_b : _GEN_3333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3335 = 10'hf5 == r_count_4_io_out ? io_r_245_b : _GEN_3334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3336 = 10'hf6 == r_count_4_io_out ? io_r_246_b : _GEN_3335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3337 = 10'hf7 == r_count_4_io_out ? io_r_247_b : _GEN_3336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3338 = 10'hf8 == r_count_4_io_out ? io_r_248_b : _GEN_3337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3339 = 10'hf9 == r_count_4_io_out ? io_r_249_b : _GEN_3338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3340 = 10'hfa == r_count_4_io_out ? io_r_250_b : _GEN_3339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3341 = 10'hfb == r_count_4_io_out ? io_r_251_b : _GEN_3340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3342 = 10'hfc == r_count_4_io_out ? io_r_252_b : _GEN_3341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3343 = 10'hfd == r_count_4_io_out ? io_r_253_b : _GEN_3342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3344 = 10'hfe == r_count_4_io_out ? io_r_254_b : _GEN_3343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3345 = 10'hff == r_count_4_io_out ? io_r_255_b : _GEN_3344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3346 = 10'h100 == r_count_4_io_out ? io_r_256_b : _GEN_3345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3347 = 10'h101 == r_count_4_io_out ? io_r_257_b : _GEN_3346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3348 = 10'h102 == r_count_4_io_out ? io_r_258_b : _GEN_3347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3349 = 10'h103 == r_count_4_io_out ? io_r_259_b : _GEN_3348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3350 = 10'h104 == r_count_4_io_out ? io_r_260_b : _GEN_3349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3351 = 10'h105 == r_count_4_io_out ? io_r_261_b : _GEN_3350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3352 = 10'h106 == r_count_4_io_out ? io_r_262_b : _GEN_3351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3353 = 10'h107 == r_count_4_io_out ? io_r_263_b : _GEN_3352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3354 = 10'h108 == r_count_4_io_out ? io_r_264_b : _GEN_3353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3355 = 10'h109 == r_count_4_io_out ? io_r_265_b : _GEN_3354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3356 = 10'h10a == r_count_4_io_out ? io_r_266_b : _GEN_3355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3357 = 10'h10b == r_count_4_io_out ? io_r_267_b : _GEN_3356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3358 = 10'h10c == r_count_4_io_out ? io_r_268_b : _GEN_3357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3359 = 10'h10d == r_count_4_io_out ? io_r_269_b : _GEN_3358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3360 = 10'h10e == r_count_4_io_out ? io_r_270_b : _GEN_3359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3361 = 10'h10f == r_count_4_io_out ? io_r_271_b : _GEN_3360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3362 = 10'h110 == r_count_4_io_out ? io_r_272_b : _GEN_3361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3363 = 10'h111 == r_count_4_io_out ? io_r_273_b : _GEN_3362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3364 = 10'h112 == r_count_4_io_out ? io_r_274_b : _GEN_3363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3365 = 10'h113 == r_count_4_io_out ? io_r_275_b : _GEN_3364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3366 = 10'h114 == r_count_4_io_out ? io_r_276_b : _GEN_3365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3367 = 10'h115 == r_count_4_io_out ? io_r_277_b : _GEN_3366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3368 = 10'h116 == r_count_4_io_out ? io_r_278_b : _GEN_3367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3369 = 10'h117 == r_count_4_io_out ? io_r_279_b : _GEN_3368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3370 = 10'h118 == r_count_4_io_out ? io_r_280_b : _GEN_3369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3371 = 10'h119 == r_count_4_io_out ? io_r_281_b : _GEN_3370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3372 = 10'h11a == r_count_4_io_out ? io_r_282_b : _GEN_3371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3373 = 10'h11b == r_count_4_io_out ? io_r_283_b : _GEN_3372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3374 = 10'h11c == r_count_4_io_out ? io_r_284_b : _GEN_3373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3375 = 10'h11d == r_count_4_io_out ? io_r_285_b : _GEN_3374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3376 = 10'h11e == r_count_4_io_out ? io_r_286_b : _GEN_3375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3377 = 10'h11f == r_count_4_io_out ? io_r_287_b : _GEN_3376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3378 = 10'h120 == r_count_4_io_out ? io_r_288_b : _GEN_3377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3379 = 10'h121 == r_count_4_io_out ? io_r_289_b : _GEN_3378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3380 = 10'h122 == r_count_4_io_out ? io_r_290_b : _GEN_3379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3381 = 10'h123 == r_count_4_io_out ? io_r_291_b : _GEN_3380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3382 = 10'h124 == r_count_4_io_out ? io_r_292_b : _GEN_3381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3383 = 10'h125 == r_count_4_io_out ? io_r_293_b : _GEN_3382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3384 = 10'h126 == r_count_4_io_out ? io_r_294_b : _GEN_3383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3385 = 10'h127 == r_count_4_io_out ? io_r_295_b : _GEN_3384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3386 = 10'h128 == r_count_4_io_out ? io_r_296_b : _GEN_3385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3387 = 10'h129 == r_count_4_io_out ? io_r_297_b : _GEN_3386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3388 = 10'h12a == r_count_4_io_out ? io_r_298_b : _GEN_3387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3389 = 10'h12b == r_count_4_io_out ? io_r_299_b : _GEN_3388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3390 = 10'h12c == r_count_4_io_out ? io_r_300_b : _GEN_3389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3391 = 10'h12d == r_count_4_io_out ? io_r_301_b : _GEN_3390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3392 = 10'h12e == r_count_4_io_out ? io_r_302_b : _GEN_3391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3393 = 10'h12f == r_count_4_io_out ? io_r_303_b : _GEN_3392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3394 = 10'h130 == r_count_4_io_out ? io_r_304_b : _GEN_3393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3395 = 10'h131 == r_count_4_io_out ? io_r_305_b : _GEN_3394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3396 = 10'h132 == r_count_4_io_out ? io_r_306_b : _GEN_3395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3397 = 10'h133 == r_count_4_io_out ? io_r_307_b : _GEN_3396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3398 = 10'h134 == r_count_4_io_out ? io_r_308_b : _GEN_3397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3399 = 10'h135 == r_count_4_io_out ? io_r_309_b : _GEN_3398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3400 = 10'h136 == r_count_4_io_out ? io_r_310_b : _GEN_3399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3401 = 10'h137 == r_count_4_io_out ? io_r_311_b : _GEN_3400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3402 = 10'h138 == r_count_4_io_out ? io_r_312_b : _GEN_3401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3403 = 10'h139 == r_count_4_io_out ? io_r_313_b : _GEN_3402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3404 = 10'h13a == r_count_4_io_out ? io_r_314_b : _GEN_3403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3405 = 10'h13b == r_count_4_io_out ? io_r_315_b : _GEN_3404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3406 = 10'h13c == r_count_4_io_out ? io_r_316_b : _GEN_3405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3407 = 10'h13d == r_count_4_io_out ? io_r_317_b : _GEN_3406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3408 = 10'h13e == r_count_4_io_out ? io_r_318_b : _GEN_3407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3409 = 10'h13f == r_count_4_io_out ? io_r_319_b : _GEN_3408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3410 = 10'h140 == r_count_4_io_out ? io_r_320_b : _GEN_3409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3411 = 10'h141 == r_count_4_io_out ? io_r_321_b : _GEN_3410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3412 = 10'h142 == r_count_4_io_out ? io_r_322_b : _GEN_3411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3413 = 10'h143 == r_count_4_io_out ? io_r_323_b : _GEN_3412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3414 = 10'h144 == r_count_4_io_out ? io_r_324_b : _GEN_3413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3415 = 10'h145 == r_count_4_io_out ? io_r_325_b : _GEN_3414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3416 = 10'h146 == r_count_4_io_out ? io_r_326_b : _GEN_3415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3417 = 10'h147 == r_count_4_io_out ? io_r_327_b : _GEN_3416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3418 = 10'h148 == r_count_4_io_out ? io_r_328_b : _GEN_3417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3419 = 10'h149 == r_count_4_io_out ? io_r_329_b : _GEN_3418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3420 = 10'h14a == r_count_4_io_out ? io_r_330_b : _GEN_3419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3421 = 10'h14b == r_count_4_io_out ? io_r_331_b : _GEN_3420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3422 = 10'h14c == r_count_4_io_out ? io_r_332_b : _GEN_3421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3423 = 10'h14d == r_count_4_io_out ? io_r_333_b : _GEN_3422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3424 = 10'h14e == r_count_4_io_out ? io_r_334_b : _GEN_3423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3425 = 10'h14f == r_count_4_io_out ? io_r_335_b : _GEN_3424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3426 = 10'h150 == r_count_4_io_out ? io_r_336_b : _GEN_3425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3427 = 10'h151 == r_count_4_io_out ? io_r_337_b : _GEN_3426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3428 = 10'h152 == r_count_4_io_out ? io_r_338_b : _GEN_3427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3429 = 10'h153 == r_count_4_io_out ? io_r_339_b : _GEN_3428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3430 = 10'h154 == r_count_4_io_out ? io_r_340_b : _GEN_3429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3431 = 10'h155 == r_count_4_io_out ? io_r_341_b : _GEN_3430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3432 = 10'h156 == r_count_4_io_out ? io_r_342_b : _GEN_3431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3433 = 10'h157 == r_count_4_io_out ? io_r_343_b : _GEN_3432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3434 = 10'h158 == r_count_4_io_out ? io_r_344_b : _GEN_3433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3435 = 10'h159 == r_count_4_io_out ? io_r_345_b : _GEN_3434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3436 = 10'h15a == r_count_4_io_out ? io_r_346_b : _GEN_3435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3437 = 10'h15b == r_count_4_io_out ? io_r_347_b : _GEN_3436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3438 = 10'h15c == r_count_4_io_out ? io_r_348_b : _GEN_3437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3439 = 10'h15d == r_count_4_io_out ? io_r_349_b : _GEN_3438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3440 = 10'h15e == r_count_4_io_out ? io_r_350_b : _GEN_3439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3441 = 10'h15f == r_count_4_io_out ? io_r_351_b : _GEN_3440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3442 = 10'h160 == r_count_4_io_out ? io_r_352_b : _GEN_3441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3443 = 10'h161 == r_count_4_io_out ? io_r_353_b : _GEN_3442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3444 = 10'h162 == r_count_4_io_out ? io_r_354_b : _GEN_3443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3445 = 10'h163 == r_count_4_io_out ? io_r_355_b : _GEN_3444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3446 = 10'h164 == r_count_4_io_out ? io_r_356_b : _GEN_3445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3447 = 10'h165 == r_count_4_io_out ? io_r_357_b : _GEN_3446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3448 = 10'h166 == r_count_4_io_out ? io_r_358_b : _GEN_3447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3449 = 10'h167 == r_count_4_io_out ? io_r_359_b : _GEN_3448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3450 = 10'h168 == r_count_4_io_out ? io_r_360_b : _GEN_3449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3451 = 10'h169 == r_count_4_io_out ? io_r_361_b : _GEN_3450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3452 = 10'h16a == r_count_4_io_out ? io_r_362_b : _GEN_3451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3453 = 10'h16b == r_count_4_io_out ? io_r_363_b : _GEN_3452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3454 = 10'h16c == r_count_4_io_out ? io_r_364_b : _GEN_3453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3455 = 10'h16d == r_count_4_io_out ? io_r_365_b : _GEN_3454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3456 = 10'h16e == r_count_4_io_out ? io_r_366_b : _GEN_3455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3457 = 10'h16f == r_count_4_io_out ? io_r_367_b : _GEN_3456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3458 = 10'h170 == r_count_4_io_out ? io_r_368_b : _GEN_3457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3459 = 10'h171 == r_count_4_io_out ? io_r_369_b : _GEN_3458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3460 = 10'h172 == r_count_4_io_out ? io_r_370_b : _GEN_3459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3461 = 10'h173 == r_count_4_io_out ? io_r_371_b : _GEN_3460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3462 = 10'h174 == r_count_4_io_out ? io_r_372_b : _GEN_3461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3463 = 10'h175 == r_count_4_io_out ? io_r_373_b : _GEN_3462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3464 = 10'h176 == r_count_4_io_out ? io_r_374_b : _GEN_3463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3465 = 10'h177 == r_count_4_io_out ? io_r_375_b : _GEN_3464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3466 = 10'h178 == r_count_4_io_out ? io_r_376_b : _GEN_3465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3467 = 10'h179 == r_count_4_io_out ? io_r_377_b : _GEN_3466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3468 = 10'h17a == r_count_4_io_out ? io_r_378_b : _GEN_3467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3469 = 10'h17b == r_count_4_io_out ? io_r_379_b : _GEN_3468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3470 = 10'h17c == r_count_4_io_out ? io_r_380_b : _GEN_3469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3471 = 10'h17d == r_count_4_io_out ? io_r_381_b : _GEN_3470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3472 = 10'h17e == r_count_4_io_out ? io_r_382_b : _GEN_3471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3473 = 10'h17f == r_count_4_io_out ? io_r_383_b : _GEN_3472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3474 = 10'h180 == r_count_4_io_out ? io_r_384_b : _GEN_3473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3475 = 10'h181 == r_count_4_io_out ? io_r_385_b : _GEN_3474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3476 = 10'h182 == r_count_4_io_out ? io_r_386_b : _GEN_3475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3477 = 10'h183 == r_count_4_io_out ? io_r_387_b : _GEN_3476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3478 = 10'h184 == r_count_4_io_out ? io_r_388_b : _GEN_3477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3479 = 10'h185 == r_count_4_io_out ? io_r_389_b : _GEN_3478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3480 = 10'h186 == r_count_4_io_out ? io_r_390_b : _GEN_3479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3481 = 10'h187 == r_count_4_io_out ? io_r_391_b : _GEN_3480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3482 = 10'h188 == r_count_4_io_out ? io_r_392_b : _GEN_3481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3483 = 10'h189 == r_count_4_io_out ? io_r_393_b : _GEN_3482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3484 = 10'h18a == r_count_4_io_out ? io_r_394_b : _GEN_3483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3485 = 10'h18b == r_count_4_io_out ? io_r_395_b : _GEN_3484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3486 = 10'h18c == r_count_4_io_out ? io_r_396_b : _GEN_3485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3487 = 10'h18d == r_count_4_io_out ? io_r_397_b : _GEN_3486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3488 = 10'h18e == r_count_4_io_out ? io_r_398_b : _GEN_3487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3489 = 10'h18f == r_count_4_io_out ? io_r_399_b : _GEN_3488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3490 = 10'h190 == r_count_4_io_out ? io_r_400_b : _GEN_3489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3491 = 10'h191 == r_count_4_io_out ? io_r_401_b : _GEN_3490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3492 = 10'h192 == r_count_4_io_out ? io_r_402_b : _GEN_3491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3493 = 10'h193 == r_count_4_io_out ? io_r_403_b : _GEN_3492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3494 = 10'h194 == r_count_4_io_out ? io_r_404_b : _GEN_3493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3495 = 10'h195 == r_count_4_io_out ? io_r_405_b : _GEN_3494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3496 = 10'h196 == r_count_4_io_out ? io_r_406_b : _GEN_3495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3497 = 10'h197 == r_count_4_io_out ? io_r_407_b : _GEN_3496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3498 = 10'h198 == r_count_4_io_out ? io_r_408_b : _GEN_3497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3499 = 10'h199 == r_count_4_io_out ? io_r_409_b : _GEN_3498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3500 = 10'h19a == r_count_4_io_out ? io_r_410_b : _GEN_3499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3501 = 10'h19b == r_count_4_io_out ? io_r_411_b : _GEN_3500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3502 = 10'h19c == r_count_4_io_out ? io_r_412_b : _GEN_3501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3503 = 10'h19d == r_count_4_io_out ? io_r_413_b : _GEN_3502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3504 = 10'h19e == r_count_4_io_out ? io_r_414_b : _GEN_3503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3505 = 10'h19f == r_count_4_io_out ? io_r_415_b : _GEN_3504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3506 = 10'h1a0 == r_count_4_io_out ? io_r_416_b : _GEN_3505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3507 = 10'h1a1 == r_count_4_io_out ? io_r_417_b : _GEN_3506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3508 = 10'h1a2 == r_count_4_io_out ? io_r_418_b : _GEN_3507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3509 = 10'h1a3 == r_count_4_io_out ? io_r_419_b : _GEN_3508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3510 = 10'h1a4 == r_count_4_io_out ? io_r_420_b : _GEN_3509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3511 = 10'h1a5 == r_count_4_io_out ? io_r_421_b : _GEN_3510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3512 = 10'h1a6 == r_count_4_io_out ? io_r_422_b : _GEN_3511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3513 = 10'h1a7 == r_count_4_io_out ? io_r_423_b : _GEN_3512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3514 = 10'h1a8 == r_count_4_io_out ? io_r_424_b : _GEN_3513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3515 = 10'h1a9 == r_count_4_io_out ? io_r_425_b : _GEN_3514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3516 = 10'h1aa == r_count_4_io_out ? io_r_426_b : _GEN_3515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3517 = 10'h1ab == r_count_4_io_out ? io_r_427_b : _GEN_3516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3518 = 10'h1ac == r_count_4_io_out ? io_r_428_b : _GEN_3517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3519 = 10'h1ad == r_count_4_io_out ? io_r_429_b : _GEN_3518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3520 = 10'h1ae == r_count_4_io_out ? io_r_430_b : _GEN_3519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3521 = 10'h1af == r_count_4_io_out ? io_r_431_b : _GEN_3520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3522 = 10'h1b0 == r_count_4_io_out ? io_r_432_b : _GEN_3521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3523 = 10'h1b1 == r_count_4_io_out ? io_r_433_b : _GEN_3522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3524 = 10'h1b2 == r_count_4_io_out ? io_r_434_b : _GEN_3523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3525 = 10'h1b3 == r_count_4_io_out ? io_r_435_b : _GEN_3524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3526 = 10'h1b4 == r_count_4_io_out ? io_r_436_b : _GEN_3525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3527 = 10'h1b5 == r_count_4_io_out ? io_r_437_b : _GEN_3526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3528 = 10'h1b6 == r_count_4_io_out ? io_r_438_b : _GEN_3527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3529 = 10'h1b7 == r_count_4_io_out ? io_r_439_b : _GEN_3528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3530 = 10'h1b8 == r_count_4_io_out ? io_r_440_b : _GEN_3529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3531 = 10'h1b9 == r_count_4_io_out ? io_r_441_b : _GEN_3530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3532 = 10'h1ba == r_count_4_io_out ? io_r_442_b : _GEN_3531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3533 = 10'h1bb == r_count_4_io_out ? io_r_443_b : _GEN_3532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3534 = 10'h1bc == r_count_4_io_out ? io_r_444_b : _GEN_3533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3535 = 10'h1bd == r_count_4_io_out ? io_r_445_b : _GEN_3534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3536 = 10'h1be == r_count_4_io_out ? io_r_446_b : _GEN_3535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3537 = 10'h1bf == r_count_4_io_out ? io_r_447_b : _GEN_3536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3538 = 10'h1c0 == r_count_4_io_out ? io_r_448_b : _GEN_3537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3539 = 10'h1c1 == r_count_4_io_out ? io_r_449_b : _GEN_3538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3540 = 10'h1c2 == r_count_4_io_out ? io_r_450_b : _GEN_3539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3541 = 10'h1c3 == r_count_4_io_out ? io_r_451_b : _GEN_3540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3542 = 10'h1c4 == r_count_4_io_out ? io_r_452_b : _GEN_3541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3543 = 10'h1c5 == r_count_4_io_out ? io_r_453_b : _GEN_3542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3544 = 10'h1c6 == r_count_4_io_out ? io_r_454_b : _GEN_3543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3545 = 10'h1c7 == r_count_4_io_out ? io_r_455_b : _GEN_3544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3546 = 10'h1c8 == r_count_4_io_out ? io_r_456_b : _GEN_3545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3547 = 10'h1c9 == r_count_4_io_out ? io_r_457_b : _GEN_3546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3548 = 10'h1ca == r_count_4_io_out ? io_r_458_b : _GEN_3547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3549 = 10'h1cb == r_count_4_io_out ? io_r_459_b : _GEN_3548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3550 = 10'h1cc == r_count_4_io_out ? io_r_460_b : _GEN_3549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3551 = 10'h1cd == r_count_4_io_out ? io_r_461_b : _GEN_3550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3552 = 10'h1ce == r_count_4_io_out ? io_r_462_b : _GEN_3551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3553 = 10'h1cf == r_count_4_io_out ? io_r_463_b : _GEN_3552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3554 = 10'h1d0 == r_count_4_io_out ? io_r_464_b : _GEN_3553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3555 = 10'h1d1 == r_count_4_io_out ? io_r_465_b : _GEN_3554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3556 = 10'h1d2 == r_count_4_io_out ? io_r_466_b : _GEN_3555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3557 = 10'h1d3 == r_count_4_io_out ? io_r_467_b : _GEN_3556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3558 = 10'h1d4 == r_count_4_io_out ? io_r_468_b : _GEN_3557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3559 = 10'h1d5 == r_count_4_io_out ? io_r_469_b : _GEN_3558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3560 = 10'h1d6 == r_count_4_io_out ? io_r_470_b : _GEN_3559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3561 = 10'h1d7 == r_count_4_io_out ? io_r_471_b : _GEN_3560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3562 = 10'h1d8 == r_count_4_io_out ? io_r_472_b : _GEN_3561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3563 = 10'h1d9 == r_count_4_io_out ? io_r_473_b : _GEN_3562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3564 = 10'h1da == r_count_4_io_out ? io_r_474_b : _GEN_3563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3565 = 10'h1db == r_count_4_io_out ? io_r_475_b : _GEN_3564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3566 = 10'h1dc == r_count_4_io_out ? io_r_476_b : _GEN_3565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3567 = 10'h1dd == r_count_4_io_out ? io_r_477_b : _GEN_3566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3568 = 10'h1de == r_count_4_io_out ? io_r_478_b : _GEN_3567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3569 = 10'h1df == r_count_4_io_out ? io_r_479_b : _GEN_3568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3570 = 10'h1e0 == r_count_4_io_out ? io_r_480_b : _GEN_3569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3571 = 10'h1e1 == r_count_4_io_out ? io_r_481_b : _GEN_3570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3572 = 10'h1e2 == r_count_4_io_out ? io_r_482_b : _GEN_3571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3573 = 10'h1e3 == r_count_4_io_out ? io_r_483_b : _GEN_3572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3574 = 10'h1e4 == r_count_4_io_out ? io_r_484_b : _GEN_3573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3575 = 10'h1e5 == r_count_4_io_out ? io_r_485_b : _GEN_3574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3576 = 10'h1e6 == r_count_4_io_out ? io_r_486_b : _GEN_3575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3577 = 10'h1e7 == r_count_4_io_out ? io_r_487_b : _GEN_3576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3578 = 10'h1e8 == r_count_4_io_out ? io_r_488_b : _GEN_3577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3579 = 10'h1e9 == r_count_4_io_out ? io_r_489_b : _GEN_3578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3580 = 10'h1ea == r_count_4_io_out ? io_r_490_b : _GEN_3579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3581 = 10'h1eb == r_count_4_io_out ? io_r_491_b : _GEN_3580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3582 = 10'h1ec == r_count_4_io_out ? io_r_492_b : _GEN_3581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3583 = 10'h1ed == r_count_4_io_out ? io_r_493_b : _GEN_3582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3584 = 10'h1ee == r_count_4_io_out ? io_r_494_b : _GEN_3583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3585 = 10'h1ef == r_count_4_io_out ? io_r_495_b : _GEN_3584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3586 = 10'h1f0 == r_count_4_io_out ? io_r_496_b : _GEN_3585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3587 = 10'h1f1 == r_count_4_io_out ? io_r_497_b : _GEN_3586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3588 = 10'h1f2 == r_count_4_io_out ? io_r_498_b : _GEN_3587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3589 = 10'h1f3 == r_count_4_io_out ? io_r_499_b : _GEN_3588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3590 = 10'h1f4 == r_count_4_io_out ? io_r_500_b : _GEN_3589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3591 = 10'h1f5 == r_count_4_io_out ? io_r_501_b : _GEN_3590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3592 = 10'h1f6 == r_count_4_io_out ? io_r_502_b : _GEN_3591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3593 = 10'h1f7 == r_count_4_io_out ? io_r_503_b : _GEN_3592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3594 = 10'h1f8 == r_count_4_io_out ? io_r_504_b : _GEN_3593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3595 = 10'h1f9 == r_count_4_io_out ? io_r_505_b : _GEN_3594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3596 = 10'h1fa == r_count_4_io_out ? io_r_506_b : _GEN_3595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3597 = 10'h1fb == r_count_4_io_out ? io_r_507_b : _GEN_3596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3598 = 10'h1fc == r_count_4_io_out ? io_r_508_b : _GEN_3597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3599 = 10'h1fd == r_count_4_io_out ? io_r_509_b : _GEN_3598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3600 = 10'h1fe == r_count_4_io_out ? io_r_510_b : _GEN_3599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3601 = 10'h1ff == r_count_4_io_out ? io_r_511_b : _GEN_3600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3602 = 10'h200 == r_count_4_io_out ? io_r_512_b : _GEN_3601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3603 = 10'h201 == r_count_4_io_out ? io_r_513_b : _GEN_3602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3604 = 10'h202 == r_count_4_io_out ? io_r_514_b : _GEN_3603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3605 = 10'h203 == r_count_4_io_out ? io_r_515_b : _GEN_3604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3606 = 10'h204 == r_count_4_io_out ? io_r_516_b : _GEN_3605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3607 = 10'h205 == r_count_4_io_out ? io_r_517_b : _GEN_3606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3608 = 10'h206 == r_count_4_io_out ? io_r_518_b : _GEN_3607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3609 = 10'h207 == r_count_4_io_out ? io_r_519_b : _GEN_3608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3610 = 10'h208 == r_count_4_io_out ? io_r_520_b : _GEN_3609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3611 = 10'h209 == r_count_4_io_out ? io_r_521_b : _GEN_3610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3612 = 10'h20a == r_count_4_io_out ? io_r_522_b : _GEN_3611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3613 = 10'h20b == r_count_4_io_out ? io_r_523_b : _GEN_3612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3614 = 10'h20c == r_count_4_io_out ? io_r_524_b : _GEN_3613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3615 = 10'h20d == r_count_4_io_out ? io_r_525_b : _GEN_3614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3616 = 10'h20e == r_count_4_io_out ? io_r_526_b : _GEN_3615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3617 = 10'h20f == r_count_4_io_out ? io_r_527_b : _GEN_3616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3618 = 10'h210 == r_count_4_io_out ? io_r_528_b : _GEN_3617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3619 = 10'h211 == r_count_4_io_out ? io_r_529_b : _GEN_3618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3620 = 10'h212 == r_count_4_io_out ? io_r_530_b : _GEN_3619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3621 = 10'h213 == r_count_4_io_out ? io_r_531_b : _GEN_3620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3622 = 10'h214 == r_count_4_io_out ? io_r_532_b : _GEN_3621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3623 = 10'h215 == r_count_4_io_out ? io_r_533_b : _GEN_3622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3624 = 10'h216 == r_count_4_io_out ? io_r_534_b : _GEN_3623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3625 = 10'h217 == r_count_4_io_out ? io_r_535_b : _GEN_3624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3626 = 10'h218 == r_count_4_io_out ? io_r_536_b : _GEN_3625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3627 = 10'h219 == r_count_4_io_out ? io_r_537_b : _GEN_3626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3628 = 10'h21a == r_count_4_io_out ? io_r_538_b : _GEN_3627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3629 = 10'h21b == r_count_4_io_out ? io_r_539_b : _GEN_3628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3630 = 10'h21c == r_count_4_io_out ? io_r_540_b : _GEN_3629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3631 = 10'h21d == r_count_4_io_out ? io_r_541_b : _GEN_3630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3632 = 10'h21e == r_count_4_io_out ? io_r_542_b : _GEN_3631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3633 = 10'h21f == r_count_4_io_out ? io_r_543_b : _GEN_3632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3634 = 10'h220 == r_count_4_io_out ? io_r_544_b : _GEN_3633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3635 = 10'h221 == r_count_4_io_out ? io_r_545_b : _GEN_3634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3636 = 10'h222 == r_count_4_io_out ? io_r_546_b : _GEN_3635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3637 = 10'h223 == r_count_4_io_out ? io_r_547_b : _GEN_3636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3638 = 10'h224 == r_count_4_io_out ? io_r_548_b : _GEN_3637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3639 = 10'h225 == r_count_4_io_out ? io_r_549_b : _GEN_3638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3640 = 10'h226 == r_count_4_io_out ? io_r_550_b : _GEN_3639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3641 = 10'h227 == r_count_4_io_out ? io_r_551_b : _GEN_3640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3642 = 10'h228 == r_count_4_io_out ? io_r_552_b : _GEN_3641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3643 = 10'h229 == r_count_4_io_out ? io_r_553_b : _GEN_3642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3644 = 10'h22a == r_count_4_io_out ? io_r_554_b : _GEN_3643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3645 = 10'h22b == r_count_4_io_out ? io_r_555_b : _GEN_3644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3646 = 10'h22c == r_count_4_io_out ? io_r_556_b : _GEN_3645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3647 = 10'h22d == r_count_4_io_out ? io_r_557_b : _GEN_3646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3648 = 10'h22e == r_count_4_io_out ? io_r_558_b : _GEN_3647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3649 = 10'h22f == r_count_4_io_out ? io_r_559_b : _GEN_3648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3650 = 10'h230 == r_count_4_io_out ? io_r_560_b : _GEN_3649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3651 = 10'h231 == r_count_4_io_out ? io_r_561_b : _GEN_3650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3652 = 10'h232 == r_count_4_io_out ? io_r_562_b : _GEN_3651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3653 = 10'h233 == r_count_4_io_out ? io_r_563_b : _GEN_3652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3654 = 10'h234 == r_count_4_io_out ? io_r_564_b : _GEN_3653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3655 = 10'h235 == r_count_4_io_out ? io_r_565_b : _GEN_3654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3656 = 10'h236 == r_count_4_io_out ? io_r_566_b : _GEN_3655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3657 = 10'h237 == r_count_4_io_out ? io_r_567_b : _GEN_3656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3658 = 10'h238 == r_count_4_io_out ? io_r_568_b : _GEN_3657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3659 = 10'h239 == r_count_4_io_out ? io_r_569_b : _GEN_3658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3660 = 10'h23a == r_count_4_io_out ? io_r_570_b : _GEN_3659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3661 = 10'h23b == r_count_4_io_out ? io_r_571_b : _GEN_3660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3662 = 10'h23c == r_count_4_io_out ? io_r_572_b : _GEN_3661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3663 = 10'h23d == r_count_4_io_out ? io_r_573_b : _GEN_3662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3664 = 10'h23e == r_count_4_io_out ? io_r_574_b : _GEN_3663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3665 = 10'h23f == r_count_4_io_out ? io_r_575_b : _GEN_3664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3666 = 10'h240 == r_count_4_io_out ? io_r_576_b : _GEN_3665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3667 = 10'h241 == r_count_4_io_out ? io_r_577_b : _GEN_3666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3668 = 10'h242 == r_count_4_io_out ? io_r_578_b : _GEN_3667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3669 = 10'h243 == r_count_4_io_out ? io_r_579_b : _GEN_3668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3670 = 10'h244 == r_count_4_io_out ? io_r_580_b : _GEN_3669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3671 = 10'h245 == r_count_4_io_out ? io_r_581_b : _GEN_3670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3672 = 10'h246 == r_count_4_io_out ? io_r_582_b : _GEN_3671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3673 = 10'h247 == r_count_4_io_out ? io_r_583_b : _GEN_3672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3674 = 10'h248 == r_count_4_io_out ? io_r_584_b : _GEN_3673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3675 = 10'h249 == r_count_4_io_out ? io_r_585_b : _GEN_3674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3676 = 10'h24a == r_count_4_io_out ? io_r_586_b : _GEN_3675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3677 = 10'h24b == r_count_4_io_out ? io_r_587_b : _GEN_3676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3678 = 10'h24c == r_count_4_io_out ? io_r_588_b : _GEN_3677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3679 = 10'h24d == r_count_4_io_out ? io_r_589_b : _GEN_3678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3680 = 10'h24e == r_count_4_io_out ? io_r_590_b : _GEN_3679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3681 = 10'h24f == r_count_4_io_out ? io_r_591_b : _GEN_3680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3682 = 10'h250 == r_count_4_io_out ? io_r_592_b : _GEN_3681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3683 = 10'h251 == r_count_4_io_out ? io_r_593_b : _GEN_3682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3684 = 10'h252 == r_count_4_io_out ? io_r_594_b : _GEN_3683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3685 = 10'h253 == r_count_4_io_out ? io_r_595_b : _GEN_3684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3686 = 10'h254 == r_count_4_io_out ? io_r_596_b : _GEN_3685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3687 = 10'h255 == r_count_4_io_out ? io_r_597_b : _GEN_3686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3688 = 10'h256 == r_count_4_io_out ? io_r_598_b : _GEN_3687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3689 = 10'h257 == r_count_4_io_out ? io_r_599_b : _GEN_3688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3690 = 10'h258 == r_count_4_io_out ? io_r_600_b : _GEN_3689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3691 = 10'h259 == r_count_4_io_out ? io_r_601_b : _GEN_3690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3692 = 10'h25a == r_count_4_io_out ? io_r_602_b : _GEN_3691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3693 = 10'h25b == r_count_4_io_out ? io_r_603_b : _GEN_3692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3694 = 10'h25c == r_count_4_io_out ? io_r_604_b : _GEN_3693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3695 = 10'h25d == r_count_4_io_out ? io_r_605_b : _GEN_3694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3696 = 10'h25e == r_count_4_io_out ? io_r_606_b : _GEN_3695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3697 = 10'h25f == r_count_4_io_out ? io_r_607_b : _GEN_3696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3698 = 10'h260 == r_count_4_io_out ? io_r_608_b : _GEN_3697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3699 = 10'h261 == r_count_4_io_out ? io_r_609_b : _GEN_3698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3700 = 10'h262 == r_count_4_io_out ? io_r_610_b : _GEN_3699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3701 = 10'h263 == r_count_4_io_out ? io_r_611_b : _GEN_3700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3702 = 10'h264 == r_count_4_io_out ? io_r_612_b : _GEN_3701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3703 = 10'h265 == r_count_4_io_out ? io_r_613_b : _GEN_3702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3704 = 10'h266 == r_count_4_io_out ? io_r_614_b : _GEN_3703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3705 = 10'h267 == r_count_4_io_out ? io_r_615_b : _GEN_3704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3706 = 10'h268 == r_count_4_io_out ? io_r_616_b : _GEN_3705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3707 = 10'h269 == r_count_4_io_out ? io_r_617_b : _GEN_3706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3708 = 10'h26a == r_count_4_io_out ? io_r_618_b : _GEN_3707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3709 = 10'h26b == r_count_4_io_out ? io_r_619_b : _GEN_3708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3710 = 10'h26c == r_count_4_io_out ? io_r_620_b : _GEN_3709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3711 = 10'h26d == r_count_4_io_out ? io_r_621_b : _GEN_3710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3712 = 10'h26e == r_count_4_io_out ? io_r_622_b : _GEN_3711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3713 = 10'h26f == r_count_4_io_out ? io_r_623_b : _GEN_3712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3714 = 10'h270 == r_count_4_io_out ? io_r_624_b : _GEN_3713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3715 = 10'h271 == r_count_4_io_out ? io_r_625_b : _GEN_3714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3716 = 10'h272 == r_count_4_io_out ? io_r_626_b : _GEN_3715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3717 = 10'h273 == r_count_4_io_out ? io_r_627_b : _GEN_3716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3718 = 10'h274 == r_count_4_io_out ? io_r_628_b : _GEN_3717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3719 = 10'h275 == r_count_4_io_out ? io_r_629_b : _GEN_3718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3720 = 10'h276 == r_count_4_io_out ? io_r_630_b : _GEN_3719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3721 = 10'h277 == r_count_4_io_out ? io_r_631_b : _GEN_3720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3722 = 10'h278 == r_count_4_io_out ? io_r_632_b : _GEN_3721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3723 = 10'h279 == r_count_4_io_out ? io_r_633_b : _GEN_3722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3724 = 10'h27a == r_count_4_io_out ? io_r_634_b : _GEN_3723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3725 = 10'h27b == r_count_4_io_out ? io_r_635_b : _GEN_3724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3726 = 10'h27c == r_count_4_io_out ? io_r_636_b : _GEN_3725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3727 = 10'h27d == r_count_4_io_out ? io_r_637_b : _GEN_3726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3728 = 10'h27e == r_count_4_io_out ? io_r_638_b : _GEN_3727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3729 = 10'h27f == r_count_4_io_out ? io_r_639_b : _GEN_3728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3730 = 10'h280 == r_count_4_io_out ? io_r_640_b : _GEN_3729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3731 = 10'h281 == r_count_4_io_out ? io_r_641_b : _GEN_3730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3732 = 10'h282 == r_count_4_io_out ? io_r_642_b : _GEN_3731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3733 = 10'h283 == r_count_4_io_out ? io_r_643_b : _GEN_3732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3734 = 10'h284 == r_count_4_io_out ? io_r_644_b : _GEN_3733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3735 = 10'h285 == r_count_4_io_out ? io_r_645_b : _GEN_3734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3736 = 10'h286 == r_count_4_io_out ? io_r_646_b : _GEN_3735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3737 = 10'h287 == r_count_4_io_out ? io_r_647_b : _GEN_3736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3738 = 10'h288 == r_count_4_io_out ? io_r_648_b : _GEN_3737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3739 = 10'h289 == r_count_4_io_out ? io_r_649_b : _GEN_3738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3740 = 10'h28a == r_count_4_io_out ? io_r_650_b : _GEN_3739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3741 = 10'h28b == r_count_4_io_out ? io_r_651_b : _GEN_3740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3742 = 10'h28c == r_count_4_io_out ? io_r_652_b : _GEN_3741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3743 = 10'h28d == r_count_4_io_out ? io_r_653_b : _GEN_3742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3744 = 10'h28e == r_count_4_io_out ? io_r_654_b : _GEN_3743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3745 = 10'h28f == r_count_4_io_out ? io_r_655_b : _GEN_3744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3746 = 10'h290 == r_count_4_io_out ? io_r_656_b : _GEN_3745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3747 = 10'h291 == r_count_4_io_out ? io_r_657_b : _GEN_3746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3748 = 10'h292 == r_count_4_io_out ? io_r_658_b : _GEN_3747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3749 = 10'h293 == r_count_4_io_out ? io_r_659_b : _GEN_3748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3750 = 10'h294 == r_count_4_io_out ? io_r_660_b : _GEN_3749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3751 = 10'h295 == r_count_4_io_out ? io_r_661_b : _GEN_3750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3752 = 10'h296 == r_count_4_io_out ? io_r_662_b : _GEN_3751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3753 = 10'h297 == r_count_4_io_out ? io_r_663_b : _GEN_3752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3754 = 10'h298 == r_count_4_io_out ? io_r_664_b : _GEN_3753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3755 = 10'h299 == r_count_4_io_out ? io_r_665_b : _GEN_3754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3756 = 10'h29a == r_count_4_io_out ? io_r_666_b : _GEN_3755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3757 = 10'h29b == r_count_4_io_out ? io_r_667_b : _GEN_3756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3758 = 10'h29c == r_count_4_io_out ? io_r_668_b : _GEN_3757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3759 = 10'h29d == r_count_4_io_out ? io_r_669_b : _GEN_3758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3760 = 10'h29e == r_count_4_io_out ? io_r_670_b : _GEN_3759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3761 = 10'h29f == r_count_4_io_out ? io_r_671_b : _GEN_3760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3762 = 10'h2a0 == r_count_4_io_out ? io_r_672_b : _GEN_3761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3763 = 10'h2a1 == r_count_4_io_out ? io_r_673_b : _GEN_3762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3764 = 10'h2a2 == r_count_4_io_out ? io_r_674_b : _GEN_3763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3765 = 10'h2a3 == r_count_4_io_out ? io_r_675_b : _GEN_3764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3766 = 10'h2a4 == r_count_4_io_out ? io_r_676_b : _GEN_3765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3767 = 10'h2a5 == r_count_4_io_out ? io_r_677_b : _GEN_3766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3768 = 10'h2a6 == r_count_4_io_out ? io_r_678_b : _GEN_3767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3769 = 10'h2a7 == r_count_4_io_out ? io_r_679_b : _GEN_3768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3770 = 10'h2a8 == r_count_4_io_out ? io_r_680_b : _GEN_3769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3771 = 10'h2a9 == r_count_4_io_out ? io_r_681_b : _GEN_3770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3772 = 10'h2aa == r_count_4_io_out ? io_r_682_b : _GEN_3771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3773 = 10'h2ab == r_count_4_io_out ? io_r_683_b : _GEN_3772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3774 = 10'h2ac == r_count_4_io_out ? io_r_684_b : _GEN_3773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3775 = 10'h2ad == r_count_4_io_out ? io_r_685_b : _GEN_3774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3776 = 10'h2ae == r_count_4_io_out ? io_r_686_b : _GEN_3775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3777 = 10'h2af == r_count_4_io_out ? io_r_687_b : _GEN_3776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3778 = 10'h2b0 == r_count_4_io_out ? io_r_688_b : _GEN_3777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3779 = 10'h2b1 == r_count_4_io_out ? io_r_689_b : _GEN_3778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3780 = 10'h2b2 == r_count_4_io_out ? io_r_690_b : _GEN_3779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3781 = 10'h2b3 == r_count_4_io_out ? io_r_691_b : _GEN_3780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3782 = 10'h2b4 == r_count_4_io_out ? io_r_692_b : _GEN_3781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3783 = 10'h2b5 == r_count_4_io_out ? io_r_693_b : _GEN_3782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3784 = 10'h2b6 == r_count_4_io_out ? io_r_694_b : _GEN_3783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3785 = 10'h2b7 == r_count_4_io_out ? io_r_695_b : _GEN_3784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3786 = 10'h2b8 == r_count_4_io_out ? io_r_696_b : _GEN_3785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3787 = 10'h2b9 == r_count_4_io_out ? io_r_697_b : _GEN_3786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3788 = 10'h2ba == r_count_4_io_out ? io_r_698_b : _GEN_3787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3789 = 10'h2bb == r_count_4_io_out ? io_r_699_b : _GEN_3788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3790 = 10'h2bc == r_count_4_io_out ? io_r_700_b : _GEN_3789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3791 = 10'h2bd == r_count_4_io_out ? io_r_701_b : _GEN_3790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3792 = 10'h2be == r_count_4_io_out ? io_r_702_b : _GEN_3791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3793 = 10'h2bf == r_count_4_io_out ? io_r_703_b : _GEN_3792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3794 = 10'h2c0 == r_count_4_io_out ? io_r_704_b : _GEN_3793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3795 = 10'h2c1 == r_count_4_io_out ? io_r_705_b : _GEN_3794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3796 = 10'h2c2 == r_count_4_io_out ? io_r_706_b : _GEN_3795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3797 = 10'h2c3 == r_count_4_io_out ? io_r_707_b : _GEN_3796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3798 = 10'h2c4 == r_count_4_io_out ? io_r_708_b : _GEN_3797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3799 = 10'h2c5 == r_count_4_io_out ? io_r_709_b : _GEN_3798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3800 = 10'h2c6 == r_count_4_io_out ? io_r_710_b : _GEN_3799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3801 = 10'h2c7 == r_count_4_io_out ? io_r_711_b : _GEN_3800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3802 = 10'h2c8 == r_count_4_io_out ? io_r_712_b : _GEN_3801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3803 = 10'h2c9 == r_count_4_io_out ? io_r_713_b : _GEN_3802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3804 = 10'h2ca == r_count_4_io_out ? io_r_714_b : _GEN_3803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3805 = 10'h2cb == r_count_4_io_out ? io_r_715_b : _GEN_3804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3806 = 10'h2cc == r_count_4_io_out ? io_r_716_b : _GEN_3805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3807 = 10'h2cd == r_count_4_io_out ? io_r_717_b : _GEN_3806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3808 = 10'h2ce == r_count_4_io_out ? io_r_718_b : _GEN_3807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3809 = 10'h2cf == r_count_4_io_out ? io_r_719_b : _GEN_3808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3810 = 10'h2d0 == r_count_4_io_out ? io_r_720_b : _GEN_3809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3811 = 10'h2d1 == r_count_4_io_out ? io_r_721_b : _GEN_3810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3812 = 10'h2d2 == r_count_4_io_out ? io_r_722_b : _GEN_3811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3813 = 10'h2d3 == r_count_4_io_out ? io_r_723_b : _GEN_3812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3814 = 10'h2d4 == r_count_4_io_out ? io_r_724_b : _GEN_3813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3815 = 10'h2d5 == r_count_4_io_out ? io_r_725_b : _GEN_3814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3816 = 10'h2d6 == r_count_4_io_out ? io_r_726_b : _GEN_3815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3817 = 10'h2d7 == r_count_4_io_out ? io_r_727_b : _GEN_3816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3818 = 10'h2d8 == r_count_4_io_out ? io_r_728_b : _GEN_3817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3819 = 10'h2d9 == r_count_4_io_out ? io_r_729_b : _GEN_3818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3820 = 10'h2da == r_count_4_io_out ? io_r_730_b : _GEN_3819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3821 = 10'h2db == r_count_4_io_out ? io_r_731_b : _GEN_3820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3822 = 10'h2dc == r_count_4_io_out ? io_r_732_b : _GEN_3821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3823 = 10'h2dd == r_count_4_io_out ? io_r_733_b : _GEN_3822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3824 = 10'h2de == r_count_4_io_out ? io_r_734_b : _GEN_3823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3825 = 10'h2df == r_count_4_io_out ? io_r_735_b : _GEN_3824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3826 = 10'h2e0 == r_count_4_io_out ? io_r_736_b : _GEN_3825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3827 = 10'h2e1 == r_count_4_io_out ? io_r_737_b : _GEN_3826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3828 = 10'h2e2 == r_count_4_io_out ? io_r_738_b : _GEN_3827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3829 = 10'h2e3 == r_count_4_io_out ? io_r_739_b : _GEN_3828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3830 = 10'h2e4 == r_count_4_io_out ? io_r_740_b : _GEN_3829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3831 = 10'h2e5 == r_count_4_io_out ? io_r_741_b : _GEN_3830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3832 = 10'h2e6 == r_count_4_io_out ? io_r_742_b : _GEN_3831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3833 = 10'h2e7 == r_count_4_io_out ? io_r_743_b : _GEN_3832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3834 = 10'h2e8 == r_count_4_io_out ? io_r_744_b : _GEN_3833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3835 = 10'h2e9 == r_count_4_io_out ? io_r_745_b : _GEN_3834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3836 = 10'h2ea == r_count_4_io_out ? io_r_746_b : _GEN_3835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3837 = 10'h2eb == r_count_4_io_out ? io_r_747_b : _GEN_3836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3838 = 10'h2ec == r_count_4_io_out ? io_r_748_b : _GEN_3837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3841 = 10'h1 == r_count_5_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3842 = 10'h2 == r_count_5_io_out ? io_r_2_b : _GEN_3841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3843 = 10'h3 == r_count_5_io_out ? io_r_3_b : _GEN_3842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3844 = 10'h4 == r_count_5_io_out ? io_r_4_b : _GEN_3843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3845 = 10'h5 == r_count_5_io_out ? io_r_5_b : _GEN_3844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3846 = 10'h6 == r_count_5_io_out ? io_r_6_b : _GEN_3845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3847 = 10'h7 == r_count_5_io_out ? io_r_7_b : _GEN_3846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3848 = 10'h8 == r_count_5_io_out ? io_r_8_b : _GEN_3847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3849 = 10'h9 == r_count_5_io_out ? io_r_9_b : _GEN_3848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3850 = 10'ha == r_count_5_io_out ? io_r_10_b : _GEN_3849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3851 = 10'hb == r_count_5_io_out ? io_r_11_b : _GEN_3850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3852 = 10'hc == r_count_5_io_out ? io_r_12_b : _GEN_3851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3853 = 10'hd == r_count_5_io_out ? io_r_13_b : _GEN_3852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3854 = 10'he == r_count_5_io_out ? io_r_14_b : _GEN_3853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3855 = 10'hf == r_count_5_io_out ? io_r_15_b : _GEN_3854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3856 = 10'h10 == r_count_5_io_out ? io_r_16_b : _GEN_3855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3857 = 10'h11 == r_count_5_io_out ? io_r_17_b : _GEN_3856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3858 = 10'h12 == r_count_5_io_out ? io_r_18_b : _GEN_3857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3859 = 10'h13 == r_count_5_io_out ? io_r_19_b : _GEN_3858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3860 = 10'h14 == r_count_5_io_out ? io_r_20_b : _GEN_3859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3861 = 10'h15 == r_count_5_io_out ? io_r_21_b : _GEN_3860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3862 = 10'h16 == r_count_5_io_out ? io_r_22_b : _GEN_3861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3863 = 10'h17 == r_count_5_io_out ? io_r_23_b : _GEN_3862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3864 = 10'h18 == r_count_5_io_out ? io_r_24_b : _GEN_3863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3865 = 10'h19 == r_count_5_io_out ? io_r_25_b : _GEN_3864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3866 = 10'h1a == r_count_5_io_out ? io_r_26_b : _GEN_3865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3867 = 10'h1b == r_count_5_io_out ? io_r_27_b : _GEN_3866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3868 = 10'h1c == r_count_5_io_out ? io_r_28_b : _GEN_3867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3869 = 10'h1d == r_count_5_io_out ? io_r_29_b : _GEN_3868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3870 = 10'h1e == r_count_5_io_out ? io_r_30_b : _GEN_3869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3871 = 10'h1f == r_count_5_io_out ? io_r_31_b : _GEN_3870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3872 = 10'h20 == r_count_5_io_out ? io_r_32_b : _GEN_3871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3873 = 10'h21 == r_count_5_io_out ? io_r_33_b : _GEN_3872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3874 = 10'h22 == r_count_5_io_out ? io_r_34_b : _GEN_3873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3875 = 10'h23 == r_count_5_io_out ? io_r_35_b : _GEN_3874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3876 = 10'h24 == r_count_5_io_out ? io_r_36_b : _GEN_3875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3877 = 10'h25 == r_count_5_io_out ? io_r_37_b : _GEN_3876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3878 = 10'h26 == r_count_5_io_out ? io_r_38_b : _GEN_3877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3879 = 10'h27 == r_count_5_io_out ? io_r_39_b : _GEN_3878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3880 = 10'h28 == r_count_5_io_out ? io_r_40_b : _GEN_3879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3881 = 10'h29 == r_count_5_io_out ? io_r_41_b : _GEN_3880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3882 = 10'h2a == r_count_5_io_out ? io_r_42_b : _GEN_3881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3883 = 10'h2b == r_count_5_io_out ? io_r_43_b : _GEN_3882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3884 = 10'h2c == r_count_5_io_out ? io_r_44_b : _GEN_3883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3885 = 10'h2d == r_count_5_io_out ? io_r_45_b : _GEN_3884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3886 = 10'h2e == r_count_5_io_out ? io_r_46_b : _GEN_3885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3887 = 10'h2f == r_count_5_io_out ? io_r_47_b : _GEN_3886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3888 = 10'h30 == r_count_5_io_out ? io_r_48_b : _GEN_3887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3889 = 10'h31 == r_count_5_io_out ? io_r_49_b : _GEN_3888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3890 = 10'h32 == r_count_5_io_out ? io_r_50_b : _GEN_3889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3891 = 10'h33 == r_count_5_io_out ? io_r_51_b : _GEN_3890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3892 = 10'h34 == r_count_5_io_out ? io_r_52_b : _GEN_3891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3893 = 10'h35 == r_count_5_io_out ? io_r_53_b : _GEN_3892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3894 = 10'h36 == r_count_5_io_out ? io_r_54_b : _GEN_3893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3895 = 10'h37 == r_count_5_io_out ? io_r_55_b : _GEN_3894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3896 = 10'h38 == r_count_5_io_out ? io_r_56_b : _GEN_3895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3897 = 10'h39 == r_count_5_io_out ? io_r_57_b : _GEN_3896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3898 = 10'h3a == r_count_5_io_out ? io_r_58_b : _GEN_3897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3899 = 10'h3b == r_count_5_io_out ? io_r_59_b : _GEN_3898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3900 = 10'h3c == r_count_5_io_out ? io_r_60_b : _GEN_3899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3901 = 10'h3d == r_count_5_io_out ? io_r_61_b : _GEN_3900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3902 = 10'h3e == r_count_5_io_out ? io_r_62_b : _GEN_3901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3903 = 10'h3f == r_count_5_io_out ? io_r_63_b : _GEN_3902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3904 = 10'h40 == r_count_5_io_out ? io_r_64_b : _GEN_3903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3905 = 10'h41 == r_count_5_io_out ? io_r_65_b : _GEN_3904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3906 = 10'h42 == r_count_5_io_out ? io_r_66_b : _GEN_3905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3907 = 10'h43 == r_count_5_io_out ? io_r_67_b : _GEN_3906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3908 = 10'h44 == r_count_5_io_out ? io_r_68_b : _GEN_3907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3909 = 10'h45 == r_count_5_io_out ? io_r_69_b : _GEN_3908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3910 = 10'h46 == r_count_5_io_out ? io_r_70_b : _GEN_3909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3911 = 10'h47 == r_count_5_io_out ? io_r_71_b : _GEN_3910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3912 = 10'h48 == r_count_5_io_out ? io_r_72_b : _GEN_3911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3913 = 10'h49 == r_count_5_io_out ? io_r_73_b : _GEN_3912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3914 = 10'h4a == r_count_5_io_out ? io_r_74_b : _GEN_3913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3915 = 10'h4b == r_count_5_io_out ? io_r_75_b : _GEN_3914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3916 = 10'h4c == r_count_5_io_out ? io_r_76_b : _GEN_3915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3917 = 10'h4d == r_count_5_io_out ? io_r_77_b : _GEN_3916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3918 = 10'h4e == r_count_5_io_out ? io_r_78_b : _GEN_3917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3919 = 10'h4f == r_count_5_io_out ? io_r_79_b : _GEN_3918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3920 = 10'h50 == r_count_5_io_out ? io_r_80_b : _GEN_3919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3921 = 10'h51 == r_count_5_io_out ? io_r_81_b : _GEN_3920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3922 = 10'h52 == r_count_5_io_out ? io_r_82_b : _GEN_3921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3923 = 10'h53 == r_count_5_io_out ? io_r_83_b : _GEN_3922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3924 = 10'h54 == r_count_5_io_out ? io_r_84_b : _GEN_3923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3925 = 10'h55 == r_count_5_io_out ? io_r_85_b : _GEN_3924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3926 = 10'h56 == r_count_5_io_out ? io_r_86_b : _GEN_3925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3927 = 10'h57 == r_count_5_io_out ? io_r_87_b : _GEN_3926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3928 = 10'h58 == r_count_5_io_out ? io_r_88_b : _GEN_3927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3929 = 10'h59 == r_count_5_io_out ? io_r_89_b : _GEN_3928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3930 = 10'h5a == r_count_5_io_out ? io_r_90_b : _GEN_3929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3931 = 10'h5b == r_count_5_io_out ? io_r_91_b : _GEN_3930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3932 = 10'h5c == r_count_5_io_out ? io_r_92_b : _GEN_3931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3933 = 10'h5d == r_count_5_io_out ? io_r_93_b : _GEN_3932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3934 = 10'h5e == r_count_5_io_out ? io_r_94_b : _GEN_3933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3935 = 10'h5f == r_count_5_io_out ? io_r_95_b : _GEN_3934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3936 = 10'h60 == r_count_5_io_out ? io_r_96_b : _GEN_3935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3937 = 10'h61 == r_count_5_io_out ? io_r_97_b : _GEN_3936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3938 = 10'h62 == r_count_5_io_out ? io_r_98_b : _GEN_3937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3939 = 10'h63 == r_count_5_io_out ? io_r_99_b : _GEN_3938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3940 = 10'h64 == r_count_5_io_out ? io_r_100_b : _GEN_3939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3941 = 10'h65 == r_count_5_io_out ? io_r_101_b : _GEN_3940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3942 = 10'h66 == r_count_5_io_out ? io_r_102_b : _GEN_3941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3943 = 10'h67 == r_count_5_io_out ? io_r_103_b : _GEN_3942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3944 = 10'h68 == r_count_5_io_out ? io_r_104_b : _GEN_3943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3945 = 10'h69 == r_count_5_io_out ? io_r_105_b : _GEN_3944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3946 = 10'h6a == r_count_5_io_out ? io_r_106_b : _GEN_3945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3947 = 10'h6b == r_count_5_io_out ? io_r_107_b : _GEN_3946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3948 = 10'h6c == r_count_5_io_out ? io_r_108_b : _GEN_3947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3949 = 10'h6d == r_count_5_io_out ? io_r_109_b : _GEN_3948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3950 = 10'h6e == r_count_5_io_out ? io_r_110_b : _GEN_3949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3951 = 10'h6f == r_count_5_io_out ? io_r_111_b : _GEN_3950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3952 = 10'h70 == r_count_5_io_out ? io_r_112_b : _GEN_3951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3953 = 10'h71 == r_count_5_io_out ? io_r_113_b : _GEN_3952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3954 = 10'h72 == r_count_5_io_out ? io_r_114_b : _GEN_3953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3955 = 10'h73 == r_count_5_io_out ? io_r_115_b : _GEN_3954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3956 = 10'h74 == r_count_5_io_out ? io_r_116_b : _GEN_3955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3957 = 10'h75 == r_count_5_io_out ? io_r_117_b : _GEN_3956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3958 = 10'h76 == r_count_5_io_out ? io_r_118_b : _GEN_3957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3959 = 10'h77 == r_count_5_io_out ? io_r_119_b : _GEN_3958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3960 = 10'h78 == r_count_5_io_out ? io_r_120_b : _GEN_3959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3961 = 10'h79 == r_count_5_io_out ? io_r_121_b : _GEN_3960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3962 = 10'h7a == r_count_5_io_out ? io_r_122_b : _GEN_3961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3963 = 10'h7b == r_count_5_io_out ? io_r_123_b : _GEN_3962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3964 = 10'h7c == r_count_5_io_out ? io_r_124_b : _GEN_3963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3965 = 10'h7d == r_count_5_io_out ? io_r_125_b : _GEN_3964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3966 = 10'h7e == r_count_5_io_out ? io_r_126_b : _GEN_3965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3967 = 10'h7f == r_count_5_io_out ? io_r_127_b : _GEN_3966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3968 = 10'h80 == r_count_5_io_out ? io_r_128_b : _GEN_3967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3969 = 10'h81 == r_count_5_io_out ? io_r_129_b : _GEN_3968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3970 = 10'h82 == r_count_5_io_out ? io_r_130_b : _GEN_3969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3971 = 10'h83 == r_count_5_io_out ? io_r_131_b : _GEN_3970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3972 = 10'h84 == r_count_5_io_out ? io_r_132_b : _GEN_3971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3973 = 10'h85 == r_count_5_io_out ? io_r_133_b : _GEN_3972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3974 = 10'h86 == r_count_5_io_out ? io_r_134_b : _GEN_3973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3975 = 10'h87 == r_count_5_io_out ? io_r_135_b : _GEN_3974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3976 = 10'h88 == r_count_5_io_out ? io_r_136_b : _GEN_3975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3977 = 10'h89 == r_count_5_io_out ? io_r_137_b : _GEN_3976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3978 = 10'h8a == r_count_5_io_out ? io_r_138_b : _GEN_3977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3979 = 10'h8b == r_count_5_io_out ? io_r_139_b : _GEN_3978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3980 = 10'h8c == r_count_5_io_out ? io_r_140_b : _GEN_3979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3981 = 10'h8d == r_count_5_io_out ? io_r_141_b : _GEN_3980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3982 = 10'h8e == r_count_5_io_out ? io_r_142_b : _GEN_3981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3983 = 10'h8f == r_count_5_io_out ? io_r_143_b : _GEN_3982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3984 = 10'h90 == r_count_5_io_out ? io_r_144_b : _GEN_3983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3985 = 10'h91 == r_count_5_io_out ? io_r_145_b : _GEN_3984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3986 = 10'h92 == r_count_5_io_out ? io_r_146_b : _GEN_3985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3987 = 10'h93 == r_count_5_io_out ? io_r_147_b : _GEN_3986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3988 = 10'h94 == r_count_5_io_out ? io_r_148_b : _GEN_3987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3989 = 10'h95 == r_count_5_io_out ? io_r_149_b : _GEN_3988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3990 = 10'h96 == r_count_5_io_out ? io_r_150_b : _GEN_3989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3991 = 10'h97 == r_count_5_io_out ? io_r_151_b : _GEN_3990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3992 = 10'h98 == r_count_5_io_out ? io_r_152_b : _GEN_3991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3993 = 10'h99 == r_count_5_io_out ? io_r_153_b : _GEN_3992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3994 = 10'h9a == r_count_5_io_out ? io_r_154_b : _GEN_3993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3995 = 10'h9b == r_count_5_io_out ? io_r_155_b : _GEN_3994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3996 = 10'h9c == r_count_5_io_out ? io_r_156_b : _GEN_3995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3997 = 10'h9d == r_count_5_io_out ? io_r_157_b : _GEN_3996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3998 = 10'h9e == r_count_5_io_out ? io_r_158_b : _GEN_3997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3999 = 10'h9f == r_count_5_io_out ? io_r_159_b : _GEN_3998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4000 = 10'ha0 == r_count_5_io_out ? io_r_160_b : _GEN_3999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4001 = 10'ha1 == r_count_5_io_out ? io_r_161_b : _GEN_4000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4002 = 10'ha2 == r_count_5_io_out ? io_r_162_b : _GEN_4001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4003 = 10'ha3 == r_count_5_io_out ? io_r_163_b : _GEN_4002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4004 = 10'ha4 == r_count_5_io_out ? io_r_164_b : _GEN_4003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4005 = 10'ha5 == r_count_5_io_out ? io_r_165_b : _GEN_4004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4006 = 10'ha6 == r_count_5_io_out ? io_r_166_b : _GEN_4005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4007 = 10'ha7 == r_count_5_io_out ? io_r_167_b : _GEN_4006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4008 = 10'ha8 == r_count_5_io_out ? io_r_168_b : _GEN_4007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4009 = 10'ha9 == r_count_5_io_out ? io_r_169_b : _GEN_4008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4010 = 10'haa == r_count_5_io_out ? io_r_170_b : _GEN_4009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4011 = 10'hab == r_count_5_io_out ? io_r_171_b : _GEN_4010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4012 = 10'hac == r_count_5_io_out ? io_r_172_b : _GEN_4011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4013 = 10'had == r_count_5_io_out ? io_r_173_b : _GEN_4012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4014 = 10'hae == r_count_5_io_out ? io_r_174_b : _GEN_4013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4015 = 10'haf == r_count_5_io_out ? io_r_175_b : _GEN_4014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4016 = 10'hb0 == r_count_5_io_out ? io_r_176_b : _GEN_4015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4017 = 10'hb1 == r_count_5_io_out ? io_r_177_b : _GEN_4016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4018 = 10'hb2 == r_count_5_io_out ? io_r_178_b : _GEN_4017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4019 = 10'hb3 == r_count_5_io_out ? io_r_179_b : _GEN_4018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4020 = 10'hb4 == r_count_5_io_out ? io_r_180_b : _GEN_4019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4021 = 10'hb5 == r_count_5_io_out ? io_r_181_b : _GEN_4020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4022 = 10'hb6 == r_count_5_io_out ? io_r_182_b : _GEN_4021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4023 = 10'hb7 == r_count_5_io_out ? io_r_183_b : _GEN_4022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4024 = 10'hb8 == r_count_5_io_out ? io_r_184_b : _GEN_4023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4025 = 10'hb9 == r_count_5_io_out ? io_r_185_b : _GEN_4024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4026 = 10'hba == r_count_5_io_out ? io_r_186_b : _GEN_4025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4027 = 10'hbb == r_count_5_io_out ? io_r_187_b : _GEN_4026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4028 = 10'hbc == r_count_5_io_out ? io_r_188_b : _GEN_4027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4029 = 10'hbd == r_count_5_io_out ? io_r_189_b : _GEN_4028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4030 = 10'hbe == r_count_5_io_out ? io_r_190_b : _GEN_4029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4031 = 10'hbf == r_count_5_io_out ? io_r_191_b : _GEN_4030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4032 = 10'hc0 == r_count_5_io_out ? io_r_192_b : _GEN_4031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4033 = 10'hc1 == r_count_5_io_out ? io_r_193_b : _GEN_4032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4034 = 10'hc2 == r_count_5_io_out ? io_r_194_b : _GEN_4033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4035 = 10'hc3 == r_count_5_io_out ? io_r_195_b : _GEN_4034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4036 = 10'hc4 == r_count_5_io_out ? io_r_196_b : _GEN_4035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4037 = 10'hc5 == r_count_5_io_out ? io_r_197_b : _GEN_4036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4038 = 10'hc6 == r_count_5_io_out ? io_r_198_b : _GEN_4037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4039 = 10'hc7 == r_count_5_io_out ? io_r_199_b : _GEN_4038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4040 = 10'hc8 == r_count_5_io_out ? io_r_200_b : _GEN_4039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4041 = 10'hc9 == r_count_5_io_out ? io_r_201_b : _GEN_4040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4042 = 10'hca == r_count_5_io_out ? io_r_202_b : _GEN_4041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4043 = 10'hcb == r_count_5_io_out ? io_r_203_b : _GEN_4042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4044 = 10'hcc == r_count_5_io_out ? io_r_204_b : _GEN_4043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4045 = 10'hcd == r_count_5_io_out ? io_r_205_b : _GEN_4044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4046 = 10'hce == r_count_5_io_out ? io_r_206_b : _GEN_4045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4047 = 10'hcf == r_count_5_io_out ? io_r_207_b : _GEN_4046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4048 = 10'hd0 == r_count_5_io_out ? io_r_208_b : _GEN_4047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4049 = 10'hd1 == r_count_5_io_out ? io_r_209_b : _GEN_4048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4050 = 10'hd2 == r_count_5_io_out ? io_r_210_b : _GEN_4049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4051 = 10'hd3 == r_count_5_io_out ? io_r_211_b : _GEN_4050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4052 = 10'hd4 == r_count_5_io_out ? io_r_212_b : _GEN_4051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4053 = 10'hd5 == r_count_5_io_out ? io_r_213_b : _GEN_4052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4054 = 10'hd6 == r_count_5_io_out ? io_r_214_b : _GEN_4053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4055 = 10'hd7 == r_count_5_io_out ? io_r_215_b : _GEN_4054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4056 = 10'hd8 == r_count_5_io_out ? io_r_216_b : _GEN_4055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4057 = 10'hd9 == r_count_5_io_out ? io_r_217_b : _GEN_4056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4058 = 10'hda == r_count_5_io_out ? io_r_218_b : _GEN_4057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4059 = 10'hdb == r_count_5_io_out ? io_r_219_b : _GEN_4058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4060 = 10'hdc == r_count_5_io_out ? io_r_220_b : _GEN_4059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4061 = 10'hdd == r_count_5_io_out ? io_r_221_b : _GEN_4060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4062 = 10'hde == r_count_5_io_out ? io_r_222_b : _GEN_4061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4063 = 10'hdf == r_count_5_io_out ? io_r_223_b : _GEN_4062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4064 = 10'he0 == r_count_5_io_out ? io_r_224_b : _GEN_4063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4065 = 10'he1 == r_count_5_io_out ? io_r_225_b : _GEN_4064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4066 = 10'he2 == r_count_5_io_out ? io_r_226_b : _GEN_4065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4067 = 10'he3 == r_count_5_io_out ? io_r_227_b : _GEN_4066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4068 = 10'he4 == r_count_5_io_out ? io_r_228_b : _GEN_4067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4069 = 10'he5 == r_count_5_io_out ? io_r_229_b : _GEN_4068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4070 = 10'he6 == r_count_5_io_out ? io_r_230_b : _GEN_4069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4071 = 10'he7 == r_count_5_io_out ? io_r_231_b : _GEN_4070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4072 = 10'he8 == r_count_5_io_out ? io_r_232_b : _GEN_4071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4073 = 10'he9 == r_count_5_io_out ? io_r_233_b : _GEN_4072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4074 = 10'hea == r_count_5_io_out ? io_r_234_b : _GEN_4073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4075 = 10'heb == r_count_5_io_out ? io_r_235_b : _GEN_4074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4076 = 10'hec == r_count_5_io_out ? io_r_236_b : _GEN_4075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4077 = 10'hed == r_count_5_io_out ? io_r_237_b : _GEN_4076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4078 = 10'hee == r_count_5_io_out ? io_r_238_b : _GEN_4077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4079 = 10'hef == r_count_5_io_out ? io_r_239_b : _GEN_4078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4080 = 10'hf0 == r_count_5_io_out ? io_r_240_b : _GEN_4079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4081 = 10'hf1 == r_count_5_io_out ? io_r_241_b : _GEN_4080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4082 = 10'hf2 == r_count_5_io_out ? io_r_242_b : _GEN_4081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4083 = 10'hf3 == r_count_5_io_out ? io_r_243_b : _GEN_4082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4084 = 10'hf4 == r_count_5_io_out ? io_r_244_b : _GEN_4083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4085 = 10'hf5 == r_count_5_io_out ? io_r_245_b : _GEN_4084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4086 = 10'hf6 == r_count_5_io_out ? io_r_246_b : _GEN_4085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4087 = 10'hf7 == r_count_5_io_out ? io_r_247_b : _GEN_4086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4088 = 10'hf8 == r_count_5_io_out ? io_r_248_b : _GEN_4087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4089 = 10'hf9 == r_count_5_io_out ? io_r_249_b : _GEN_4088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4090 = 10'hfa == r_count_5_io_out ? io_r_250_b : _GEN_4089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4091 = 10'hfb == r_count_5_io_out ? io_r_251_b : _GEN_4090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4092 = 10'hfc == r_count_5_io_out ? io_r_252_b : _GEN_4091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4093 = 10'hfd == r_count_5_io_out ? io_r_253_b : _GEN_4092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4094 = 10'hfe == r_count_5_io_out ? io_r_254_b : _GEN_4093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4095 = 10'hff == r_count_5_io_out ? io_r_255_b : _GEN_4094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4096 = 10'h100 == r_count_5_io_out ? io_r_256_b : _GEN_4095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4097 = 10'h101 == r_count_5_io_out ? io_r_257_b : _GEN_4096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4098 = 10'h102 == r_count_5_io_out ? io_r_258_b : _GEN_4097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4099 = 10'h103 == r_count_5_io_out ? io_r_259_b : _GEN_4098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4100 = 10'h104 == r_count_5_io_out ? io_r_260_b : _GEN_4099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4101 = 10'h105 == r_count_5_io_out ? io_r_261_b : _GEN_4100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4102 = 10'h106 == r_count_5_io_out ? io_r_262_b : _GEN_4101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4103 = 10'h107 == r_count_5_io_out ? io_r_263_b : _GEN_4102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4104 = 10'h108 == r_count_5_io_out ? io_r_264_b : _GEN_4103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4105 = 10'h109 == r_count_5_io_out ? io_r_265_b : _GEN_4104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4106 = 10'h10a == r_count_5_io_out ? io_r_266_b : _GEN_4105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4107 = 10'h10b == r_count_5_io_out ? io_r_267_b : _GEN_4106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4108 = 10'h10c == r_count_5_io_out ? io_r_268_b : _GEN_4107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4109 = 10'h10d == r_count_5_io_out ? io_r_269_b : _GEN_4108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4110 = 10'h10e == r_count_5_io_out ? io_r_270_b : _GEN_4109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4111 = 10'h10f == r_count_5_io_out ? io_r_271_b : _GEN_4110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4112 = 10'h110 == r_count_5_io_out ? io_r_272_b : _GEN_4111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4113 = 10'h111 == r_count_5_io_out ? io_r_273_b : _GEN_4112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4114 = 10'h112 == r_count_5_io_out ? io_r_274_b : _GEN_4113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4115 = 10'h113 == r_count_5_io_out ? io_r_275_b : _GEN_4114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4116 = 10'h114 == r_count_5_io_out ? io_r_276_b : _GEN_4115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4117 = 10'h115 == r_count_5_io_out ? io_r_277_b : _GEN_4116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4118 = 10'h116 == r_count_5_io_out ? io_r_278_b : _GEN_4117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4119 = 10'h117 == r_count_5_io_out ? io_r_279_b : _GEN_4118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4120 = 10'h118 == r_count_5_io_out ? io_r_280_b : _GEN_4119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4121 = 10'h119 == r_count_5_io_out ? io_r_281_b : _GEN_4120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4122 = 10'h11a == r_count_5_io_out ? io_r_282_b : _GEN_4121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4123 = 10'h11b == r_count_5_io_out ? io_r_283_b : _GEN_4122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4124 = 10'h11c == r_count_5_io_out ? io_r_284_b : _GEN_4123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4125 = 10'h11d == r_count_5_io_out ? io_r_285_b : _GEN_4124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4126 = 10'h11e == r_count_5_io_out ? io_r_286_b : _GEN_4125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4127 = 10'h11f == r_count_5_io_out ? io_r_287_b : _GEN_4126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4128 = 10'h120 == r_count_5_io_out ? io_r_288_b : _GEN_4127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4129 = 10'h121 == r_count_5_io_out ? io_r_289_b : _GEN_4128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4130 = 10'h122 == r_count_5_io_out ? io_r_290_b : _GEN_4129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4131 = 10'h123 == r_count_5_io_out ? io_r_291_b : _GEN_4130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4132 = 10'h124 == r_count_5_io_out ? io_r_292_b : _GEN_4131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4133 = 10'h125 == r_count_5_io_out ? io_r_293_b : _GEN_4132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4134 = 10'h126 == r_count_5_io_out ? io_r_294_b : _GEN_4133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4135 = 10'h127 == r_count_5_io_out ? io_r_295_b : _GEN_4134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4136 = 10'h128 == r_count_5_io_out ? io_r_296_b : _GEN_4135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4137 = 10'h129 == r_count_5_io_out ? io_r_297_b : _GEN_4136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4138 = 10'h12a == r_count_5_io_out ? io_r_298_b : _GEN_4137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4139 = 10'h12b == r_count_5_io_out ? io_r_299_b : _GEN_4138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4140 = 10'h12c == r_count_5_io_out ? io_r_300_b : _GEN_4139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4141 = 10'h12d == r_count_5_io_out ? io_r_301_b : _GEN_4140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4142 = 10'h12e == r_count_5_io_out ? io_r_302_b : _GEN_4141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4143 = 10'h12f == r_count_5_io_out ? io_r_303_b : _GEN_4142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4144 = 10'h130 == r_count_5_io_out ? io_r_304_b : _GEN_4143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4145 = 10'h131 == r_count_5_io_out ? io_r_305_b : _GEN_4144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4146 = 10'h132 == r_count_5_io_out ? io_r_306_b : _GEN_4145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4147 = 10'h133 == r_count_5_io_out ? io_r_307_b : _GEN_4146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4148 = 10'h134 == r_count_5_io_out ? io_r_308_b : _GEN_4147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4149 = 10'h135 == r_count_5_io_out ? io_r_309_b : _GEN_4148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4150 = 10'h136 == r_count_5_io_out ? io_r_310_b : _GEN_4149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4151 = 10'h137 == r_count_5_io_out ? io_r_311_b : _GEN_4150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4152 = 10'h138 == r_count_5_io_out ? io_r_312_b : _GEN_4151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4153 = 10'h139 == r_count_5_io_out ? io_r_313_b : _GEN_4152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4154 = 10'h13a == r_count_5_io_out ? io_r_314_b : _GEN_4153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4155 = 10'h13b == r_count_5_io_out ? io_r_315_b : _GEN_4154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4156 = 10'h13c == r_count_5_io_out ? io_r_316_b : _GEN_4155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4157 = 10'h13d == r_count_5_io_out ? io_r_317_b : _GEN_4156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4158 = 10'h13e == r_count_5_io_out ? io_r_318_b : _GEN_4157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4159 = 10'h13f == r_count_5_io_out ? io_r_319_b : _GEN_4158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4160 = 10'h140 == r_count_5_io_out ? io_r_320_b : _GEN_4159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4161 = 10'h141 == r_count_5_io_out ? io_r_321_b : _GEN_4160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4162 = 10'h142 == r_count_5_io_out ? io_r_322_b : _GEN_4161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4163 = 10'h143 == r_count_5_io_out ? io_r_323_b : _GEN_4162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4164 = 10'h144 == r_count_5_io_out ? io_r_324_b : _GEN_4163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4165 = 10'h145 == r_count_5_io_out ? io_r_325_b : _GEN_4164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4166 = 10'h146 == r_count_5_io_out ? io_r_326_b : _GEN_4165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4167 = 10'h147 == r_count_5_io_out ? io_r_327_b : _GEN_4166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4168 = 10'h148 == r_count_5_io_out ? io_r_328_b : _GEN_4167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4169 = 10'h149 == r_count_5_io_out ? io_r_329_b : _GEN_4168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4170 = 10'h14a == r_count_5_io_out ? io_r_330_b : _GEN_4169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4171 = 10'h14b == r_count_5_io_out ? io_r_331_b : _GEN_4170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4172 = 10'h14c == r_count_5_io_out ? io_r_332_b : _GEN_4171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4173 = 10'h14d == r_count_5_io_out ? io_r_333_b : _GEN_4172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4174 = 10'h14e == r_count_5_io_out ? io_r_334_b : _GEN_4173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4175 = 10'h14f == r_count_5_io_out ? io_r_335_b : _GEN_4174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4176 = 10'h150 == r_count_5_io_out ? io_r_336_b : _GEN_4175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4177 = 10'h151 == r_count_5_io_out ? io_r_337_b : _GEN_4176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4178 = 10'h152 == r_count_5_io_out ? io_r_338_b : _GEN_4177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4179 = 10'h153 == r_count_5_io_out ? io_r_339_b : _GEN_4178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4180 = 10'h154 == r_count_5_io_out ? io_r_340_b : _GEN_4179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4181 = 10'h155 == r_count_5_io_out ? io_r_341_b : _GEN_4180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4182 = 10'h156 == r_count_5_io_out ? io_r_342_b : _GEN_4181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4183 = 10'h157 == r_count_5_io_out ? io_r_343_b : _GEN_4182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4184 = 10'h158 == r_count_5_io_out ? io_r_344_b : _GEN_4183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4185 = 10'h159 == r_count_5_io_out ? io_r_345_b : _GEN_4184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4186 = 10'h15a == r_count_5_io_out ? io_r_346_b : _GEN_4185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4187 = 10'h15b == r_count_5_io_out ? io_r_347_b : _GEN_4186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4188 = 10'h15c == r_count_5_io_out ? io_r_348_b : _GEN_4187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4189 = 10'h15d == r_count_5_io_out ? io_r_349_b : _GEN_4188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4190 = 10'h15e == r_count_5_io_out ? io_r_350_b : _GEN_4189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4191 = 10'h15f == r_count_5_io_out ? io_r_351_b : _GEN_4190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4192 = 10'h160 == r_count_5_io_out ? io_r_352_b : _GEN_4191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4193 = 10'h161 == r_count_5_io_out ? io_r_353_b : _GEN_4192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4194 = 10'h162 == r_count_5_io_out ? io_r_354_b : _GEN_4193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4195 = 10'h163 == r_count_5_io_out ? io_r_355_b : _GEN_4194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4196 = 10'h164 == r_count_5_io_out ? io_r_356_b : _GEN_4195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4197 = 10'h165 == r_count_5_io_out ? io_r_357_b : _GEN_4196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4198 = 10'h166 == r_count_5_io_out ? io_r_358_b : _GEN_4197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4199 = 10'h167 == r_count_5_io_out ? io_r_359_b : _GEN_4198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4200 = 10'h168 == r_count_5_io_out ? io_r_360_b : _GEN_4199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4201 = 10'h169 == r_count_5_io_out ? io_r_361_b : _GEN_4200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4202 = 10'h16a == r_count_5_io_out ? io_r_362_b : _GEN_4201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4203 = 10'h16b == r_count_5_io_out ? io_r_363_b : _GEN_4202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4204 = 10'h16c == r_count_5_io_out ? io_r_364_b : _GEN_4203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4205 = 10'h16d == r_count_5_io_out ? io_r_365_b : _GEN_4204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4206 = 10'h16e == r_count_5_io_out ? io_r_366_b : _GEN_4205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4207 = 10'h16f == r_count_5_io_out ? io_r_367_b : _GEN_4206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4208 = 10'h170 == r_count_5_io_out ? io_r_368_b : _GEN_4207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4209 = 10'h171 == r_count_5_io_out ? io_r_369_b : _GEN_4208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4210 = 10'h172 == r_count_5_io_out ? io_r_370_b : _GEN_4209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4211 = 10'h173 == r_count_5_io_out ? io_r_371_b : _GEN_4210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4212 = 10'h174 == r_count_5_io_out ? io_r_372_b : _GEN_4211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4213 = 10'h175 == r_count_5_io_out ? io_r_373_b : _GEN_4212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4214 = 10'h176 == r_count_5_io_out ? io_r_374_b : _GEN_4213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4215 = 10'h177 == r_count_5_io_out ? io_r_375_b : _GEN_4214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4216 = 10'h178 == r_count_5_io_out ? io_r_376_b : _GEN_4215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4217 = 10'h179 == r_count_5_io_out ? io_r_377_b : _GEN_4216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4218 = 10'h17a == r_count_5_io_out ? io_r_378_b : _GEN_4217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4219 = 10'h17b == r_count_5_io_out ? io_r_379_b : _GEN_4218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4220 = 10'h17c == r_count_5_io_out ? io_r_380_b : _GEN_4219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4221 = 10'h17d == r_count_5_io_out ? io_r_381_b : _GEN_4220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4222 = 10'h17e == r_count_5_io_out ? io_r_382_b : _GEN_4221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4223 = 10'h17f == r_count_5_io_out ? io_r_383_b : _GEN_4222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4224 = 10'h180 == r_count_5_io_out ? io_r_384_b : _GEN_4223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4225 = 10'h181 == r_count_5_io_out ? io_r_385_b : _GEN_4224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4226 = 10'h182 == r_count_5_io_out ? io_r_386_b : _GEN_4225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4227 = 10'h183 == r_count_5_io_out ? io_r_387_b : _GEN_4226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4228 = 10'h184 == r_count_5_io_out ? io_r_388_b : _GEN_4227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4229 = 10'h185 == r_count_5_io_out ? io_r_389_b : _GEN_4228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4230 = 10'h186 == r_count_5_io_out ? io_r_390_b : _GEN_4229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4231 = 10'h187 == r_count_5_io_out ? io_r_391_b : _GEN_4230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4232 = 10'h188 == r_count_5_io_out ? io_r_392_b : _GEN_4231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4233 = 10'h189 == r_count_5_io_out ? io_r_393_b : _GEN_4232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4234 = 10'h18a == r_count_5_io_out ? io_r_394_b : _GEN_4233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4235 = 10'h18b == r_count_5_io_out ? io_r_395_b : _GEN_4234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4236 = 10'h18c == r_count_5_io_out ? io_r_396_b : _GEN_4235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4237 = 10'h18d == r_count_5_io_out ? io_r_397_b : _GEN_4236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4238 = 10'h18e == r_count_5_io_out ? io_r_398_b : _GEN_4237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4239 = 10'h18f == r_count_5_io_out ? io_r_399_b : _GEN_4238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4240 = 10'h190 == r_count_5_io_out ? io_r_400_b : _GEN_4239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4241 = 10'h191 == r_count_5_io_out ? io_r_401_b : _GEN_4240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4242 = 10'h192 == r_count_5_io_out ? io_r_402_b : _GEN_4241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4243 = 10'h193 == r_count_5_io_out ? io_r_403_b : _GEN_4242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4244 = 10'h194 == r_count_5_io_out ? io_r_404_b : _GEN_4243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4245 = 10'h195 == r_count_5_io_out ? io_r_405_b : _GEN_4244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4246 = 10'h196 == r_count_5_io_out ? io_r_406_b : _GEN_4245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4247 = 10'h197 == r_count_5_io_out ? io_r_407_b : _GEN_4246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4248 = 10'h198 == r_count_5_io_out ? io_r_408_b : _GEN_4247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4249 = 10'h199 == r_count_5_io_out ? io_r_409_b : _GEN_4248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4250 = 10'h19a == r_count_5_io_out ? io_r_410_b : _GEN_4249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4251 = 10'h19b == r_count_5_io_out ? io_r_411_b : _GEN_4250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4252 = 10'h19c == r_count_5_io_out ? io_r_412_b : _GEN_4251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4253 = 10'h19d == r_count_5_io_out ? io_r_413_b : _GEN_4252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4254 = 10'h19e == r_count_5_io_out ? io_r_414_b : _GEN_4253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4255 = 10'h19f == r_count_5_io_out ? io_r_415_b : _GEN_4254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4256 = 10'h1a0 == r_count_5_io_out ? io_r_416_b : _GEN_4255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4257 = 10'h1a1 == r_count_5_io_out ? io_r_417_b : _GEN_4256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4258 = 10'h1a2 == r_count_5_io_out ? io_r_418_b : _GEN_4257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4259 = 10'h1a3 == r_count_5_io_out ? io_r_419_b : _GEN_4258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4260 = 10'h1a4 == r_count_5_io_out ? io_r_420_b : _GEN_4259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4261 = 10'h1a5 == r_count_5_io_out ? io_r_421_b : _GEN_4260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4262 = 10'h1a6 == r_count_5_io_out ? io_r_422_b : _GEN_4261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4263 = 10'h1a7 == r_count_5_io_out ? io_r_423_b : _GEN_4262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4264 = 10'h1a8 == r_count_5_io_out ? io_r_424_b : _GEN_4263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4265 = 10'h1a9 == r_count_5_io_out ? io_r_425_b : _GEN_4264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4266 = 10'h1aa == r_count_5_io_out ? io_r_426_b : _GEN_4265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4267 = 10'h1ab == r_count_5_io_out ? io_r_427_b : _GEN_4266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4268 = 10'h1ac == r_count_5_io_out ? io_r_428_b : _GEN_4267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4269 = 10'h1ad == r_count_5_io_out ? io_r_429_b : _GEN_4268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4270 = 10'h1ae == r_count_5_io_out ? io_r_430_b : _GEN_4269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4271 = 10'h1af == r_count_5_io_out ? io_r_431_b : _GEN_4270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4272 = 10'h1b0 == r_count_5_io_out ? io_r_432_b : _GEN_4271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4273 = 10'h1b1 == r_count_5_io_out ? io_r_433_b : _GEN_4272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4274 = 10'h1b2 == r_count_5_io_out ? io_r_434_b : _GEN_4273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4275 = 10'h1b3 == r_count_5_io_out ? io_r_435_b : _GEN_4274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4276 = 10'h1b4 == r_count_5_io_out ? io_r_436_b : _GEN_4275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4277 = 10'h1b5 == r_count_5_io_out ? io_r_437_b : _GEN_4276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4278 = 10'h1b6 == r_count_5_io_out ? io_r_438_b : _GEN_4277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4279 = 10'h1b7 == r_count_5_io_out ? io_r_439_b : _GEN_4278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4280 = 10'h1b8 == r_count_5_io_out ? io_r_440_b : _GEN_4279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4281 = 10'h1b9 == r_count_5_io_out ? io_r_441_b : _GEN_4280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4282 = 10'h1ba == r_count_5_io_out ? io_r_442_b : _GEN_4281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4283 = 10'h1bb == r_count_5_io_out ? io_r_443_b : _GEN_4282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4284 = 10'h1bc == r_count_5_io_out ? io_r_444_b : _GEN_4283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4285 = 10'h1bd == r_count_5_io_out ? io_r_445_b : _GEN_4284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4286 = 10'h1be == r_count_5_io_out ? io_r_446_b : _GEN_4285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4287 = 10'h1bf == r_count_5_io_out ? io_r_447_b : _GEN_4286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4288 = 10'h1c0 == r_count_5_io_out ? io_r_448_b : _GEN_4287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4289 = 10'h1c1 == r_count_5_io_out ? io_r_449_b : _GEN_4288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4290 = 10'h1c2 == r_count_5_io_out ? io_r_450_b : _GEN_4289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4291 = 10'h1c3 == r_count_5_io_out ? io_r_451_b : _GEN_4290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4292 = 10'h1c4 == r_count_5_io_out ? io_r_452_b : _GEN_4291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4293 = 10'h1c5 == r_count_5_io_out ? io_r_453_b : _GEN_4292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4294 = 10'h1c6 == r_count_5_io_out ? io_r_454_b : _GEN_4293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4295 = 10'h1c7 == r_count_5_io_out ? io_r_455_b : _GEN_4294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4296 = 10'h1c8 == r_count_5_io_out ? io_r_456_b : _GEN_4295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4297 = 10'h1c9 == r_count_5_io_out ? io_r_457_b : _GEN_4296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4298 = 10'h1ca == r_count_5_io_out ? io_r_458_b : _GEN_4297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4299 = 10'h1cb == r_count_5_io_out ? io_r_459_b : _GEN_4298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4300 = 10'h1cc == r_count_5_io_out ? io_r_460_b : _GEN_4299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4301 = 10'h1cd == r_count_5_io_out ? io_r_461_b : _GEN_4300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4302 = 10'h1ce == r_count_5_io_out ? io_r_462_b : _GEN_4301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4303 = 10'h1cf == r_count_5_io_out ? io_r_463_b : _GEN_4302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4304 = 10'h1d0 == r_count_5_io_out ? io_r_464_b : _GEN_4303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4305 = 10'h1d1 == r_count_5_io_out ? io_r_465_b : _GEN_4304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4306 = 10'h1d2 == r_count_5_io_out ? io_r_466_b : _GEN_4305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4307 = 10'h1d3 == r_count_5_io_out ? io_r_467_b : _GEN_4306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4308 = 10'h1d4 == r_count_5_io_out ? io_r_468_b : _GEN_4307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4309 = 10'h1d5 == r_count_5_io_out ? io_r_469_b : _GEN_4308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4310 = 10'h1d6 == r_count_5_io_out ? io_r_470_b : _GEN_4309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4311 = 10'h1d7 == r_count_5_io_out ? io_r_471_b : _GEN_4310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4312 = 10'h1d8 == r_count_5_io_out ? io_r_472_b : _GEN_4311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4313 = 10'h1d9 == r_count_5_io_out ? io_r_473_b : _GEN_4312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4314 = 10'h1da == r_count_5_io_out ? io_r_474_b : _GEN_4313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4315 = 10'h1db == r_count_5_io_out ? io_r_475_b : _GEN_4314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4316 = 10'h1dc == r_count_5_io_out ? io_r_476_b : _GEN_4315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4317 = 10'h1dd == r_count_5_io_out ? io_r_477_b : _GEN_4316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4318 = 10'h1de == r_count_5_io_out ? io_r_478_b : _GEN_4317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4319 = 10'h1df == r_count_5_io_out ? io_r_479_b : _GEN_4318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4320 = 10'h1e0 == r_count_5_io_out ? io_r_480_b : _GEN_4319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4321 = 10'h1e1 == r_count_5_io_out ? io_r_481_b : _GEN_4320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4322 = 10'h1e2 == r_count_5_io_out ? io_r_482_b : _GEN_4321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4323 = 10'h1e3 == r_count_5_io_out ? io_r_483_b : _GEN_4322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4324 = 10'h1e4 == r_count_5_io_out ? io_r_484_b : _GEN_4323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4325 = 10'h1e5 == r_count_5_io_out ? io_r_485_b : _GEN_4324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4326 = 10'h1e6 == r_count_5_io_out ? io_r_486_b : _GEN_4325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4327 = 10'h1e7 == r_count_5_io_out ? io_r_487_b : _GEN_4326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4328 = 10'h1e8 == r_count_5_io_out ? io_r_488_b : _GEN_4327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4329 = 10'h1e9 == r_count_5_io_out ? io_r_489_b : _GEN_4328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4330 = 10'h1ea == r_count_5_io_out ? io_r_490_b : _GEN_4329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4331 = 10'h1eb == r_count_5_io_out ? io_r_491_b : _GEN_4330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4332 = 10'h1ec == r_count_5_io_out ? io_r_492_b : _GEN_4331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4333 = 10'h1ed == r_count_5_io_out ? io_r_493_b : _GEN_4332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4334 = 10'h1ee == r_count_5_io_out ? io_r_494_b : _GEN_4333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4335 = 10'h1ef == r_count_5_io_out ? io_r_495_b : _GEN_4334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4336 = 10'h1f0 == r_count_5_io_out ? io_r_496_b : _GEN_4335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4337 = 10'h1f1 == r_count_5_io_out ? io_r_497_b : _GEN_4336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4338 = 10'h1f2 == r_count_5_io_out ? io_r_498_b : _GEN_4337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4339 = 10'h1f3 == r_count_5_io_out ? io_r_499_b : _GEN_4338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4340 = 10'h1f4 == r_count_5_io_out ? io_r_500_b : _GEN_4339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4341 = 10'h1f5 == r_count_5_io_out ? io_r_501_b : _GEN_4340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4342 = 10'h1f6 == r_count_5_io_out ? io_r_502_b : _GEN_4341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4343 = 10'h1f7 == r_count_5_io_out ? io_r_503_b : _GEN_4342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4344 = 10'h1f8 == r_count_5_io_out ? io_r_504_b : _GEN_4343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4345 = 10'h1f9 == r_count_5_io_out ? io_r_505_b : _GEN_4344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4346 = 10'h1fa == r_count_5_io_out ? io_r_506_b : _GEN_4345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4347 = 10'h1fb == r_count_5_io_out ? io_r_507_b : _GEN_4346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4348 = 10'h1fc == r_count_5_io_out ? io_r_508_b : _GEN_4347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4349 = 10'h1fd == r_count_5_io_out ? io_r_509_b : _GEN_4348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4350 = 10'h1fe == r_count_5_io_out ? io_r_510_b : _GEN_4349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4351 = 10'h1ff == r_count_5_io_out ? io_r_511_b : _GEN_4350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4352 = 10'h200 == r_count_5_io_out ? io_r_512_b : _GEN_4351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4353 = 10'h201 == r_count_5_io_out ? io_r_513_b : _GEN_4352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4354 = 10'h202 == r_count_5_io_out ? io_r_514_b : _GEN_4353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4355 = 10'h203 == r_count_5_io_out ? io_r_515_b : _GEN_4354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4356 = 10'h204 == r_count_5_io_out ? io_r_516_b : _GEN_4355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4357 = 10'h205 == r_count_5_io_out ? io_r_517_b : _GEN_4356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4358 = 10'h206 == r_count_5_io_out ? io_r_518_b : _GEN_4357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4359 = 10'h207 == r_count_5_io_out ? io_r_519_b : _GEN_4358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4360 = 10'h208 == r_count_5_io_out ? io_r_520_b : _GEN_4359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4361 = 10'h209 == r_count_5_io_out ? io_r_521_b : _GEN_4360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4362 = 10'h20a == r_count_5_io_out ? io_r_522_b : _GEN_4361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4363 = 10'h20b == r_count_5_io_out ? io_r_523_b : _GEN_4362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4364 = 10'h20c == r_count_5_io_out ? io_r_524_b : _GEN_4363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4365 = 10'h20d == r_count_5_io_out ? io_r_525_b : _GEN_4364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4366 = 10'h20e == r_count_5_io_out ? io_r_526_b : _GEN_4365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4367 = 10'h20f == r_count_5_io_out ? io_r_527_b : _GEN_4366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4368 = 10'h210 == r_count_5_io_out ? io_r_528_b : _GEN_4367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4369 = 10'h211 == r_count_5_io_out ? io_r_529_b : _GEN_4368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4370 = 10'h212 == r_count_5_io_out ? io_r_530_b : _GEN_4369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4371 = 10'h213 == r_count_5_io_out ? io_r_531_b : _GEN_4370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4372 = 10'h214 == r_count_5_io_out ? io_r_532_b : _GEN_4371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4373 = 10'h215 == r_count_5_io_out ? io_r_533_b : _GEN_4372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4374 = 10'h216 == r_count_5_io_out ? io_r_534_b : _GEN_4373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4375 = 10'h217 == r_count_5_io_out ? io_r_535_b : _GEN_4374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4376 = 10'h218 == r_count_5_io_out ? io_r_536_b : _GEN_4375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4377 = 10'h219 == r_count_5_io_out ? io_r_537_b : _GEN_4376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4378 = 10'h21a == r_count_5_io_out ? io_r_538_b : _GEN_4377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4379 = 10'h21b == r_count_5_io_out ? io_r_539_b : _GEN_4378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4380 = 10'h21c == r_count_5_io_out ? io_r_540_b : _GEN_4379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4381 = 10'h21d == r_count_5_io_out ? io_r_541_b : _GEN_4380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4382 = 10'h21e == r_count_5_io_out ? io_r_542_b : _GEN_4381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4383 = 10'h21f == r_count_5_io_out ? io_r_543_b : _GEN_4382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4384 = 10'h220 == r_count_5_io_out ? io_r_544_b : _GEN_4383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4385 = 10'h221 == r_count_5_io_out ? io_r_545_b : _GEN_4384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4386 = 10'h222 == r_count_5_io_out ? io_r_546_b : _GEN_4385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4387 = 10'h223 == r_count_5_io_out ? io_r_547_b : _GEN_4386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4388 = 10'h224 == r_count_5_io_out ? io_r_548_b : _GEN_4387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4389 = 10'h225 == r_count_5_io_out ? io_r_549_b : _GEN_4388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4390 = 10'h226 == r_count_5_io_out ? io_r_550_b : _GEN_4389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4391 = 10'h227 == r_count_5_io_out ? io_r_551_b : _GEN_4390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4392 = 10'h228 == r_count_5_io_out ? io_r_552_b : _GEN_4391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4393 = 10'h229 == r_count_5_io_out ? io_r_553_b : _GEN_4392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4394 = 10'h22a == r_count_5_io_out ? io_r_554_b : _GEN_4393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4395 = 10'h22b == r_count_5_io_out ? io_r_555_b : _GEN_4394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4396 = 10'h22c == r_count_5_io_out ? io_r_556_b : _GEN_4395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4397 = 10'h22d == r_count_5_io_out ? io_r_557_b : _GEN_4396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4398 = 10'h22e == r_count_5_io_out ? io_r_558_b : _GEN_4397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4399 = 10'h22f == r_count_5_io_out ? io_r_559_b : _GEN_4398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4400 = 10'h230 == r_count_5_io_out ? io_r_560_b : _GEN_4399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4401 = 10'h231 == r_count_5_io_out ? io_r_561_b : _GEN_4400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4402 = 10'h232 == r_count_5_io_out ? io_r_562_b : _GEN_4401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4403 = 10'h233 == r_count_5_io_out ? io_r_563_b : _GEN_4402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4404 = 10'h234 == r_count_5_io_out ? io_r_564_b : _GEN_4403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4405 = 10'h235 == r_count_5_io_out ? io_r_565_b : _GEN_4404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4406 = 10'h236 == r_count_5_io_out ? io_r_566_b : _GEN_4405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4407 = 10'h237 == r_count_5_io_out ? io_r_567_b : _GEN_4406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4408 = 10'h238 == r_count_5_io_out ? io_r_568_b : _GEN_4407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4409 = 10'h239 == r_count_5_io_out ? io_r_569_b : _GEN_4408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4410 = 10'h23a == r_count_5_io_out ? io_r_570_b : _GEN_4409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4411 = 10'h23b == r_count_5_io_out ? io_r_571_b : _GEN_4410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4412 = 10'h23c == r_count_5_io_out ? io_r_572_b : _GEN_4411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4413 = 10'h23d == r_count_5_io_out ? io_r_573_b : _GEN_4412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4414 = 10'h23e == r_count_5_io_out ? io_r_574_b : _GEN_4413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4415 = 10'h23f == r_count_5_io_out ? io_r_575_b : _GEN_4414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4416 = 10'h240 == r_count_5_io_out ? io_r_576_b : _GEN_4415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4417 = 10'h241 == r_count_5_io_out ? io_r_577_b : _GEN_4416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4418 = 10'h242 == r_count_5_io_out ? io_r_578_b : _GEN_4417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4419 = 10'h243 == r_count_5_io_out ? io_r_579_b : _GEN_4418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4420 = 10'h244 == r_count_5_io_out ? io_r_580_b : _GEN_4419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4421 = 10'h245 == r_count_5_io_out ? io_r_581_b : _GEN_4420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4422 = 10'h246 == r_count_5_io_out ? io_r_582_b : _GEN_4421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4423 = 10'h247 == r_count_5_io_out ? io_r_583_b : _GEN_4422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4424 = 10'h248 == r_count_5_io_out ? io_r_584_b : _GEN_4423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4425 = 10'h249 == r_count_5_io_out ? io_r_585_b : _GEN_4424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4426 = 10'h24a == r_count_5_io_out ? io_r_586_b : _GEN_4425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4427 = 10'h24b == r_count_5_io_out ? io_r_587_b : _GEN_4426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4428 = 10'h24c == r_count_5_io_out ? io_r_588_b : _GEN_4427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4429 = 10'h24d == r_count_5_io_out ? io_r_589_b : _GEN_4428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4430 = 10'h24e == r_count_5_io_out ? io_r_590_b : _GEN_4429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4431 = 10'h24f == r_count_5_io_out ? io_r_591_b : _GEN_4430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4432 = 10'h250 == r_count_5_io_out ? io_r_592_b : _GEN_4431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4433 = 10'h251 == r_count_5_io_out ? io_r_593_b : _GEN_4432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4434 = 10'h252 == r_count_5_io_out ? io_r_594_b : _GEN_4433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4435 = 10'h253 == r_count_5_io_out ? io_r_595_b : _GEN_4434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4436 = 10'h254 == r_count_5_io_out ? io_r_596_b : _GEN_4435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4437 = 10'h255 == r_count_5_io_out ? io_r_597_b : _GEN_4436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4438 = 10'h256 == r_count_5_io_out ? io_r_598_b : _GEN_4437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4439 = 10'h257 == r_count_5_io_out ? io_r_599_b : _GEN_4438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4440 = 10'h258 == r_count_5_io_out ? io_r_600_b : _GEN_4439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4441 = 10'h259 == r_count_5_io_out ? io_r_601_b : _GEN_4440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4442 = 10'h25a == r_count_5_io_out ? io_r_602_b : _GEN_4441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4443 = 10'h25b == r_count_5_io_out ? io_r_603_b : _GEN_4442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4444 = 10'h25c == r_count_5_io_out ? io_r_604_b : _GEN_4443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4445 = 10'h25d == r_count_5_io_out ? io_r_605_b : _GEN_4444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4446 = 10'h25e == r_count_5_io_out ? io_r_606_b : _GEN_4445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4447 = 10'h25f == r_count_5_io_out ? io_r_607_b : _GEN_4446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4448 = 10'h260 == r_count_5_io_out ? io_r_608_b : _GEN_4447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4449 = 10'h261 == r_count_5_io_out ? io_r_609_b : _GEN_4448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4450 = 10'h262 == r_count_5_io_out ? io_r_610_b : _GEN_4449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4451 = 10'h263 == r_count_5_io_out ? io_r_611_b : _GEN_4450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4452 = 10'h264 == r_count_5_io_out ? io_r_612_b : _GEN_4451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4453 = 10'h265 == r_count_5_io_out ? io_r_613_b : _GEN_4452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4454 = 10'h266 == r_count_5_io_out ? io_r_614_b : _GEN_4453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4455 = 10'h267 == r_count_5_io_out ? io_r_615_b : _GEN_4454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4456 = 10'h268 == r_count_5_io_out ? io_r_616_b : _GEN_4455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4457 = 10'h269 == r_count_5_io_out ? io_r_617_b : _GEN_4456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4458 = 10'h26a == r_count_5_io_out ? io_r_618_b : _GEN_4457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4459 = 10'h26b == r_count_5_io_out ? io_r_619_b : _GEN_4458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4460 = 10'h26c == r_count_5_io_out ? io_r_620_b : _GEN_4459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4461 = 10'h26d == r_count_5_io_out ? io_r_621_b : _GEN_4460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4462 = 10'h26e == r_count_5_io_out ? io_r_622_b : _GEN_4461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4463 = 10'h26f == r_count_5_io_out ? io_r_623_b : _GEN_4462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4464 = 10'h270 == r_count_5_io_out ? io_r_624_b : _GEN_4463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4465 = 10'h271 == r_count_5_io_out ? io_r_625_b : _GEN_4464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4466 = 10'h272 == r_count_5_io_out ? io_r_626_b : _GEN_4465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4467 = 10'h273 == r_count_5_io_out ? io_r_627_b : _GEN_4466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4468 = 10'h274 == r_count_5_io_out ? io_r_628_b : _GEN_4467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4469 = 10'h275 == r_count_5_io_out ? io_r_629_b : _GEN_4468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4470 = 10'h276 == r_count_5_io_out ? io_r_630_b : _GEN_4469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4471 = 10'h277 == r_count_5_io_out ? io_r_631_b : _GEN_4470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4472 = 10'h278 == r_count_5_io_out ? io_r_632_b : _GEN_4471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4473 = 10'h279 == r_count_5_io_out ? io_r_633_b : _GEN_4472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4474 = 10'h27a == r_count_5_io_out ? io_r_634_b : _GEN_4473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4475 = 10'h27b == r_count_5_io_out ? io_r_635_b : _GEN_4474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4476 = 10'h27c == r_count_5_io_out ? io_r_636_b : _GEN_4475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4477 = 10'h27d == r_count_5_io_out ? io_r_637_b : _GEN_4476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4478 = 10'h27e == r_count_5_io_out ? io_r_638_b : _GEN_4477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4479 = 10'h27f == r_count_5_io_out ? io_r_639_b : _GEN_4478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4480 = 10'h280 == r_count_5_io_out ? io_r_640_b : _GEN_4479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4481 = 10'h281 == r_count_5_io_out ? io_r_641_b : _GEN_4480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4482 = 10'h282 == r_count_5_io_out ? io_r_642_b : _GEN_4481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4483 = 10'h283 == r_count_5_io_out ? io_r_643_b : _GEN_4482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4484 = 10'h284 == r_count_5_io_out ? io_r_644_b : _GEN_4483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4485 = 10'h285 == r_count_5_io_out ? io_r_645_b : _GEN_4484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4486 = 10'h286 == r_count_5_io_out ? io_r_646_b : _GEN_4485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4487 = 10'h287 == r_count_5_io_out ? io_r_647_b : _GEN_4486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4488 = 10'h288 == r_count_5_io_out ? io_r_648_b : _GEN_4487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4489 = 10'h289 == r_count_5_io_out ? io_r_649_b : _GEN_4488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4490 = 10'h28a == r_count_5_io_out ? io_r_650_b : _GEN_4489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4491 = 10'h28b == r_count_5_io_out ? io_r_651_b : _GEN_4490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4492 = 10'h28c == r_count_5_io_out ? io_r_652_b : _GEN_4491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4493 = 10'h28d == r_count_5_io_out ? io_r_653_b : _GEN_4492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4494 = 10'h28e == r_count_5_io_out ? io_r_654_b : _GEN_4493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4495 = 10'h28f == r_count_5_io_out ? io_r_655_b : _GEN_4494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4496 = 10'h290 == r_count_5_io_out ? io_r_656_b : _GEN_4495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4497 = 10'h291 == r_count_5_io_out ? io_r_657_b : _GEN_4496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4498 = 10'h292 == r_count_5_io_out ? io_r_658_b : _GEN_4497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4499 = 10'h293 == r_count_5_io_out ? io_r_659_b : _GEN_4498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4500 = 10'h294 == r_count_5_io_out ? io_r_660_b : _GEN_4499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4501 = 10'h295 == r_count_5_io_out ? io_r_661_b : _GEN_4500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4502 = 10'h296 == r_count_5_io_out ? io_r_662_b : _GEN_4501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4503 = 10'h297 == r_count_5_io_out ? io_r_663_b : _GEN_4502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4504 = 10'h298 == r_count_5_io_out ? io_r_664_b : _GEN_4503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4505 = 10'h299 == r_count_5_io_out ? io_r_665_b : _GEN_4504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4506 = 10'h29a == r_count_5_io_out ? io_r_666_b : _GEN_4505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4507 = 10'h29b == r_count_5_io_out ? io_r_667_b : _GEN_4506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4508 = 10'h29c == r_count_5_io_out ? io_r_668_b : _GEN_4507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4509 = 10'h29d == r_count_5_io_out ? io_r_669_b : _GEN_4508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4510 = 10'h29e == r_count_5_io_out ? io_r_670_b : _GEN_4509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4511 = 10'h29f == r_count_5_io_out ? io_r_671_b : _GEN_4510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4512 = 10'h2a0 == r_count_5_io_out ? io_r_672_b : _GEN_4511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4513 = 10'h2a1 == r_count_5_io_out ? io_r_673_b : _GEN_4512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4514 = 10'h2a2 == r_count_5_io_out ? io_r_674_b : _GEN_4513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4515 = 10'h2a3 == r_count_5_io_out ? io_r_675_b : _GEN_4514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4516 = 10'h2a4 == r_count_5_io_out ? io_r_676_b : _GEN_4515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4517 = 10'h2a5 == r_count_5_io_out ? io_r_677_b : _GEN_4516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4518 = 10'h2a6 == r_count_5_io_out ? io_r_678_b : _GEN_4517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4519 = 10'h2a7 == r_count_5_io_out ? io_r_679_b : _GEN_4518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4520 = 10'h2a8 == r_count_5_io_out ? io_r_680_b : _GEN_4519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4521 = 10'h2a9 == r_count_5_io_out ? io_r_681_b : _GEN_4520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4522 = 10'h2aa == r_count_5_io_out ? io_r_682_b : _GEN_4521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4523 = 10'h2ab == r_count_5_io_out ? io_r_683_b : _GEN_4522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4524 = 10'h2ac == r_count_5_io_out ? io_r_684_b : _GEN_4523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4525 = 10'h2ad == r_count_5_io_out ? io_r_685_b : _GEN_4524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4526 = 10'h2ae == r_count_5_io_out ? io_r_686_b : _GEN_4525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4527 = 10'h2af == r_count_5_io_out ? io_r_687_b : _GEN_4526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4528 = 10'h2b0 == r_count_5_io_out ? io_r_688_b : _GEN_4527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4529 = 10'h2b1 == r_count_5_io_out ? io_r_689_b : _GEN_4528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4530 = 10'h2b2 == r_count_5_io_out ? io_r_690_b : _GEN_4529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4531 = 10'h2b3 == r_count_5_io_out ? io_r_691_b : _GEN_4530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4532 = 10'h2b4 == r_count_5_io_out ? io_r_692_b : _GEN_4531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4533 = 10'h2b5 == r_count_5_io_out ? io_r_693_b : _GEN_4532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4534 = 10'h2b6 == r_count_5_io_out ? io_r_694_b : _GEN_4533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4535 = 10'h2b7 == r_count_5_io_out ? io_r_695_b : _GEN_4534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4536 = 10'h2b8 == r_count_5_io_out ? io_r_696_b : _GEN_4535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4537 = 10'h2b9 == r_count_5_io_out ? io_r_697_b : _GEN_4536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4538 = 10'h2ba == r_count_5_io_out ? io_r_698_b : _GEN_4537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4539 = 10'h2bb == r_count_5_io_out ? io_r_699_b : _GEN_4538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4540 = 10'h2bc == r_count_5_io_out ? io_r_700_b : _GEN_4539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4541 = 10'h2bd == r_count_5_io_out ? io_r_701_b : _GEN_4540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4542 = 10'h2be == r_count_5_io_out ? io_r_702_b : _GEN_4541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4543 = 10'h2bf == r_count_5_io_out ? io_r_703_b : _GEN_4542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4544 = 10'h2c0 == r_count_5_io_out ? io_r_704_b : _GEN_4543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4545 = 10'h2c1 == r_count_5_io_out ? io_r_705_b : _GEN_4544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4546 = 10'h2c2 == r_count_5_io_out ? io_r_706_b : _GEN_4545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4547 = 10'h2c3 == r_count_5_io_out ? io_r_707_b : _GEN_4546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4548 = 10'h2c4 == r_count_5_io_out ? io_r_708_b : _GEN_4547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4549 = 10'h2c5 == r_count_5_io_out ? io_r_709_b : _GEN_4548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4550 = 10'h2c6 == r_count_5_io_out ? io_r_710_b : _GEN_4549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4551 = 10'h2c7 == r_count_5_io_out ? io_r_711_b : _GEN_4550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4552 = 10'h2c8 == r_count_5_io_out ? io_r_712_b : _GEN_4551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4553 = 10'h2c9 == r_count_5_io_out ? io_r_713_b : _GEN_4552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4554 = 10'h2ca == r_count_5_io_out ? io_r_714_b : _GEN_4553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4555 = 10'h2cb == r_count_5_io_out ? io_r_715_b : _GEN_4554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4556 = 10'h2cc == r_count_5_io_out ? io_r_716_b : _GEN_4555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4557 = 10'h2cd == r_count_5_io_out ? io_r_717_b : _GEN_4556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4558 = 10'h2ce == r_count_5_io_out ? io_r_718_b : _GEN_4557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4559 = 10'h2cf == r_count_5_io_out ? io_r_719_b : _GEN_4558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4560 = 10'h2d0 == r_count_5_io_out ? io_r_720_b : _GEN_4559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4561 = 10'h2d1 == r_count_5_io_out ? io_r_721_b : _GEN_4560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4562 = 10'h2d2 == r_count_5_io_out ? io_r_722_b : _GEN_4561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4563 = 10'h2d3 == r_count_5_io_out ? io_r_723_b : _GEN_4562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4564 = 10'h2d4 == r_count_5_io_out ? io_r_724_b : _GEN_4563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4565 = 10'h2d5 == r_count_5_io_out ? io_r_725_b : _GEN_4564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4566 = 10'h2d6 == r_count_5_io_out ? io_r_726_b : _GEN_4565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4567 = 10'h2d7 == r_count_5_io_out ? io_r_727_b : _GEN_4566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4568 = 10'h2d8 == r_count_5_io_out ? io_r_728_b : _GEN_4567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4569 = 10'h2d9 == r_count_5_io_out ? io_r_729_b : _GEN_4568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4570 = 10'h2da == r_count_5_io_out ? io_r_730_b : _GEN_4569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4571 = 10'h2db == r_count_5_io_out ? io_r_731_b : _GEN_4570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4572 = 10'h2dc == r_count_5_io_out ? io_r_732_b : _GEN_4571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4573 = 10'h2dd == r_count_5_io_out ? io_r_733_b : _GEN_4572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4574 = 10'h2de == r_count_5_io_out ? io_r_734_b : _GEN_4573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4575 = 10'h2df == r_count_5_io_out ? io_r_735_b : _GEN_4574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4576 = 10'h2e0 == r_count_5_io_out ? io_r_736_b : _GEN_4575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4577 = 10'h2e1 == r_count_5_io_out ? io_r_737_b : _GEN_4576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4578 = 10'h2e2 == r_count_5_io_out ? io_r_738_b : _GEN_4577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4579 = 10'h2e3 == r_count_5_io_out ? io_r_739_b : _GEN_4578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4580 = 10'h2e4 == r_count_5_io_out ? io_r_740_b : _GEN_4579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4581 = 10'h2e5 == r_count_5_io_out ? io_r_741_b : _GEN_4580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4582 = 10'h2e6 == r_count_5_io_out ? io_r_742_b : _GEN_4581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4583 = 10'h2e7 == r_count_5_io_out ? io_r_743_b : _GEN_4582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4584 = 10'h2e8 == r_count_5_io_out ? io_r_744_b : _GEN_4583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4585 = 10'h2e9 == r_count_5_io_out ? io_r_745_b : _GEN_4584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4586 = 10'h2ea == r_count_5_io_out ? io_r_746_b : _GEN_4585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4587 = 10'h2eb == r_count_5_io_out ? io_r_747_b : _GEN_4586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4588 = 10'h2ec == r_count_5_io_out ? io_r_748_b : _GEN_4587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4591 = 10'h1 == r_count_6_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4592 = 10'h2 == r_count_6_io_out ? io_r_2_b : _GEN_4591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4593 = 10'h3 == r_count_6_io_out ? io_r_3_b : _GEN_4592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4594 = 10'h4 == r_count_6_io_out ? io_r_4_b : _GEN_4593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4595 = 10'h5 == r_count_6_io_out ? io_r_5_b : _GEN_4594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4596 = 10'h6 == r_count_6_io_out ? io_r_6_b : _GEN_4595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4597 = 10'h7 == r_count_6_io_out ? io_r_7_b : _GEN_4596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4598 = 10'h8 == r_count_6_io_out ? io_r_8_b : _GEN_4597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4599 = 10'h9 == r_count_6_io_out ? io_r_9_b : _GEN_4598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4600 = 10'ha == r_count_6_io_out ? io_r_10_b : _GEN_4599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4601 = 10'hb == r_count_6_io_out ? io_r_11_b : _GEN_4600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4602 = 10'hc == r_count_6_io_out ? io_r_12_b : _GEN_4601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4603 = 10'hd == r_count_6_io_out ? io_r_13_b : _GEN_4602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4604 = 10'he == r_count_6_io_out ? io_r_14_b : _GEN_4603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4605 = 10'hf == r_count_6_io_out ? io_r_15_b : _GEN_4604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4606 = 10'h10 == r_count_6_io_out ? io_r_16_b : _GEN_4605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4607 = 10'h11 == r_count_6_io_out ? io_r_17_b : _GEN_4606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4608 = 10'h12 == r_count_6_io_out ? io_r_18_b : _GEN_4607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4609 = 10'h13 == r_count_6_io_out ? io_r_19_b : _GEN_4608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4610 = 10'h14 == r_count_6_io_out ? io_r_20_b : _GEN_4609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4611 = 10'h15 == r_count_6_io_out ? io_r_21_b : _GEN_4610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4612 = 10'h16 == r_count_6_io_out ? io_r_22_b : _GEN_4611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4613 = 10'h17 == r_count_6_io_out ? io_r_23_b : _GEN_4612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4614 = 10'h18 == r_count_6_io_out ? io_r_24_b : _GEN_4613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4615 = 10'h19 == r_count_6_io_out ? io_r_25_b : _GEN_4614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4616 = 10'h1a == r_count_6_io_out ? io_r_26_b : _GEN_4615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4617 = 10'h1b == r_count_6_io_out ? io_r_27_b : _GEN_4616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4618 = 10'h1c == r_count_6_io_out ? io_r_28_b : _GEN_4617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4619 = 10'h1d == r_count_6_io_out ? io_r_29_b : _GEN_4618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4620 = 10'h1e == r_count_6_io_out ? io_r_30_b : _GEN_4619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4621 = 10'h1f == r_count_6_io_out ? io_r_31_b : _GEN_4620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4622 = 10'h20 == r_count_6_io_out ? io_r_32_b : _GEN_4621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4623 = 10'h21 == r_count_6_io_out ? io_r_33_b : _GEN_4622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4624 = 10'h22 == r_count_6_io_out ? io_r_34_b : _GEN_4623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4625 = 10'h23 == r_count_6_io_out ? io_r_35_b : _GEN_4624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4626 = 10'h24 == r_count_6_io_out ? io_r_36_b : _GEN_4625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4627 = 10'h25 == r_count_6_io_out ? io_r_37_b : _GEN_4626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4628 = 10'h26 == r_count_6_io_out ? io_r_38_b : _GEN_4627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4629 = 10'h27 == r_count_6_io_out ? io_r_39_b : _GEN_4628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4630 = 10'h28 == r_count_6_io_out ? io_r_40_b : _GEN_4629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4631 = 10'h29 == r_count_6_io_out ? io_r_41_b : _GEN_4630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4632 = 10'h2a == r_count_6_io_out ? io_r_42_b : _GEN_4631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4633 = 10'h2b == r_count_6_io_out ? io_r_43_b : _GEN_4632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4634 = 10'h2c == r_count_6_io_out ? io_r_44_b : _GEN_4633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4635 = 10'h2d == r_count_6_io_out ? io_r_45_b : _GEN_4634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4636 = 10'h2e == r_count_6_io_out ? io_r_46_b : _GEN_4635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4637 = 10'h2f == r_count_6_io_out ? io_r_47_b : _GEN_4636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4638 = 10'h30 == r_count_6_io_out ? io_r_48_b : _GEN_4637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4639 = 10'h31 == r_count_6_io_out ? io_r_49_b : _GEN_4638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4640 = 10'h32 == r_count_6_io_out ? io_r_50_b : _GEN_4639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4641 = 10'h33 == r_count_6_io_out ? io_r_51_b : _GEN_4640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4642 = 10'h34 == r_count_6_io_out ? io_r_52_b : _GEN_4641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4643 = 10'h35 == r_count_6_io_out ? io_r_53_b : _GEN_4642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4644 = 10'h36 == r_count_6_io_out ? io_r_54_b : _GEN_4643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4645 = 10'h37 == r_count_6_io_out ? io_r_55_b : _GEN_4644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4646 = 10'h38 == r_count_6_io_out ? io_r_56_b : _GEN_4645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4647 = 10'h39 == r_count_6_io_out ? io_r_57_b : _GEN_4646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4648 = 10'h3a == r_count_6_io_out ? io_r_58_b : _GEN_4647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4649 = 10'h3b == r_count_6_io_out ? io_r_59_b : _GEN_4648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4650 = 10'h3c == r_count_6_io_out ? io_r_60_b : _GEN_4649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4651 = 10'h3d == r_count_6_io_out ? io_r_61_b : _GEN_4650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4652 = 10'h3e == r_count_6_io_out ? io_r_62_b : _GEN_4651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4653 = 10'h3f == r_count_6_io_out ? io_r_63_b : _GEN_4652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4654 = 10'h40 == r_count_6_io_out ? io_r_64_b : _GEN_4653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4655 = 10'h41 == r_count_6_io_out ? io_r_65_b : _GEN_4654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4656 = 10'h42 == r_count_6_io_out ? io_r_66_b : _GEN_4655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4657 = 10'h43 == r_count_6_io_out ? io_r_67_b : _GEN_4656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4658 = 10'h44 == r_count_6_io_out ? io_r_68_b : _GEN_4657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4659 = 10'h45 == r_count_6_io_out ? io_r_69_b : _GEN_4658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4660 = 10'h46 == r_count_6_io_out ? io_r_70_b : _GEN_4659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4661 = 10'h47 == r_count_6_io_out ? io_r_71_b : _GEN_4660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4662 = 10'h48 == r_count_6_io_out ? io_r_72_b : _GEN_4661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4663 = 10'h49 == r_count_6_io_out ? io_r_73_b : _GEN_4662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4664 = 10'h4a == r_count_6_io_out ? io_r_74_b : _GEN_4663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4665 = 10'h4b == r_count_6_io_out ? io_r_75_b : _GEN_4664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4666 = 10'h4c == r_count_6_io_out ? io_r_76_b : _GEN_4665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4667 = 10'h4d == r_count_6_io_out ? io_r_77_b : _GEN_4666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4668 = 10'h4e == r_count_6_io_out ? io_r_78_b : _GEN_4667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4669 = 10'h4f == r_count_6_io_out ? io_r_79_b : _GEN_4668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4670 = 10'h50 == r_count_6_io_out ? io_r_80_b : _GEN_4669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4671 = 10'h51 == r_count_6_io_out ? io_r_81_b : _GEN_4670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4672 = 10'h52 == r_count_6_io_out ? io_r_82_b : _GEN_4671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4673 = 10'h53 == r_count_6_io_out ? io_r_83_b : _GEN_4672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4674 = 10'h54 == r_count_6_io_out ? io_r_84_b : _GEN_4673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4675 = 10'h55 == r_count_6_io_out ? io_r_85_b : _GEN_4674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4676 = 10'h56 == r_count_6_io_out ? io_r_86_b : _GEN_4675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4677 = 10'h57 == r_count_6_io_out ? io_r_87_b : _GEN_4676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4678 = 10'h58 == r_count_6_io_out ? io_r_88_b : _GEN_4677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4679 = 10'h59 == r_count_6_io_out ? io_r_89_b : _GEN_4678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4680 = 10'h5a == r_count_6_io_out ? io_r_90_b : _GEN_4679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4681 = 10'h5b == r_count_6_io_out ? io_r_91_b : _GEN_4680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4682 = 10'h5c == r_count_6_io_out ? io_r_92_b : _GEN_4681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4683 = 10'h5d == r_count_6_io_out ? io_r_93_b : _GEN_4682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4684 = 10'h5e == r_count_6_io_out ? io_r_94_b : _GEN_4683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4685 = 10'h5f == r_count_6_io_out ? io_r_95_b : _GEN_4684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4686 = 10'h60 == r_count_6_io_out ? io_r_96_b : _GEN_4685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4687 = 10'h61 == r_count_6_io_out ? io_r_97_b : _GEN_4686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4688 = 10'h62 == r_count_6_io_out ? io_r_98_b : _GEN_4687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4689 = 10'h63 == r_count_6_io_out ? io_r_99_b : _GEN_4688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4690 = 10'h64 == r_count_6_io_out ? io_r_100_b : _GEN_4689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4691 = 10'h65 == r_count_6_io_out ? io_r_101_b : _GEN_4690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4692 = 10'h66 == r_count_6_io_out ? io_r_102_b : _GEN_4691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4693 = 10'h67 == r_count_6_io_out ? io_r_103_b : _GEN_4692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4694 = 10'h68 == r_count_6_io_out ? io_r_104_b : _GEN_4693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4695 = 10'h69 == r_count_6_io_out ? io_r_105_b : _GEN_4694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4696 = 10'h6a == r_count_6_io_out ? io_r_106_b : _GEN_4695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4697 = 10'h6b == r_count_6_io_out ? io_r_107_b : _GEN_4696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4698 = 10'h6c == r_count_6_io_out ? io_r_108_b : _GEN_4697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4699 = 10'h6d == r_count_6_io_out ? io_r_109_b : _GEN_4698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4700 = 10'h6e == r_count_6_io_out ? io_r_110_b : _GEN_4699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4701 = 10'h6f == r_count_6_io_out ? io_r_111_b : _GEN_4700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4702 = 10'h70 == r_count_6_io_out ? io_r_112_b : _GEN_4701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4703 = 10'h71 == r_count_6_io_out ? io_r_113_b : _GEN_4702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4704 = 10'h72 == r_count_6_io_out ? io_r_114_b : _GEN_4703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4705 = 10'h73 == r_count_6_io_out ? io_r_115_b : _GEN_4704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4706 = 10'h74 == r_count_6_io_out ? io_r_116_b : _GEN_4705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4707 = 10'h75 == r_count_6_io_out ? io_r_117_b : _GEN_4706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4708 = 10'h76 == r_count_6_io_out ? io_r_118_b : _GEN_4707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4709 = 10'h77 == r_count_6_io_out ? io_r_119_b : _GEN_4708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4710 = 10'h78 == r_count_6_io_out ? io_r_120_b : _GEN_4709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4711 = 10'h79 == r_count_6_io_out ? io_r_121_b : _GEN_4710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4712 = 10'h7a == r_count_6_io_out ? io_r_122_b : _GEN_4711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4713 = 10'h7b == r_count_6_io_out ? io_r_123_b : _GEN_4712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4714 = 10'h7c == r_count_6_io_out ? io_r_124_b : _GEN_4713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4715 = 10'h7d == r_count_6_io_out ? io_r_125_b : _GEN_4714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4716 = 10'h7e == r_count_6_io_out ? io_r_126_b : _GEN_4715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4717 = 10'h7f == r_count_6_io_out ? io_r_127_b : _GEN_4716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4718 = 10'h80 == r_count_6_io_out ? io_r_128_b : _GEN_4717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4719 = 10'h81 == r_count_6_io_out ? io_r_129_b : _GEN_4718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4720 = 10'h82 == r_count_6_io_out ? io_r_130_b : _GEN_4719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4721 = 10'h83 == r_count_6_io_out ? io_r_131_b : _GEN_4720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4722 = 10'h84 == r_count_6_io_out ? io_r_132_b : _GEN_4721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4723 = 10'h85 == r_count_6_io_out ? io_r_133_b : _GEN_4722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4724 = 10'h86 == r_count_6_io_out ? io_r_134_b : _GEN_4723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4725 = 10'h87 == r_count_6_io_out ? io_r_135_b : _GEN_4724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4726 = 10'h88 == r_count_6_io_out ? io_r_136_b : _GEN_4725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4727 = 10'h89 == r_count_6_io_out ? io_r_137_b : _GEN_4726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4728 = 10'h8a == r_count_6_io_out ? io_r_138_b : _GEN_4727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4729 = 10'h8b == r_count_6_io_out ? io_r_139_b : _GEN_4728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4730 = 10'h8c == r_count_6_io_out ? io_r_140_b : _GEN_4729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4731 = 10'h8d == r_count_6_io_out ? io_r_141_b : _GEN_4730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4732 = 10'h8e == r_count_6_io_out ? io_r_142_b : _GEN_4731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4733 = 10'h8f == r_count_6_io_out ? io_r_143_b : _GEN_4732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4734 = 10'h90 == r_count_6_io_out ? io_r_144_b : _GEN_4733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4735 = 10'h91 == r_count_6_io_out ? io_r_145_b : _GEN_4734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4736 = 10'h92 == r_count_6_io_out ? io_r_146_b : _GEN_4735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4737 = 10'h93 == r_count_6_io_out ? io_r_147_b : _GEN_4736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4738 = 10'h94 == r_count_6_io_out ? io_r_148_b : _GEN_4737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4739 = 10'h95 == r_count_6_io_out ? io_r_149_b : _GEN_4738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4740 = 10'h96 == r_count_6_io_out ? io_r_150_b : _GEN_4739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4741 = 10'h97 == r_count_6_io_out ? io_r_151_b : _GEN_4740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4742 = 10'h98 == r_count_6_io_out ? io_r_152_b : _GEN_4741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4743 = 10'h99 == r_count_6_io_out ? io_r_153_b : _GEN_4742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4744 = 10'h9a == r_count_6_io_out ? io_r_154_b : _GEN_4743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4745 = 10'h9b == r_count_6_io_out ? io_r_155_b : _GEN_4744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4746 = 10'h9c == r_count_6_io_out ? io_r_156_b : _GEN_4745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4747 = 10'h9d == r_count_6_io_out ? io_r_157_b : _GEN_4746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4748 = 10'h9e == r_count_6_io_out ? io_r_158_b : _GEN_4747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4749 = 10'h9f == r_count_6_io_out ? io_r_159_b : _GEN_4748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4750 = 10'ha0 == r_count_6_io_out ? io_r_160_b : _GEN_4749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4751 = 10'ha1 == r_count_6_io_out ? io_r_161_b : _GEN_4750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4752 = 10'ha2 == r_count_6_io_out ? io_r_162_b : _GEN_4751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4753 = 10'ha3 == r_count_6_io_out ? io_r_163_b : _GEN_4752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4754 = 10'ha4 == r_count_6_io_out ? io_r_164_b : _GEN_4753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4755 = 10'ha5 == r_count_6_io_out ? io_r_165_b : _GEN_4754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4756 = 10'ha6 == r_count_6_io_out ? io_r_166_b : _GEN_4755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4757 = 10'ha7 == r_count_6_io_out ? io_r_167_b : _GEN_4756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4758 = 10'ha8 == r_count_6_io_out ? io_r_168_b : _GEN_4757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4759 = 10'ha9 == r_count_6_io_out ? io_r_169_b : _GEN_4758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4760 = 10'haa == r_count_6_io_out ? io_r_170_b : _GEN_4759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4761 = 10'hab == r_count_6_io_out ? io_r_171_b : _GEN_4760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4762 = 10'hac == r_count_6_io_out ? io_r_172_b : _GEN_4761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4763 = 10'had == r_count_6_io_out ? io_r_173_b : _GEN_4762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4764 = 10'hae == r_count_6_io_out ? io_r_174_b : _GEN_4763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4765 = 10'haf == r_count_6_io_out ? io_r_175_b : _GEN_4764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4766 = 10'hb0 == r_count_6_io_out ? io_r_176_b : _GEN_4765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4767 = 10'hb1 == r_count_6_io_out ? io_r_177_b : _GEN_4766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4768 = 10'hb2 == r_count_6_io_out ? io_r_178_b : _GEN_4767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4769 = 10'hb3 == r_count_6_io_out ? io_r_179_b : _GEN_4768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4770 = 10'hb4 == r_count_6_io_out ? io_r_180_b : _GEN_4769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4771 = 10'hb5 == r_count_6_io_out ? io_r_181_b : _GEN_4770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4772 = 10'hb6 == r_count_6_io_out ? io_r_182_b : _GEN_4771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4773 = 10'hb7 == r_count_6_io_out ? io_r_183_b : _GEN_4772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4774 = 10'hb8 == r_count_6_io_out ? io_r_184_b : _GEN_4773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4775 = 10'hb9 == r_count_6_io_out ? io_r_185_b : _GEN_4774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4776 = 10'hba == r_count_6_io_out ? io_r_186_b : _GEN_4775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4777 = 10'hbb == r_count_6_io_out ? io_r_187_b : _GEN_4776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4778 = 10'hbc == r_count_6_io_out ? io_r_188_b : _GEN_4777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4779 = 10'hbd == r_count_6_io_out ? io_r_189_b : _GEN_4778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4780 = 10'hbe == r_count_6_io_out ? io_r_190_b : _GEN_4779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4781 = 10'hbf == r_count_6_io_out ? io_r_191_b : _GEN_4780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4782 = 10'hc0 == r_count_6_io_out ? io_r_192_b : _GEN_4781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4783 = 10'hc1 == r_count_6_io_out ? io_r_193_b : _GEN_4782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4784 = 10'hc2 == r_count_6_io_out ? io_r_194_b : _GEN_4783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4785 = 10'hc3 == r_count_6_io_out ? io_r_195_b : _GEN_4784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4786 = 10'hc4 == r_count_6_io_out ? io_r_196_b : _GEN_4785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4787 = 10'hc5 == r_count_6_io_out ? io_r_197_b : _GEN_4786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4788 = 10'hc6 == r_count_6_io_out ? io_r_198_b : _GEN_4787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4789 = 10'hc7 == r_count_6_io_out ? io_r_199_b : _GEN_4788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4790 = 10'hc8 == r_count_6_io_out ? io_r_200_b : _GEN_4789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4791 = 10'hc9 == r_count_6_io_out ? io_r_201_b : _GEN_4790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4792 = 10'hca == r_count_6_io_out ? io_r_202_b : _GEN_4791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4793 = 10'hcb == r_count_6_io_out ? io_r_203_b : _GEN_4792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4794 = 10'hcc == r_count_6_io_out ? io_r_204_b : _GEN_4793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4795 = 10'hcd == r_count_6_io_out ? io_r_205_b : _GEN_4794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4796 = 10'hce == r_count_6_io_out ? io_r_206_b : _GEN_4795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4797 = 10'hcf == r_count_6_io_out ? io_r_207_b : _GEN_4796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4798 = 10'hd0 == r_count_6_io_out ? io_r_208_b : _GEN_4797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4799 = 10'hd1 == r_count_6_io_out ? io_r_209_b : _GEN_4798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4800 = 10'hd2 == r_count_6_io_out ? io_r_210_b : _GEN_4799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4801 = 10'hd3 == r_count_6_io_out ? io_r_211_b : _GEN_4800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4802 = 10'hd4 == r_count_6_io_out ? io_r_212_b : _GEN_4801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4803 = 10'hd5 == r_count_6_io_out ? io_r_213_b : _GEN_4802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4804 = 10'hd6 == r_count_6_io_out ? io_r_214_b : _GEN_4803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4805 = 10'hd7 == r_count_6_io_out ? io_r_215_b : _GEN_4804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4806 = 10'hd8 == r_count_6_io_out ? io_r_216_b : _GEN_4805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4807 = 10'hd9 == r_count_6_io_out ? io_r_217_b : _GEN_4806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4808 = 10'hda == r_count_6_io_out ? io_r_218_b : _GEN_4807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4809 = 10'hdb == r_count_6_io_out ? io_r_219_b : _GEN_4808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4810 = 10'hdc == r_count_6_io_out ? io_r_220_b : _GEN_4809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4811 = 10'hdd == r_count_6_io_out ? io_r_221_b : _GEN_4810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4812 = 10'hde == r_count_6_io_out ? io_r_222_b : _GEN_4811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4813 = 10'hdf == r_count_6_io_out ? io_r_223_b : _GEN_4812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4814 = 10'he0 == r_count_6_io_out ? io_r_224_b : _GEN_4813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4815 = 10'he1 == r_count_6_io_out ? io_r_225_b : _GEN_4814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4816 = 10'he2 == r_count_6_io_out ? io_r_226_b : _GEN_4815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4817 = 10'he3 == r_count_6_io_out ? io_r_227_b : _GEN_4816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4818 = 10'he4 == r_count_6_io_out ? io_r_228_b : _GEN_4817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4819 = 10'he5 == r_count_6_io_out ? io_r_229_b : _GEN_4818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4820 = 10'he6 == r_count_6_io_out ? io_r_230_b : _GEN_4819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4821 = 10'he7 == r_count_6_io_out ? io_r_231_b : _GEN_4820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4822 = 10'he8 == r_count_6_io_out ? io_r_232_b : _GEN_4821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4823 = 10'he9 == r_count_6_io_out ? io_r_233_b : _GEN_4822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4824 = 10'hea == r_count_6_io_out ? io_r_234_b : _GEN_4823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4825 = 10'heb == r_count_6_io_out ? io_r_235_b : _GEN_4824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4826 = 10'hec == r_count_6_io_out ? io_r_236_b : _GEN_4825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4827 = 10'hed == r_count_6_io_out ? io_r_237_b : _GEN_4826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4828 = 10'hee == r_count_6_io_out ? io_r_238_b : _GEN_4827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4829 = 10'hef == r_count_6_io_out ? io_r_239_b : _GEN_4828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4830 = 10'hf0 == r_count_6_io_out ? io_r_240_b : _GEN_4829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4831 = 10'hf1 == r_count_6_io_out ? io_r_241_b : _GEN_4830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4832 = 10'hf2 == r_count_6_io_out ? io_r_242_b : _GEN_4831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4833 = 10'hf3 == r_count_6_io_out ? io_r_243_b : _GEN_4832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4834 = 10'hf4 == r_count_6_io_out ? io_r_244_b : _GEN_4833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4835 = 10'hf5 == r_count_6_io_out ? io_r_245_b : _GEN_4834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4836 = 10'hf6 == r_count_6_io_out ? io_r_246_b : _GEN_4835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4837 = 10'hf7 == r_count_6_io_out ? io_r_247_b : _GEN_4836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4838 = 10'hf8 == r_count_6_io_out ? io_r_248_b : _GEN_4837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4839 = 10'hf9 == r_count_6_io_out ? io_r_249_b : _GEN_4838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4840 = 10'hfa == r_count_6_io_out ? io_r_250_b : _GEN_4839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4841 = 10'hfb == r_count_6_io_out ? io_r_251_b : _GEN_4840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4842 = 10'hfc == r_count_6_io_out ? io_r_252_b : _GEN_4841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4843 = 10'hfd == r_count_6_io_out ? io_r_253_b : _GEN_4842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4844 = 10'hfe == r_count_6_io_out ? io_r_254_b : _GEN_4843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4845 = 10'hff == r_count_6_io_out ? io_r_255_b : _GEN_4844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4846 = 10'h100 == r_count_6_io_out ? io_r_256_b : _GEN_4845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4847 = 10'h101 == r_count_6_io_out ? io_r_257_b : _GEN_4846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4848 = 10'h102 == r_count_6_io_out ? io_r_258_b : _GEN_4847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4849 = 10'h103 == r_count_6_io_out ? io_r_259_b : _GEN_4848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4850 = 10'h104 == r_count_6_io_out ? io_r_260_b : _GEN_4849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4851 = 10'h105 == r_count_6_io_out ? io_r_261_b : _GEN_4850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4852 = 10'h106 == r_count_6_io_out ? io_r_262_b : _GEN_4851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4853 = 10'h107 == r_count_6_io_out ? io_r_263_b : _GEN_4852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4854 = 10'h108 == r_count_6_io_out ? io_r_264_b : _GEN_4853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4855 = 10'h109 == r_count_6_io_out ? io_r_265_b : _GEN_4854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4856 = 10'h10a == r_count_6_io_out ? io_r_266_b : _GEN_4855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4857 = 10'h10b == r_count_6_io_out ? io_r_267_b : _GEN_4856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4858 = 10'h10c == r_count_6_io_out ? io_r_268_b : _GEN_4857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4859 = 10'h10d == r_count_6_io_out ? io_r_269_b : _GEN_4858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4860 = 10'h10e == r_count_6_io_out ? io_r_270_b : _GEN_4859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4861 = 10'h10f == r_count_6_io_out ? io_r_271_b : _GEN_4860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4862 = 10'h110 == r_count_6_io_out ? io_r_272_b : _GEN_4861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4863 = 10'h111 == r_count_6_io_out ? io_r_273_b : _GEN_4862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4864 = 10'h112 == r_count_6_io_out ? io_r_274_b : _GEN_4863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4865 = 10'h113 == r_count_6_io_out ? io_r_275_b : _GEN_4864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4866 = 10'h114 == r_count_6_io_out ? io_r_276_b : _GEN_4865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4867 = 10'h115 == r_count_6_io_out ? io_r_277_b : _GEN_4866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4868 = 10'h116 == r_count_6_io_out ? io_r_278_b : _GEN_4867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4869 = 10'h117 == r_count_6_io_out ? io_r_279_b : _GEN_4868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4870 = 10'h118 == r_count_6_io_out ? io_r_280_b : _GEN_4869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4871 = 10'h119 == r_count_6_io_out ? io_r_281_b : _GEN_4870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4872 = 10'h11a == r_count_6_io_out ? io_r_282_b : _GEN_4871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4873 = 10'h11b == r_count_6_io_out ? io_r_283_b : _GEN_4872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4874 = 10'h11c == r_count_6_io_out ? io_r_284_b : _GEN_4873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4875 = 10'h11d == r_count_6_io_out ? io_r_285_b : _GEN_4874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4876 = 10'h11e == r_count_6_io_out ? io_r_286_b : _GEN_4875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4877 = 10'h11f == r_count_6_io_out ? io_r_287_b : _GEN_4876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4878 = 10'h120 == r_count_6_io_out ? io_r_288_b : _GEN_4877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4879 = 10'h121 == r_count_6_io_out ? io_r_289_b : _GEN_4878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4880 = 10'h122 == r_count_6_io_out ? io_r_290_b : _GEN_4879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4881 = 10'h123 == r_count_6_io_out ? io_r_291_b : _GEN_4880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4882 = 10'h124 == r_count_6_io_out ? io_r_292_b : _GEN_4881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4883 = 10'h125 == r_count_6_io_out ? io_r_293_b : _GEN_4882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4884 = 10'h126 == r_count_6_io_out ? io_r_294_b : _GEN_4883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4885 = 10'h127 == r_count_6_io_out ? io_r_295_b : _GEN_4884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4886 = 10'h128 == r_count_6_io_out ? io_r_296_b : _GEN_4885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4887 = 10'h129 == r_count_6_io_out ? io_r_297_b : _GEN_4886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4888 = 10'h12a == r_count_6_io_out ? io_r_298_b : _GEN_4887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4889 = 10'h12b == r_count_6_io_out ? io_r_299_b : _GEN_4888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4890 = 10'h12c == r_count_6_io_out ? io_r_300_b : _GEN_4889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4891 = 10'h12d == r_count_6_io_out ? io_r_301_b : _GEN_4890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4892 = 10'h12e == r_count_6_io_out ? io_r_302_b : _GEN_4891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4893 = 10'h12f == r_count_6_io_out ? io_r_303_b : _GEN_4892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4894 = 10'h130 == r_count_6_io_out ? io_r_304_b : _GEN_4893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4895 = 10'h131 == r_count_6_io_out ? io_r_305_b : _GEN_4894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4896 = 10'h132 == r_count_6_io_out ? io_r_306_b : _GEN_4895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4897 = 10'h133 == r_count_6_io_out ? io_r_307_b : _GEN_4896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4898 = 10'h134 == r_count_6_io_out ? io_r_308_b : _GEN_4897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4899 = 10'h135 == r_count_6_io_out ? io_r_309_b : _GEN_4898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4900 = 10'h136 == r_count_6_io_out ? io_r_310_b : _GEN_4899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4901 = 10'h137 == r_count_6_io_out ? io_r_311_b : _GEN_4900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4902 = 10'h138 == r_count_6_io_out ? io_r_312_b : _GEN_4901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4903 = 10'h139 == r_count_6_io_out ? io_r_313_b : _GEN_4902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4904 = 10'h13a == r_count_6_io_out ? io_r_314_b : _GEN_4903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4905 = 10'h13b == r_count_6_io_out ? io_r_315_b : _GEN_4904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4906 = 10'h13c == r_count_6_io_out ? io_r_316_b : _GEN_4905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4907 = 10'h13d == r_count_6_io_out ? io_r_317_b : _GEN_4906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4908 = 10'h13e == r_count_6_io_out ? io_r_318_b : _GEN_4907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4909 = 10'h13f == r_count_6_io_out ? io_r_319_b : _GEN_4908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4910 = 10'h140 == r_count_6_io_out ? io_r_320_b : _GEN_4909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4911 = 10'h141 == r_count_6_io_out ? io_r_321_b : _GEN_4910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4912 = 10'h142 == r_count_6_io_out ? io_r_322_b : _GEN_4911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4913 = 10'h143 == r_count_6_io_out ? io_r_323_b : _GEN_4912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4914 = 10'h144 == r_count_6_io_out ? io_r_324_b : _GEN_4913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4915 = 10'h145 == r_count_6_io_out ? io_r_325_b : _GEN_4914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4916 = 10'h146 == r_count_6_io_out ? io_r_326_b : _GEN_4915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4917 = 10'h147 == r_count_6_io_out ? io_r_327_b : _GEN_4916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4918 = 10'h148 == r_count_6_io_out ? io_r_328_b : _GEN_4917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4919 = 10'h149 == r_count_6_io_out ? io_r_329_b : _GEN_4918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4920 = 10'h14a == r_count_6_io_out ? io_r_330_b : _GEN_4919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4921 = 10'h14b == r_count_6_io_out ? io_r_331_b : _GEN_4920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4922 = 10'h14c == r_count_6_io_out ? io_r_332_b : _GEN_4921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4923 = 10'h14d == r_count_6_io_out ? io_r_333_b : _GEN_4922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4924 = 10'h14e == r_count_6_io_out ? io_r_334_b : _GEN_4923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4925 = 10'h14f == r_count_6_io_out ? io_r_335_b : _GEN_4924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4926 = 10'h150 == r_count_6_io_out ? io_r_336_b : _GEN_4925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4927 = 10'h151 == r_count_6_io_out ? io_r_337_b : _GEN_4926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4928 = 10'h152 == r_count_6_io_out ? io_r_338_b : _GEN_4927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4929 = 10'h153 == r_count_6_io_out ? io_r_339_b : _GEN_4928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4930 = 10'h154 == r_count_6_io_out ? io_r_340_b : _GEN_4929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4931 = 10'h155 == r_count_6_io_out ? io_r_341_b : _GEN_4930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4932 = 10'h156 == r_count_6_io_out ? io_r_342_b : _GEN_4931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4933 = 10'h157 == r_count_6_io_out ? io_r_343_b : _GEN_4932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4934 = 10'h158 == r_count_6_io_out ? io_r_344_b : _GEN_4933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4935 = 10'h159 == r_count_6_io_out ? io_r_345_b : _GEN_4934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4936 = 10'h15a == r_count_6_io_out ? io_r_346_b : _GEN_4935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4937 = 10'h15b == r_count_6_io_out ? io_r_347_b : _GEN_4936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4938 = 10'h15c == r_count_6_io_out ? io_r_348_b : _GEN_4937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4939 = 10'h15d == r_count_6_io_out ? io_r_349_b : _GEN_4938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4940 = 10'h15e == r_count_6_io_out ? io_r_350_b : _GEN_4939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4941 = 10'h15f == r_count_6_io_out ? io_r_351_b : _GEN_4940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4942 = 10'h160 == r_count_6_io_out ? io_r_352_b : _GEN_4941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4943 = 10'h161 == r_count_6_io_out ? io_r_353_b : _GEN_4942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4944 = 10'h162 == r_count_6_io_out ? io_r_354_b : _GEN_4943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4945 = 10'h163 == r_count_6_io_out ? io_r_355_b : _GEN_4944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4946 = 10'h164 == r_count_6_io_out ? io_r_356_b : _GEN_4945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4947 = 10'h165 == r_count_6_io_out ? io_r_357_b : _GEN_4946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4948 = 10'h166 == r_count_6_io_out ? io_r_358_b : _GEN_4947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4949 = 10'h167 == r_count_6_io_out ? io_r_359_b : _GEN_4948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4950 = 10'h168 == r_count_6_io_out ? io_r_360_b : _GEN_4949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4951 = 10'h169 == r_count_6_io_out ? io_r_361_b : _GEN_4950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4952 = 10'h16a == r_count_6_io_out ? io_r_362_b : _GEN_4951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4953 = 10'h16b == r_count_6_io_out ? io_r_363_b : _GEN_4952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4954 = 10'h16c == r_count_6_io_out ? io_r_364_b : _GEN_4953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4955 = 10'h16d == r_count_6_io_out ? io_r_365_b : _GEN_4954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4956 = 10'h16e == r_count_6_io_out ? io_r_366_b : _GEN_4955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4957 = 10'h16f == r_count_6_io_out ? io_r_367_b : _GEN_4956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4958 = 10'h170 == r_count_6_io_out ? io_r_368_b : _GEN_4957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4959 = 10'h171 == r_count_6_io_out ? io_r_369_b : _GEN_4958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4960 = 10'h172 == r_count_6_io_out ? io_r_370_b : _GEN_4959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4961 = 10'h173 == r_count_6_io_out ? io_r_371_b : _GEN_4960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4962 = 10'h174 == r_count_6_io_out ? io_r_372_b : _GEN_4961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4963 = 10'h175 == r_count_6_io_out ? io_r_373_b : _GEN_4962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4964 = 10'h176 == r_count_6_io_out ? io_r_374_b : _GEN_4963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4965 = 10'h177 == r_count_6_io_out ? io_r_375_b : _GEN_4964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4966 = 10'h178 == r_count_6_io_out ? io_r_376_b : _GEN_4965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4967 = 10'h179 == r_count_6_io_out ? io_r_377_b : _GEN_4966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4968 = 10'h17a == r_count_6_io_out ? io_r_378_b : _GEN_4967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4969 = 10'h17b == r_count_6_io_out ? io_r_379_b : _GEN_4968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4970 = 10'h17c == r_count_6_io_out ? io_r_380_b : _GEN_4969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4971 = 10'h17d == r_count_6_io_out ? io_r_381_b : _GEN_4970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4972 = 10'h17e == r_count_6_io_out ? io_r_382_b : _GEN_4971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4973 = 10'h17f == r_count_6_io_out ? io_r_383_b : _GEN_4972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4974 = 10'h180 == r_count_6_io_out ? io_r_384_b : _GEN_4973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4975 = 10'h181 == r_count_6_io_out ? io_r_385_b : _GEN_4974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4976 = 10'h182 == r_count_6_io_out ? io_r_386_b : _GEN_4975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4977 = 10'h183 == r_count_6_io_out ? io_r_387_b : _GEN_4976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4978 = 10'h184 == r_count_6_io_out ? io_r_388_b : _GEN_4977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4979 = 10'h185 == r_count_6_io_out ? io_r_389_b : _GEN_4978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4980 = 10'h186 == r_count_6_io_out ? io_r_390_b : _GEN_4979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4981 = 10'h187 == r_count_6_io_out ? io_r_391_b : _GEN_4980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4982 = 10'h188 == r_count_6_io_out ? io_r_392_b : _GEN_4981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4983 = 10'h189 == r_count_6_io_out ? io_r_393_b : _GEN_4982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4984 = 10'h18a == r_count_6_io_out ? io_r_394_b : _GEN_4983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4985 = 10'h18b == r_count_6_io_out ? io_r_395_b : _GEN_4984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4986 = 10'h18c == r_count_6_io_out ? io_r_396_b : _GEN_4985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4987 = 10'h18d == r_count_6_io_out ? io_r_397_b : _GEN_4986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4988 = 10'h18e == r_count_6_io_out ? io_r_398_b : _GEN_4987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4989 = 10'h18f == r_count_6_io_out ? io_r_399_b : _GEN_4988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4990 = 10'h190 == r_count_6_io_out ? io_r_400_b : _GEN_4989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4991 = 10'h191 == r_count_6_io_out ? io_r_401_b : _GEN_4990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4992 = 10'h192 == r_count_6_io_out ? io_r_402_b : _GEN_4991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4993 = 10'h193 == r_count_6_io_out ? io_r_403_b : _GEN_4992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4994 = 10'h194 == r_count_6_io_out ? io_r_404_b : _GEN_4993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4995 = 10'h195 == r_count_6_io_out ? io_r_405_b : _GEN_4994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4996 = 10'h196 == r_count_6_io_out ? io_r_406_b : _GEN_4995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4997 = 10'h197 == r_count_6_io_out ? io_r_407_b : _GEN_4996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4998 = 10'h198 == r_count_6_io_out ? io_r_408_b : _GEN_4997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4999 = 10'h199 == r_count_6_io_out ? io_r_409_b : _GEN_4998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5000 = 10'h19a == r_count_6_io_out ? io_r_410_b : _GEN_4999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5001 = 10'h19b == r_count_6_io_out ? io_r_411_b : _GEN_5000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5002 = 10'h19c == r_count_6_io_out ? io_r_412_b : _GEN_5001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5003 = 10'h19d == r_count_6_io_out ? io_r_413_b : _GEN_5002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5004 = 10'h19e == r_count_6_io_out ? io_r_414_b : _GEN_5003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5005 = 10'h19f == r_count_6_io_out ? io_r_415_b : _GEN_5004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5006 = 10'h1a0 == r_count_6_io_out ? io_r_416_b : _GEN_5005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5007 = 10'h1a1 == r_count_6_io_out ? io_r_417_b : _GEN_5006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5008 = 10'h1a2 == r_count_6_io_out ? io_r_418_b : _GEN_5007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5009 = 10'h1a3 == r_count_6_io_out ? io_r_419_b : _GEN_5008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5010 = 10'h1a4 == r_count_6_io_out ? io_r_420_b : _GEN_5009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5011 = 10'h1a5 == r_count_6_io_out ? io_r_421_b : _GEN_5010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5012 = 10'h1a6 == r_count_6_io_out ? io_r_422_b : _GEN_5011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5013 = 10'h1a7 == r_count_6_io_out ? io_r_423_b : _GEN_5012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5014 = 10'h1a8 == r_count_6_io_out ? io_r_424_b : _GEN_5013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5015 = 10'h1a9 == r_count_6_io_out ? io_r_425_b : _GEN_5014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5016 = 10'h1aa == r_count_6_io_out ? io_r_426_b : _GEN_5015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5017 = 10'h1ab == r_count_6_io_out ? io_r_427_b : _GEN_5016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5018 = 10'h1ac == r_count_6_io_out ? io_r_428_b : _GEN_5017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5019 = 10'h1ad == r_count_6_io_out ? io_r_429_b : _GEN_5018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5020 = 10'h1ae == r_count_6_io_out ? io_r_430_b : _GEN_5019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5021 = 10'h1af == r_count_6_io_out ? io_r_431_b : _GEN_5020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5022 = 10'h1b0 == r_count_6_io_out ? io_r_432_b : _GEN_5021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5023 = 10'h1b1 == r_count_6_io_out ? io_r_433_b : _GEN_5022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5024 = 10'h1b2 == r_count_6_io_out ? io_r_434_b : _GEN_5023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5025 = 10'h1b3 == r_count_6_io_out ? io_r_435_b : _GEN_5024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5026 = 10'h1b4 == r_count_6_io_out ? io_r_436_b : _GEN_5025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5027 = 10'h1b5 == r_count_6_io_out ? io_r_437_b : _GEN_5026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5028 = 10'h1b6 == r_count_6_io_out ? io_r_438_b : _GEN_5027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5029 = 10'h1b7 == r_count_6_io_out ? io_r_439_b : _GEN_5028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5030 = 10'h1b8 == r_count_6_io_out ? io_r_440_b : _GEN_5029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5031 = 10'h1b9 == r_count_6_io_out ? io_r_441_b : _GEN_5030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5032 = 10'h1ba == r_count_6_io_out ? io_r_442_b : _GEN_5031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5033 = 10'h1bb == r_count_6_io_out ? io_r_443_b : _GEN_5032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5034 = 10'h1bc == r_count_6_io_out ? io_r_444_b : _GEN_5033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5035 = 10'h1bd == r_count_6_io_out ? io_r_445_b : _GEN_5034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5036 = 10'h1be == r_count_6_io_out ? io_r_446_b : _GEN_5035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5037 = 10'h1bf == r_count_6_io_out ? io_r_447_b : _GEN_5036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5038 = 10'h1c0 == r_count_6_io_out ? io_r_448_b : _GEN_5037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5039 = 10'h1c1 == r_count_6_io_out ? io_r_449_b : _GEN_5038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5040 = 10'h1c2 == r_count_6_io_out ? io_r_450_b : _GEN_5039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5041 = 10'h1c3 == r_count_6_io_out ? io_r_451_b : _GEN_5040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5042 = 10'h1c4 == r_count_6_io_out ? io_r_452_b : _GEN_5041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5043 = 10'h1c5 == r_count_6_io_out ? io_r_453_b : _GEN_5042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5044 = 10'h1c6 == r_count_6_io_out ? io_r_454_b : _GEN_5043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5045 = 10'h1c7 == r_count_6_io_out ? io_r_455_b : _GEN_5044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5046 = 10'h1c8 == r_count_6_io_out ? io_r_456_b : _GEN_5045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5047 = 10'h1c9 == r_count_6_io_out ? io_r_457_b : _GEN_5046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5048 = 10'h1ca == r_count_6_io_out ? io_r_458_b : _GEN_5047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5049 = 10'h1cb == r_count_6_io_out ? io_r_459_b : _GEN_5048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5050 = 10'h1cc == r_count_6_io_out ? io_r_460_b : _GEN_5049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5051 = 10'h1cd == r_count_6_io_out ? io_r_461_b : _GEN_5050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5052 = 10'h1ce == r_count_6_io_out ? io_r_462_b : _GEN_5051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5053 = 10'h1cf == r_count_6_io_out ? io_r_463_b : _GEN_5052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5054 = 10'h1d0 == r_count_6_io_out ? io_r_464_b : _GEN_5053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5055 = 10'h1d1 == r_count_6_io_out ? io_r_465_b : _GEN_5054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5056 = 10'h1d2 == r_count_6_io_out ? io_r_466_b : _GEN_5055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5057 = 10'h1d3 == r_count_6_io_out ? io_r_467_b : _GEN_5056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5058 = 10'h1d4 == r_count_6_io_out ? io_r_468_b : _GEN_5057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5059 = 10'h1d5 == r_count_6_io_out ? io_r_469_b : _GEN_5058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5060 = 10'h1d6 == r_count_6_io_out ? io_r_470_b : _GEN_5059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5061 = 10'h1d7 == r_count_6_io_out ? io_r_471_b : _GEN_5060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5062 = 10'h1d8 == r_count_6_io_out ? io_r_472_b : _GEN_5061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5063 = 10'h1d9 == r_count_6_io_out ? io_r_473_b : _GEN_5062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5064 = 10'h1da == r_count_6_io_out ? io_r_474_b : _GEN_5063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5065 = 10'h1db == r_count_6_io_out ? io_r_475_b : _GEN_5064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5066 = 10'h1dc == r_count_6_io_out ? io_r_476_b : _GEN_5065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5067 = 10'h1dd == r_count_6_io_out ? io_r_477_b : _GEN_5066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5068 = 10'h1de == r_count_6_io_out ? io_r_478_b : _GEN_5067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5069 = 10'h1df == r_count_6_io_out ? io_r_479_b : _GEN_5068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5070 = 10'h1e0 == r_count_6_io_out ? io_r_480_b : _GEN_5069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5071 = 10'h1e1 == r_count_6_io_out ? io_r_481_b : _GEN_5070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5072 = 10'h1e2 == r_count_6_io_out ? io_r_482_b : _GEN_5071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5073 = 10'h1e3 == r_count_6_io_out ? io_r_483_b : _GEN_5072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5074 = 10'h1e4 == r_count_6_io_out ? io_r_484_b : _GEN_5073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5075 = 10'h1e5 == r_count_6_io_out ? io_r_485_b : _GEN_5074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5076 = 10'h1e6 == r_count_6_io_out ? io_r_486_b : _GEN_5075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5077 = 10'h1e7 == r_count_6_io_out ? io_r_487_b : _GEN_5076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5078 = 10'h1e8 == r_count_6_io_out ? io_r_488_b : _GEN_5077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5079 = 10'h1e9 == r_count_6_io_out ? io_r_489_b : _GEN_5078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5080 = 10'h1ea == r_count_6_io_out ? io_r_490_b : _GEN_5079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5081 = 10'h1eb == r_count_6_io_out ? io_r_491_b : _GEN_5080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5082 = 10'h1ec == r_count_6_io_out ? io_r_492_b : _GEN_5081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5083 = 10'h1ed == r_count_6_io_out ? io_r_493_b : _GEN_5082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5084 = 10'h1ee == r_count_6_io_out ? io_r_494_b : _GEN_5083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5085 = 10'h1ef == r_count_6_io_out ? io_r_495_b : _GEN_5084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5086 = 10'h1f0 == r_count_6_io_out ? io_r_496_b : _GEN_5085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5087 = 10'h1f1 == r_count_6_io_out ? io_r_497_b : _GEN_5086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5088 = 10'h1f2 == r_count_6_io_out ? io_r_498_b : _GEN_5087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5089 = 10'h1f3 == r_count_6_io_out ? io_r_499_b : _GEN_5088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5090 = 10'h1f4 == r_count_6_io_out ? io_r_500_b : _GEN_5089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5091 = 10'h1f5 == r_count_6_io_out ? io_r_501_b : _GEN_5090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5092 = 10'h1f6 == r_count_6_io_out ? io_r_502_b : _GEN_5091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5093 = 10'h1f7 == r_count_6_io_out ? io_r_503_b : _GEN_5092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5094 = 10'h1f8 == r_count_6_io_out ? io_r_504_b : _GEN_5093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5095 = 10'h1f9 == r_count_6_io_out ? io_r_505_b : _GEN_5094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5096 = 10'h1fa == r_count_6_io_out ? io_r_506_b : _GEN_5095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5097 = 10'h1fb == r_count_6_io_out ? io_r_507_b : _GEN_5096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5098 = 10'h1fc == r_count_6_io_out ? io_r_508_b : _GEN_5097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5099 = 10'h1fd == r_count_6_io_out ? io_r_509_b : _GEN_5098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5100 = 10'h1fe == r_count_6_io_out ? io_r_510_b : _GEN_5099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5101 = 10'h1ff == r_count_6_io_out ? io_r_511_b : _GEN_5100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5102 = 10'h200 == r_count_6_io_out ? io_r_512_b : _GEN_5101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5103 = 10'h201 == r_count_6_io_out ? io_r_513_b : _GEN_5102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5104 = 10'h202 == r_count_6_io_out ? io_r_514_b : _GEN_5103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5105 = 10'h203 == r_count_6_io_out ? io_r_515_b : _GEN_5104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5106 = 10'h204 == r_count_6_io_out ? io_r_516_b : _GEN_5105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5107 = 10'h205 == r_count_6_io_out ? io_r_517_b : _GEN_5106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5108 = 10'h206 == r_count_6_io_out ? io_r_518_b : _GEN_5107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5109 = 10'h207 == r_count_6_io_out ? io_r_519_b : _GEN_5108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5110 = 10'h208 == r_count_6_io_out ? io_r_520_b : _GEN_5109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5111 = 10'h209 == r_count_6_io_out ? io_r_521_b : _GEN_5110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5112 = 10'h20a == r_count_6_io_out ? io_r_522_b : _GEN_5111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5113 = 10'h20b == r_count_6_io_out ? io_r_523_b : _GEN_5112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5114 = 10'h20c == r_count_6_io_out ? io_r_524_b : _GEN_5113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5115 = 10'h20d == r_count_6_io_out ? io_r_525_b : _GEN_5114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5116 = 10'h20e == r_count_6_io_out ? io_r_526_b : _GEN_5115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5117 = 10'h20f == r_count_6_io_out ? io_r_527_b : _GEN_5116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5118 = 10'h210 == r_count_6_io_out ? io_r_528_b : _GEN_5117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5119 = 10'h211 == r_count_6_io_out ? io_r_529_b : _GEN_5118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5120 = 10'h212 == r_count_6_io_out ? io_r_530_b : _GEN_5119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5121 = 10'h213 == r_count_6_io_out ? io_r_531_b : _GEN_5120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5122 = 10'h214 == r_count_6_io_out ? io_r_532_b : _GEN_5121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5123 = 10'h215 == r_count_6_io_out ? io_r_533_b : _GEN_5122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5124 = 10'h216 == r_count_6_io_out ? io_r_534_b : _GEN_5123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5125 = 10'h217 == r_count_6_io_out ? io_r_535_b : _GEN_5124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5126 = 10'h218 == r_count_6_io_out ? io_r_536_b : _GEN_5125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5127 = 10'h219 == r_count_6_io_out ? io_r_537_b : _GEN_5126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5128 = 10'h21a == r_count_6_io_out ? io_r_538_b : _GEN_5127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5129 = 10'h21b == r_count_6_io_out ? io_r_539_b : _GEN_5128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5130 = 10'h21c == r_count_6_io_out ? io_r_540_b : _GEN_5129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5131 = 10'h21d == r_count_6_io_out ? io_r_541_b : _GEN_5130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5132 = 10'h21e == r_count_6_io_out ? io_r_542_b : _GEN_5131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5133 = 10'h21f == r_count_6_io_out ? io_r_543_b : _GEN_5132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5134 = 10'h220 == r_count_6_io_out ? io_r_544_b : _GEN_5133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5135 = 10'h221 == r_count_6_io_out ? io_r_545_b : _GEN_5134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5136 = 10'h222 == r_count_6_io_out ? io_r_546_b : _GEN_5135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5137 = 10'h223 == r_count_6_io_out ? io_r_547_b : _GEN_5136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5138 = 10'h224 == r_count_6_io_out ? io_r_548_b : _GEN_5137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5139 = 10'h225 == r_count_6_io_out ? io_r_549_b : _GEN_5138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5140 = 10'h226 == r_count_6_io_out ? io_r_550_b : _GEN_5139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5141 = 10'h227 == r_count_6_io_out ? io_r_551_b : _GEN_5140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5142 = 10'h228 == r_count_6_io_out ? io_r_552_b : _GEN_5141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5143 = 10'h229 == r_count_6_io_out ? io_r_553_b : _GEN_5142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5144 = 10'h22a == r_count_6_io_out ? io_r_554_b : _GEN_5143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5145 = 10'h22b == r_count_6_io_out ? io_r_555_b : _GEN_5144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5146 = 10'h22c == r_count_6_io_out ? io_r_556_b : _GEN_5145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5147 = 10'h22d == r_count_6_io_out ? io_r_557_b : _GEN_5146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5148 = 10'h22e == r_count_6_io_out ? io_r_558_b : _GEN_5147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5149 = 10'h22f == r_count_6_io_out ? io_r_559_b : _GEN_5148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5150 = 10'h230 == r_count_6_io_out ? io_r_560_b : _GEN_5149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5151 = 10'h231 == r_count_6_io_out ? io_r_561_b : _GEN_5150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5152 = 10'h232 == r_count_6_io_out ? io_r_562_b : _GEN_5151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5153 = 10'h233 == r_count_6_io_out ? io_r_563_b : _GEN_5152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5154 = 10'h234 == r_count_6_io_out ? io_r_564_b : _GEN_5153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5155 = 10'h235 == r_count_6_io_out ? io_r_565_b : _GEN_5154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5156 = 10'h236 == r_count_6_io_out ? io_r_566_b : _GEN_5155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5157 = 10'h237 == r_count_6_io_out ? io_r_567_b : _GEN_5156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5158 = 10'h238 == r_count_6_io_out ? io_r_568_b : _GEN_5157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5159 = 10'h239 == r_count_6_io_out ? io_r_569_b : _GEN_5158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5160 = 10'h23a == r_count_6_io_out ? io_r_570_b : _GEN_5159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5161 = 10'h23b == r_count_6_io_out ? io_r_571_b : _GEN_5160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5162 = 10'h23c == r_count_6_io_out ? io_r_572_b : _GEN_5161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5163 = 10'h23d == r_count_6_io_out ? io_r_573_b : _GEN_5162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5164 = 10'h23e == r_count_6_io_out ? io_r_574_b : _GEN_5163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5165 = 10'h23f == r_count_6_io_out ? io_r_575_b : _GEN_5164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5166 = 10'h240 == r_count_6_io_out ? io_r_576_b : _GEN_5165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5167 = 10'h241 == r_count_6_io_out ? io_r_577_b : _GEN_5166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5168 = 10'h242 == r_count_6_io_out ? io_r_578_b : _GEN_5167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5169 = 10'h243 == r_count_6_io_out ? io_r_579_b : _GEN_5168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5170 = 10'h244 == r_count_6_io_out ? io_r_580_b : _GEN_5169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5171 = 10'h245 == r_count_6_io_out ? io_r_581_b : _GEN_5170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5172 = 10'h246 == r_count_6_io_out ? io_r_582_b : _GEN_5171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5173 = 10'h247 == r_count_6_io_out ? io_r_583_b : _GEN_5172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5174 = 10'h248 == r_count_6_io_out ? io_r_584_b : _GEN_5173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5175 = 10'h249 == r_count_6_io_out ? io_r_585_b : _GEN_5174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5176 = 10'h24a == r_count_6_io_out ? io_r_586_b : _GEN_5175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5177 = 10'h24b == r_count_6_io_out ? io_r_587_b : _GEN_5176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5178 = 10'h24c == r_count_6_io_out ? io_r_588_b : _GEN_5177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5179 = 10'h24d == r_count_6_io_out ? io_r_589_b : _GEN_5178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5180 = 10'h24e == r_count_6_io_out ? io_r_590_b : _GEN_5179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5181 = 10'h24f == r_count_6_io_out ? io_r_591_b : _GEN_5180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5182 = 10'h250 == r_count_6_io_out ? io_r_592_b : _GEN_5181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5183 = 10'h251 == r_count_6_io_out ? io_r_593_b : _GEN_5182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5184 = 10'h252 == r_count_6_io_out ? io_r_594_b : _GEN_5183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5185 = 10'h253 == r_count_6_io_out ? io_r_595_b : _GEN_5184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5186 = 10'h254 == r_count_6_io_out ? io_r_596_b : _GEN_5185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5187 = 10'h255 == r_count_6_io_out ? io_r_597_b : _GEN_5186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5188 = 10'h256 == r_count_6_io_out ? io_r_598_b : _GEN_5187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5189 = 10'h257 == r_count_6_io_out ? io_r_599_b : _GEN_5188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5190 = 10'h258 == r_count_6_io_out ? io_r_600_b : _GEN_5189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5191 = 10'h259 == r_count_6_io_out ? io_r_601_b : _GEN_5190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5192 = 10'h25a == r_count_6_io_out ? io_r_602_b : _GEN_5191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5193 = 10'h25b == r_count_6_io_out ? io_r_603_b : _GEN_5192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5194 = 10'h25c == r_count_6_io_out ? io_r_604_b : _GEN_5193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5195 = 10'h25d == r_count_6_io_out ? io_r_605_b : _GEN_5194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5196 = 10'h25e == r_count_6_io_out ? io_r_606_b : _GEN_5195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5197 = 10'h25f == r_count_6_io_out ? io_r_607_b : _GEN_5196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5198 = 10'h260 == r_count_6_io_out ? io_r_608_b : _GEN_5197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5199 = 10'h261 == r_count_6_io_out ? io_r_609_b : _GEN_5198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5200 = 10'h262 == r_count_6_io_out ? io_r_610_b : _GEN_5199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5201 = 10'h263 == r_count_6_io_out ? io_r_611_b : _GEN_5200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5202 = 10'h264 == r_count_6_io_out ? io_r_612_b : _GEN_5201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5203 = 10'h265 == r_count_6_io_out ? io_r_613_b : _GEN_5202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5204 = 10'h266 == r_count_6_io_out ? io_r_614_b : _GEN_5203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5205 = 10'h267 == r_count_6_io_out ? io_r_615_b : _GEN_5204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5206 = 10'h268 == r_count_6_io_out ? io_r_616_b : _GEN_5205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5207 = 10'h269 == r_count_6_io_out ? io_r_617_b : _GEN_5206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5208 = 10'h26a == r_count_6_io_out ? io_r_618_b : _GEN_5207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5209 = 10'h26b == r_count_6_io_out ? io_r_619_b : _GEN_5208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5210 = 10'h26c == r_count_6_io_out ? io_r_620_b : _GEN_5209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5211 = 10'h26d == r_count_6_io_out ? io_r_621_b : _GEN_5210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5212 = 10'h26e == r_count_6_io_out ? io_r_622_b : _GEN_5211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5213 = 10'h26f == r_count_6_io_out ? io_r_623_b : _GEN_5212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5214 = 10'h270 == r_count_6_io_out ? io_r_624_b : _GEN_5213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5215 = 10'h271 == r_count_6_io_out ? io_r_625_b : _GEN_5214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5216 = 10'h272 == r_count_6_io_out ? io_r_626_b : _GEN_5215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5217 = 10'h273 == r_count_6_io_out ? io_r_627_b : _GEN_5216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5218 = 10'h274 == r_count_6_io_out ? io_r_628_b : _GEN_5217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5219 = 10'h275 == r_count_6_io_out ? io_r_629_b : _GEN_5218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5220 = 10'h276 == r_count_6_io_out ? io_r_630_b : _GEN_5219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5221 = 10'h277 == r_count_6_io_out ? io_r_631_b : _GEN_5220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5222 = 10'h278 == r_count_6_io_out ? io_r_632_b : _GEN_5221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5223 = 10'h279 == r_count_6_io_out ? io_r_633_b : _GEN_5222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5224 = 10'h27a == r_count_6_io_out ? io_r_634_b : _GEN_5223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5225 = 10'h27b == r_count_6_io_out ? io_r_635_b : _GEN_5224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5226 = 10'h27c == r_count_6_io_out ? io_r_636_b : _GEN_5225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5227 = 10'h27d == r_count_6_io_out ? io_r_637_b : _GEN_5226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5228 = 10'h27e == r_count_6_io_out ? io_r_638_b : _GEN_5227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5229 = 10'h27f == r_count_6_io_out ? io_r_639_b : _GEN_5228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5230 = 10'h280 == r_count_6_io_out ? io_r_640_b : _GEN_5229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5231 = 10'h281 == r_count_6_io_out ? io_r_641_b : _GEN_5230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5232 = 10'h282 == r_count_6_io_out ? io_r_642_b : _GEN_5231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5233 = 10'h283 == r_count_6_io_out ? io_r_643_b : _GEN_5232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5234 = 10'h284 == r_count_6_io_out ? io_r_644_b : _GEN_5233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5235 = 10'h285 == r_count_6_io_out ? io_r_645_b : _GEN_5234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5236 = 10'h286 == r_count_6_io_out ? io_r_646_b : _GEN_5235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5237 = 10'h287 == r_count_6_io_out ? io_r_647_b : _GEN_5236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5238 = 10'h288 == r_count_6_io_out ? io_r_648_b : _GEN_5237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5239 = 10'h289 == r_count_6_io_out ? io_r_649_b : _GEN_5238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5240 = 10'h28a == r_count_6_io_out ? io_r_650_b : _GEN_5239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5241 = 10'h28b == r_count_6_io_out ? io_r_651_b : _GEN_5240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5242 = 10'h28c == r_count_6_io_out ? io_r_652_b : _GEN_5241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5243 = 10'h28d == r_count_6_io_out ? io_r_653_b : _GEN_5242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5244 = 10'h28e == r_count_6_io_out ? io_r_654_b : _GEN_5243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5245 = 10'h28f == r_count_6_io_out ? io_r_655_b : _GEN_5244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5246 = 10'h290 == r_count_6_io_out ? io_r_656_b : _GEN_5245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5247 = 10'h291 == r_count_6_io_out ? io_r_657_b : _GEN_5246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5248 = 10'h292 == r_count_6_io_out ? io_r_658_b : _GEN_5247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5249 = 10'h293 == r_count_6_io_out ? io_r_659_b : _GEN_5248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5250 = 10'h294 == r_count_6_io_out ? io_r_660_b : _GEN_5249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5251 = 10'h295 == r_count_6_io_out ? io_r_661_b : _GEN_5250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5252 = 10'h296 == r_count_6_io_out ? io_r_662_b : _GEN_5251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5253 = 10'h297 == r_count_6_io_out ? io_r_663_b : _GEN_5252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5254 = 10'h298 == r_count_6_io_out ? io_r_664_b : _GEN_5253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5255 = 10'h299 == r_count_6_io_out ? io_r_665_b : _GEN_5254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5256 = 10'h29a == r_count_6_io_out ? io_r_666_b : _GEN_5255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5257 = 10'h29b == r_count_6_io_out ? io_r_667_b : _GEN_5256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5258 = 10'h29c == r_count_6_io_out ? io_r_668_b : _GEN_5257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5259 = 10'h29d == r_count_6_io_out ? io_r_669_b : _GEN_5258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5260 = 10'h29e == r_count_6_io_out ? io_r_670_b : _GEN_5259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5261 = 10'h29f == r_count_6_io_out ? io_r_671_b : _GEN_5260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5262 = 10'h2a0 == r_count_6_io_out ? io_r_672_b : _GEN_5261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5263 = 10'h2a1 == r_count_6_io_out ? io_r_673_b : _GEN_5262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5264 = 10'h2a2 == r_count_6_io_out ? io_r_674_b : _GEN_5263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5265 = 10'h2a3 == r_count_6_io_out ? io_r_675_b : _GEN_5264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5266 = 10'h2a4 == r_count_6_io_out ? io_r_676_b : _GEN_5265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5267 = 10'h2a5 == r_count_6_io_out ? io_r_677_b : _GEN_5266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5268 = 10'h2a6 == r_count_6_io_out ? io_r_678_b : _GEN_5267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5269 = 10'h2a7 == r_count_6_io_out ? io_r_679_b : _GEN_5268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5270 = 10'h2a8 == r_count_6_io_out ? io_r_680_b : _GEN_5269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5271 = 10'h2a9 == r_count_6_io_out ? io_r_681_b : _GEN_5270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5272 = 10'h2aa == r_count_6_io_out ? io_r_682_b : _GEN_5271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5273 = 10'h2ab == r_count_6_io_out ? io_r_683_b : _GEN_5272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5274 = 10'h2ac == r_count_6_io_out ? io_r_684_b : _GEN_5273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5275 = 10'h2ad == r_count_6_io_out ? io_r_685_b : _GEN_5274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5276 = 10'h2ae == r_count_6_io_out ? io_r_686_b : _GEN_5275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5277 = 10'h2af == r_count_6_io_out ? io_r_687_b : _GEN_5276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5278 = 10'h2b0 == r_count_6_io_out ? io_r_688_b : _GEN_5277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5279 = 10'h2b1 == r_count_6_io_out ? io_r_689_b : _GEN_5278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5280 = 10'h2b2 == r_count_6_io_out ? io_r_690_b : _GEN_5279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5281 = 10'h2b3 == r_count_6_io_out ? io_r_691_b : _GEN_5280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5282 = 10'h2b4 == r_count_6_io_out ? io_r_692_b : _GEN_5281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5283 = 10'h2b5 == r_count_6_io_out ? io_r_693_b : _GEN_5282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5284 = 10'h2b6 == r_count_6_io_out ? io_r_694_b : _GEN_5283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5285 = 10'h2b7 == r_count_6_io_out ? io_r_695_b : _GEN_5284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5286 = 10'h2b8 == r_count_6_io_out ? io_r_696_b : _GEN_5285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5287 = 10'h2b9 == r_count_6_io_out ? io_r_697_b : _GEN_5286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5288 = 10'h2ba == r_count_6_io_out ? io_r_698_b : _GEN_5287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5289 = 10'h2bb == r_count_6_io_out ? io_r_699_b : _GEN_5288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5290 = 10'h2bc == r_count_6_io_out ? io_r_700_b : _GEN_5289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5291 = 10'h2bd == r_count_6_io_out ? io_r_701_b : _GEN_5290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5292 = 10'h2be == r_count_6_io_out ? io_r_702_b : _GEN_5291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5293 = 10'h2bf == r_count_6_io_out ? io_r_703_b : _GEN_5292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5294 = 10'h2c0 == r_count_6_io_out ? io_r_704_b : _GEN_5293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5295 = 10'h2c1 == r_count_6_io_out ? io_r_705_b : _GEN_5294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5296 = 10'h2c2 == r_count_6_io_out ? io_r_706_b : _GEN_5295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5297 = 10'h2c3 == r_count_6_io_out ? io_r_707_b : _GEN_5296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5298 = 10'h2c4 == r_count_6_io_out ? io_r_708_b : _GEN_5297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5299 = 10'h2c5 == r_count_6_io_out ? io_r_709_b : _GEN_5298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5300 = 10'h2c6 == r_count_6_io_out ? io_r_710_b : _GEN_5299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5301 = 10'h2c7 == r_count_6_io_out ? io_r_711_b : _GEN_5300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5302 = 10'h2c8 == r_count_6_io_out ? io_r_712_b : _GEN_5301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5303 = 10'h2c9 == r_count_6_io_out ? io_r_713_b : _GEN_5302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5304 = 10'h2ca == r_count_6_io_out ? io_r_714_b : _GEN_5303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5305 = 10'h2cb == r_count_6_io_out ? io_r_715_b : _GEN_5304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5306 = 10'h2cc == r_count_6_io_out ? io_r_716_b : _GEN_5305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5307 = 10'h2cd == r_count_6_io_out ? io_r_717_b : _GEN_5306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5308 = 10'h2ce == r_count_6_io_out ? io_r_718_b : _GEN_5307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5309 = 10'h2cf == r_count_6_io_out ? io_r_719_b : _GEN_5308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5310 = 10'h2d0 == r_count_6_io_out ? io_r_720_b : _GEN_5309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5311 = 10'h2d1 == r_count_6_io_out ? io_r_721_b : _GEN_5310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5312 = 10'h2d2 == r_count_6_io_out ? io_r_722_b : _GEN_5311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5313 = 10'h2d3 == r_count_6_io_out ? io_r_723_b : _GEN_5312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5314 = 10'h2d4 == r_count_6_io_out ? io_r_724_b : _GEN_5313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5315 = 10'h2d5 == r_count_6_io_out ? io_r_725_b : _GEN_5314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5316 = 10'h2d6 == r_count_6_io_out ? io_r_726_b : _GEN_5315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5317 = 10'h2d7 == r_count_6_io_out ? io_r_727_b : _GEN_5316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5318 = 10'h2d8 == r_count_6_io_out ? io_r_728_b : _GEN_5317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5319 = 10'h2d9 == r_count_6_io_out ? io_r_729_b : _GEN_5318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5320 = 10'h2da == r_count_6_io_out ? io_r_730_b : _GEN_5319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5321 = 10'h2db == r_count_6_io_out ? io_r_731_b : _GEN_5320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5322 = 10'h2dc == r_count_6_io_out ? io_r_732_b : _GEN_5321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5323 = 10'h2dd == r_count_6_io_out ? io_r_733_b : _GEN_5322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5324 = 10'h2de == r_count_6_io_out ? io_r_734_b : _GEN_5323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5325 = 10'h2df == r_count_6_io_out ? io_r_735_b : _GEN_5324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5326 = 10'h2e0 == r_count_6_io_out ? io_r_736_b : _GEN_5325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5327 = 10'h2e1 == r_count_6_io_out ? io_r_737_b : _GEN_5326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5328 = 10'h2e2 == r_count_6_io_out ? io_r_738_b : _GEN_5327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5329 = 10'h2e3 == r_count_6_io_out ? io_r_739_b : _GEN_5328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5330 = 10'h2e4 == r_count_6_io_out ? io_r_740_b : _GEN_5329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5331 = 10'h2e5 == r_count_6_io_out ? io_r_741_b : _GEN_5330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5332 = 10'h2e6 == r_count_6_io_out ? io_r_742_b : _GEN_5331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5333 = 10'h2e7 == r_count_6_io_out ? io_r_743_b : _GEN_5332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5334 = 10'h2e8 == r_count_6_io_out ? io_r_744_b : _GEN_5333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5335 = 10'h2e9 == r_count_6_io_out ? io_r_745_b : _GEN_5334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5336 = 10'h2ea == r_count_6_io_out ? io_r_746_b : _GEN_5335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5337 = 10'h2eb == r_count_6_io_out ? io_r_747_b : _GEN_5336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5338 = 10'h2ec == r_count_6_io_out ? io_r_748_b : _GEN_5337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5341 = 10'h1 == r_count_7_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5342 = 10'h2 == r_count_7_io_out ? io_r_2_b : _GEN_5341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5343 = 10'h3 == r_count_7_io_out ? io_r_3_b : _GEN_5342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5344 = 10'h4 == r_count_7_io_out ? io_r_4_b : _GEN_5343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5345 = 10'h5 == r_count_7_io_out ? io_r_5_b : _GEN_5344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5346 = 10'h6 == r_count_7_io_out ? io_r_6_b : _GEN_5345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5347 = 10'h7 == r_count_7_io_out ? io_r_7_b : _GEN_5346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5348 = 10'h8 == r_count_7_io_out ? io_r_8_b : _GEN_5347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5349 = 10'h9 == r_count_7_io_out ? io_r_9_b : _GEN_5348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5350 = 10'ha == r_count_7_io_out ? io_r_10_b : _GEN_5349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5351 = 10'hb == r_count_7_io_out ? io_r_11_b : _GEN_5350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5352 = 10'hc == r_count_7_io_out ? io_r_12_b : _GEN_5351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5353 = 10'hd == r_count_7_io_out ? io_r_13_b : _GEN_5352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5354 = 10'he == r_count_7_io_out ? io_r_14_b : _GEN_5353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5355 = 10'hf == r_count_7_io_out ? io_r_15_b : _GEN_5354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5356 = 10'h10 == r_count_7_io_out ? io_r_16_b : _GEN_5355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5357 = 10'h11 == r_count_7_io_out ? io_r_17_b : _GEN_5356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5358 = 10'h12 == r_count_7_io_out ? io_r_18_b : _GEN_5357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5359 = 10'h13 == r_count_7_io_out ? io_r_19_b : _GEN_5358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5360 = 10'h14 == r_count_7_io_out ? io_r_20_b : _GEN_5359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5361 = 10'h15 == r_count_7_io_out ? io_r_21_b : _GEN_5360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5362 = 10'h16 == r_count_7_io_out ? io_r_22_b : _GEN_5361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5363 = 10'h17 == r_count_7_io_out ? io_r_23_b : _GEN_5362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5364 = 10'h18 == r_count_7_io_out ? io_r_24_b : _GEN_5363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5365 = 10'h19 == r_count_7_io_out ? io_r_25_b : _GEN_5364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5366 = 10'h1a == r_count_7_io_out ? io_r_26_b : _GEN_5365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5367 = 10'h1b == r_count_7_io_out ? io_r_27_b : _GEN_5366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5368 = 10'h1c == r_count_7_io_out ? io_r_28_b : _GEN_5367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5369 = 10'h1d == r_count_7_io_out ? io_r_29_b : _GEN_5368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5370 = 10'h1e == r_count_7_io_out ? io_r_30_b : _GEN_5369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5371 = 10'h1f == r_count_7_io_out ? io_r_31_b : _GEN_5370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5372 = 10'h20 == r_count_7_io_out ? io_r_32_b : _GEN_5371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5373 = 10'h21 == r_count_7_io_out ? io_r_33_b : _GEN_5372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5374 = 10'h22 == r_count_7_io_out ? io_r_34_b : _GEN_5373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5375 = 10'h23 == r_count_7_io_out ? io_r_35_b : _GEN_5374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5376 = 10'h24 == r_count_7_io_out ? io_r_36_b : _GEN_5375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5377 = 10'h25 == r_count_7_io_out ? io_r_37_b : _GEN_5376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5378 = 10'h26 == r_count_7_io_out ? io_r_38_b : _GEN_5377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5379 = 10'h27 == r_count_7_io_out ? io_r_39_b : _GEN_5378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5380 = 10'h28 == r_count_7_io_out ? io_r_40_b : _GEN_5379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5381 = 10'h29 == r_count_7_io_out ? io_r_41_b : _GEN_5380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5382 = 10'h2a == r_count_7_io_out ? io_r_42_b : _GEN_5381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5383 = 10'h2b == r_count_7_io_out ? io_r_43_b : _GEN_5382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5384 = 10'h2c == r_count_7_io_out ? io_r_44_b : _GEN_5383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5385 = 10'h2d == r_count_7_io_out ? io_r_45_b : _GEN_5384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5386 = 10'h2e == r_count_7_io_out ? io_r_46_b : _GEN_5385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5387 = 10'h2f == r_count_7_io_out ? io_r_47_b : _GEN_5386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5388 = 10'h30 == r_count_7_io_out ? io_r_48_b : _GEN_5387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5389 = 10'h31 == r_count_7_io_out ? io_r_49_b : _GEN_5388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5390 = 10'h32 == r_count_7_io_out ? io_r_50_b : _GEN_5389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5391 = 10'h33 == r_count_7_io_out ? io_r_51_b : _GEN_5390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5392 = 10'h34 == r_count_7_io_out ? io_r_52_b : _GEN_5391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5393 = 10'h35 == r_count_7_io_out ? io_r_53_b : _GEN_5392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5394 = 10'h36 == r_count_7_io_out ? io_r_54_b : _GEN_5393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5395 = 10'h37 == r_count_7_io_out ? io_r_55_b : _GEN_5394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5396 = 10'h38 == r_count_7_io_out ? io_r_56_b : _GEN_5395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5397 = 10'h39 == r_count_7_io_out ? io_r_57_b : _GEN_5396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5398 = 10'h3a == r_count_7_io_out ? io_r_58_b : _GEN_5397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5399 = 10'h3b == r_count_7_io_out ? io_r_59_b : _GEN_5398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5400 = 10'h3c == r_count_7_io_out ? io_r_60_b : _GEN_5399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5401 = 10'h3d == r_count_7_io_out ? io_r_61_b : _GEN_5400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5402 = 10'h3e == r_count_7_io_out ? io_r_62_b : _GEN_5401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5403 = 10'h3f == r_count_7_io_out ? io_r_63_b : _GEN_5402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5404 = 10'h40 == r_count_7_io_out ? io_r_64_b : _GEN_5403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5405 = 10'h41 == r_count_7_io_out ? io_r_65_b : _GEN_5404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5406 = 10'h42 == r_count_7_io_out ? io_r_66_b : _GEN_5405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5407 = 10'h43 == r_count_7_io_out ? io_r_67_b : _GEN_5406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5408 = 10'h44 == r_count_7_io_out ? io_r_68_b : _GEN_5407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5409 = 10'h45 == r_count_7_io_out ? io_r_69_b : _GEN_5408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5410 = 10'h46 == r_count_7_io_out ? io_r_70_b : _GEN_5409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5411 = 10'h47 == r_count_7_io_out ? io_r_71_b : _GEN_5410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5412 = 10'h48 == r_count_7_io_out ? io_r_72_b : _GEN_5411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5413 = 10'h49 == r_count_7_io_out ? io_r_73_b : _GEN_5412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5414 = 10'h4a == r_count_7_io_out ? io_r_74_b : _GEN_5413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5415 = 10'h4b == r_count_7_io_out ? io_r_75_b : _GEN_5414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5416 = 10'h4c == r_count_7_io_out ? io_r_76_b : _GEN_5415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5417 = 10'h4d == r_count_7_io_out ? io_r_77_b : _GEN_5416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5418 = 10'h4e == r_count_7_io_out ? io_r_78_b : _GEN_5417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5419 = 10'h4f == r_count_7_io_out ? io_r_79_b : _GEN_5418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5420 = 10'h50 == r_count_7_io_out ? io_r_80_b : _GEN_5419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5421 = 10'h51 == r_count_7_io_out ? io_r_81_b : _GEN_5420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5422 = 10'h52 == r_count_7_io_out ? io_r_82_b : _GEN_5421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5423 = 10'h53 == r_count_7_io_out ? io_r_83_b : _GEN_5422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5424 = 10'h54 == r_count_7_io_out ? io_r_84_b : _GEN_5423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5425 = 10'h55 == r_count_7_io_out ? io_r_85_b : _GEN_5424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5426 = 10'h56 == r_count_7_io_out ? io_r_86_b : _GEN_5425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5427 = 10'h57 == r_count_7_io_out ? io_r_87_b : _GEN_5426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5428 = 10'h58 == r_count_7_io_out ? io_r_88_b : _GEN_5427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5429 = 10'h59 == r_count_7_io_out ? io_r_89_b : _GEN_5428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5430 = 10'h5a == r_count_7_io_out ? io_r_90_b : _GEN_5429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5431 = 10'h5b == r_count_7_io_out ? io_r_91_b : _GEN_5430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5432 = 10'h5c == r_count_7_io_out ? io_r_92_b : _GEN_5431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5433 = 10'h5d == r_count_7_io_out ? io_r_93_b : _GEN_5432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5434 = 10'h5e == r_count_7_io_out ? io_r_94_b : _GEN_5433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5435 = 10'h5f == r_count_7_io_out ? io_r_95_b : _GEN_5434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5436 = 10'h60 == r_count_7_io_out ? io_r_96_b : _GEN_5435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5437 = 10'h61 == r_count_7_io_out ? io_r_97_b : _GEN_5436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5438 = 10'h62 == r_count_7_io_out ? io_r_98_b : _GEN_5437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5439 = 10'h63 == r_count_7_io_out ? io_r_99_b : _GEN_5438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5440 = 10'h64 == r_count_7_io_out ? io_r_100_b : _GEN_5439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5441 = 10'h65 == r_count_7_io_out ? io_r_101_b : _GEN_5440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5442 = 10'h66 == r_count_7_io_out ? io_r_102_b : _GEN_5441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5443 = 10'h67 == r_count_7_io_out ? io_r_103_b : _GEN_5442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5444 = 10'h68 == r_count_7_io_out ? io_r_104_b : _GEN_5443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5445 = 10'h69 == r_count_7_io_out ? io_r_105_b : _GEN_5444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5446 = 10'h6a == r_count_7_io_out ? io_r_106_b : _GEN_5445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5447 = 10'h6b == r_count_7_io_out ? io_r_107_b : _GEN_5446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5448 = 10'h6c == r_count_7_io_out ? io_r_108_b : _GEN_5447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5449 = 10'h6d == r_count_7_io_out ? io_r_109_b : _GEN_5448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5450 = 10'h6e == r_count_7_io_out ? io_r_110_b : _GEN_5449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5451 = 10'h6f == r_count_7_io_out ? io_r_111_b : _GEN_5450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5452 = 10'h70 == r_count_7_io_out ? io_r_112_b : _GEN_5451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5453 = 10'h71 == r_count_7_io_out ? io_r_113_b : _GEN_5452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5454 = 10'h72 == r_count_7_io_out ? io_r_114_b : _GEN_5453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5455 = 10'h73 == r_count_7_io_out ? io_r_115_b : _GEN_5454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5456 = 10'h74 == r_count_7_io_out ? io_r_116_b : _GEN_5455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5457 = 10'h75 == r_count_7_io_out ? io_r_117_b : _GEN_5456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5458 = 10'h76 == r_count_7_io_out ? io_r_118_b : _GEN_5457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5459 = 10'h77 == r_count_7_io_out ? io_r_119_b : _GEN_5458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5460 = 10'h78 == r_count_7_io_out ? io_r_120_b : _GEN_5459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5461 = 10'h79 == r_count_7_io_out ? io_r_121_b : _GEN_5460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5462 = 10'h7a == r_count_7_io_out ? io_r_122_b : _GEN_5461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5463 = 10'h7b == r_count_7_io_out ? io_r_123_b : _GEN_5462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5464 = 10'h7c == r_count_7_io_out ? io_r_124_b : _GEN_5463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5465 = 10'h7d == r_count_7_io_out ? io_r_125_b : _GEN_5464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5466 = 10'h7e == r_count_7_io_out ? io_r_126_b : _GEN_5465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5467 = 10'h7f == r_count_7_io_out ? io_r_127_b : _GEN_5466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5468 = 10'h80 == r_count_7_io_out ? io_r_128_b : _GEN_5467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5469 = 10'h81 == r_count_7_io_out ? io_r_129_b : _GEN_5468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5470 = 10'h82 == r_count_7_io_out ? io_r_130_b : _GEN_5469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5471 = 10'h83 == r_count_7_io_out ? io_r_131_b : _GEN_5470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5472 = 10'h84 == r_count_7_io_out ? io_r_132_b : _GEN_5471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5473 = 10'h85 == r_count_7_io_out ? io_r_133_b : _GEN_5472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5474 = 10'h86 == r_count_7_io_out ? io_r_134_b : _GEN_5473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5475 = 10'h87 == r_count_7_io_out ? io_r_135_b : _GEN_5474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5476 = 10'h88 == r_count_7_io_out ? io_r_136_b : _GEN_5475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5477 = 10'h89 == r_count_7_io_out ? io_r_137_b : _GEN_5476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5478 = 10'h8a == r_count_7_io_out ? io_r_138_b : _GEN_5477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5479 = 10'h8b == r_count_7_io_out ? io_r_139_b : _GEN_5478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5480 = 10'h8c == r_count_7_io_out ? io_r_140_b : _GEN_5479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5481 = 10'h8d == r_count_7_io_out ? io_r_141_b : _GEN_5480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5482 = 10'h8e == r_count_7_io_out ? io_r_142_b : _GEN_5481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5483 = 10'h8f == r_count_7_io_out ? io_r_143_b : _GEN_5482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5484 = 10'h90 == r_count_7_io_out ? io_r_144_b : _GEN_5483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5485 = 10'h91 == r_count_7_io_out ? io_r_145_b : _GEN_5484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5486 = 10'h92 == r_count_7_io_out ? io_r_146_b : _GEN_5485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5487 = 10'h93 == r_count_7_io_out ? io_r_147_b : _GEN_5486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5488 = 10'h94 == r_count_7_io_out ? io_r_148_b : _GEN_5487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5489 = 10'h95 == r_count_7_io_out ? io_r_149_b : _GEN_5488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5490 = 10'h96 == r_count_7_io_out ? io_r_150_b : _GEN_5489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5491 = 10'h97 == r_count_7_io_out ? io_r_151_b : _GEN_5490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5492 = 10'h98 == r_count_7_io_out ? io_r_152_b : _GEN_5491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5493 = 10'h99 == r_count_7_io_out ? io_r_153_b : _GEN_5492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5494 = 10'h9a == r_count_7_io_out ? io_r_154_b : _GEN_5493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5495 = 10'h9b == r_count_7_io_out ? io_r_155_b : _GEN_5494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5496 = 10'h9c == r_count_7_io_out ? io_r_156_b : _GEN_5495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5497 = 10'h9d == r_count_7_io_out ? io_r_157_b : _GEN_5496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5498 = 10'h9e == r_count_7_io_out ? io_r_158_b : _GEN_5497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5499 = 10'h9f == r_count_7_io_out ? io_r_159_b : _GEN_5498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5500 = 10'ha0 == r_count_7_io_out ? io_r_160_b : _GEN_5499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5501 = 10'ha1 == r_count_7_io_out ? io_r_161_b : _GEN_5500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5502 = 10'ha2 == r_count_7_io_out ? io_r_162_b : _GEN_5501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5503 = 10'ha3 == r_count_7_io_out ? io_r_163_b : _GEN_5502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5504 = 10'ha4 == r_count_7_io_out ? io_r_164_b : _GEN_5503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5505 = 10'ha5 == r_count_7_io_out ? io_r_165_b : _GEN_5504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5506 = 10'ha6 == r_count_7_io_out ? io_r_166_b : _GEN_5505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5507 = 10'ha7 == r_count_7_io_out ? io_r_167_b : _GEN_5506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5508 = 10'ha8 == r_count_7_io_out ? io_r_168_b : _GEN_5507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5509 = 10'ha9 == r_count_7_io_out ? io_r_169_b : _GEN_5508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5510 = 10'haa == r_count_7_io_out ? io_r_170_b : _GEN_5509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5511 = 10'hab == r_count_7_io_out ? io_r_171_b : _GEN_5510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5512 = 10'hac == r_count_7_io_out ? io_r_172_b : _GEN_5511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5513 = 10'had == r_count_7_io_out ? io_r_173_b : _GEN_5512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5514 = 10'hae == r_count_7_io_out ? io_r_174_b : _GEN_5513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5515 = 10'haf == r_count_7_io_out ? io_r_175_b : _GEN_5514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5516 = 10'hb0 == r_count_7_io_out ? io_r_176_b : _GEN_5515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5517 = 10'hb1 == r_count_7_io_out ? io_r_177_b : _GEN_5516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5518 = 10'hb2 == r_count_7_io_out ? io_r_178_b : _GEN_5517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5519 = 10'hb3 == r_count_7_io_out ? io_r_179_b : _GEN_5518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5520 = 10'hb4 == r_count_7_io_out ? io_r_180_b : _GEN_5519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5521 = 10'hb5 == r_count_7_io_out ? io_r_181_b : _GEN_5520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5522 = 10'hb6 == r_count_7_io_out ? io_r_182_b : _GEN_5521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5523 = 10'hb7 == r_count_7_io_out ? io_r_183_b : _GEN_5522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5524 = 10'hb8 == r_count_7_io_out ? io_r_184_b : _GEN_5523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5525 = 10'hb9 == r_count_7_io_out ? io_r_185_b : _GEN_5524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5526 = 10'hba == r_count_7_io_out ? io_r_186_b : _GEN_5525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5527 = 10'hbb == r_count_7_io_out ? io_r_187_b : _GEN_5526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5528 = 10'hbc == r_count_7_io_out ? io_r_188_b : _GEN_5527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5529 = 10'hbd == r_count_7_io_out ? io_r_189_b : _GEN_5528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5530 = 10'hbe == r_count_7_io_out ? io_r_190_b : _GEN_5529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5531 = 10'hbf == r_count_7_io_out ? io_r_191_b : _GEN_5530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5532 = 10'hc0 == r_count_7_io_out ? io_r_192_b : _GEN_5531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5533 = 10'hc1 == r_count_7_io_out ? io_r_193_b : _GEN_5532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5534 = 10'hc2 == r_count_7_io_out ? io_r_194_b : _GEN_5533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5535 = 10'hc3 == r_count_7_io_out ? io_r_195_b : _GEN_5534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5536 = 10'hc4 == r_count_7_io_out ? io_r_196_b : _GEN_5535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5537 = 10'hc5 == r_count_7_io_out ? io_r_197_b : _GEN_5536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5538 = 10'hc6 == r_count_7_io_out ? io_r_198_b : _GEN_5537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5539 = 10'hc7 == r_count_7_io_out ? io_r_199_b : _GEN_5538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5540 = 10'hc8 == r_count_7_io_out ? io_r_200_b : _GEN_5539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5541 = 10'hc9 == r_count_7_io_out ? io_r_201_b : _GEN_5540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5542 = 10'hca == r_count_7_io_out ? io_r_202_b : _GEN_5541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5543 = 10'hcb == r_count_7_io_out ? io_r_203_b : _GEN_5542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5544 = 10'hcc == r_count_7_io_out ? io_r_204_b : _GEN_5543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5545 = 10'hcd == r_count_7_io_out ? io_r_205_b : _GEN_5544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5546 = 10'hce == r_count_7_io_out ? io_r_206_b : _GEN_5545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5547 = 10'hcf == r_count_7_io_out ? io_r_207_b : _GEN_5546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5548 = 10'hd0 == r_count_7_io_out ? io_r_208_b : _GEN_5547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5549 = 10'hd1 == r_count_7_io_out ? io_r_209_b : _GEN_5548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5550 = 10'hd2 == r_count_7_io_out ? io_r_210_b : _GEN_5549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5551 = 10'hd3 == r_count_7_io_out ? io_r_211_b : _GEN_5550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5552 = 10'hd4 == r_count_7_io_out ? io_r_212_b : _GEN_5551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5553 = 10'hd5 == r_count_7_io_out ? io_r_213_b : _GEN_5552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5554 = 10'hd6 == r_count_7_io_out ? io_r_214_b : _GEN_5553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5555 = 10'hd7 == r_count_7_io_out ? io_r_215_b : _GEN_5554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5556 = 10'hd8 == r_count_7_io_out ? io_r_216_b : _GEN_5555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5557 = 10'hd9 == r_count_7_io_out ? io_r_217_b : _GEN_5556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5558 = 10'hda == r_count_7_io_out ? io_r_218_b : _GEN_5557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5559 = 10'hdb == r_count_7_io_out ? io_r_219_b : _GEN_5558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5560 = 10'hdc == r_count_7_io_out ? io_r_220_b : _GEN_5559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5561 = 10'hdd == r_count_7_io_out ? io_r_221_b : _GEN_5560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5562 = 10'hde == r_count_7_io_out ? io_r_222_b : _GEN_5561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5563 = 10'hdf == r_count_7_io_out ? io_r_223_b : _GEN_5562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5564 = 10'he0 == r_count_7_io_out ? io_r_224_b : _GEN_5563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5565 = 10'he1 == r_count_7_io_out ? io_r_225_b : _GEN_5564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5566 = 10'he2 == r_count_7_io_out ? io_r_226_b : _GEN_5565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5567 = 10'he3 == r_count_7_io_out ? io_r_227_b : _GEN_5566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5568 = 10'he4 == r_count_7_io_out ? io_r_228_b : _GEN_5567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5569 = 10'he5 == r_count_7_io_out ? io_r_229_b : _GEN_5568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5570 = 10'he6 == r_count_7_io_out ? io_r_230_b : _GEN_5569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5571 = 10'he7 == r_count_7_io_out ? io_r_231_b : _GEN_5570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5572 = 10'he8 == r_count_7_io_out ? io_r_232_b : _GEN_5571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5573 = 10'he9 == r_count_7_io_out ? io_r_233_b : _GEN_5572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5574 = 10'hea == r_count_7_io_out ? io_r_234_b : _GEN_5573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5575 = 10'heb == r_count_7_io_out ? io_r_235_b : _GEN_5574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5576 = 10'hec == r_count_7_io_out ? io_r_236_b : _GEN_5575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5577 = 10'hed == r_count_7_io_out ? io_r_237_b : _GEN_5576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5578 = 10'hee == r_count_7_io_out ? io_r_238_b : _GEN_5577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5579 = 10'hef == r_count_7_io_out ? io_r_239_b : _GEN_5578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5580 = 10'hf0 == r_count_7_io_out ? io_r_240_b : _GEN_5579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5581 = 10'hf1 == r_count_7_io_out ? io_r_241_b : _GEN_5580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5582 = 10'hf2 == r_count_7_io_out ? io_r_242_b : _GEN_5581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5583 = 10'hf3 == r_count_7_io_out ? io_r_243_b : _GEN_5582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5584 = 10'hf4 == r_count_7_io_out ? io_r_244_b : _GEN_5583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5585 = 10'hf5 == r_count_7_io_out ? io_r_245_b : _GEN_5584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5586 = 10'hf6 == r_count_7_io_out ? io_r_246_b : _GEN_5585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5587 = 10'hf7 == r_count_7_io_out ? io_r_247_b : _GEN_5586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5588 = 10'hf8 == r_count_7_io_out ? io_r_248_b : _GEN_5587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5589 = 10'hf9 == r_count_7_io_out ? io_r_249_b : _GEN_5588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5590 = 10'hfa == r_count_7_io_out ? io_r_250_b : _GEN_5589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5591 = 10'hfb == r_count_7_io_out ? io_r_251_b : _GEN_5590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5592 = 10'hfc == r_count_7_io_out ? io_r_252_b : _GEN_5591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5593 = 10'hfd == r_count_7_io_out ? io_r_253_b : _GEN_5592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5594 = 10'hfe == r_count_7_io_out ? io_r_254_b : _GEN_5593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5595 = 10'hff == r_count_7_io_out ? io_r_255_b : _GEN_5594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5596 = 10'h100 == r_count_7_io_out ? io_r_256_b : _GEN_5595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5597 = 10'h101 == r_count_7_io_out ? io_r_257_b : _GEN_5596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5598 = 10'h102 == r_count_7_io_out ? io_r_258_b : _GEN_5597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5599 = 10'h103 == r_count_7_io_out ? io_r_259_b : _GEN_5598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5600 = 10'h104 == r_count_7_io_out ? io_r_260_b : _GEN_5599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5601 = 10'h105 == r_count_7_io_out ? io_r_261_b : _GEN_5600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5602 = 10'h106 == r_count_7_io_out ? io_r_262_b : _GEN_5601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5603 = 10'h107 == r_count_7_io_out ? io_r_263_b : _GEN_5602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5604 = 10'h108 == r_count_7_io_out ? io_r_264_b : _GEN_5603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5605 = 10'h109 == r_count_7_io_out ? io_r_265_b : _GEN_5604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5606 = 10'h10a == r_count_7_io_out ? io_r_266_b : _GEN_5605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5607 = 10'h10b == r_count_7_io_out ? io_r_267_b : _GEN_5606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5608 = 10'h10c == r_count_7_io_out ? io_r_268_b : _GEN_5607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5609 = 10'h10d == r_count_7_io_out ? io_r_269_b : _GEN_5608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5610 = 10'h10e == r_count_7_io_out ? io_r_270_b : _GEN_5609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5611 = 10'h10f == r_count_7_io_out ? io_r_271_b : _GEN_5610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5612 = 10'h110 == r_count_7_io_out ? io_r_272_b : _GEN_5611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5613 = 10'h111 == r_count_7_io_out ? io_r_273_b : _GEN_5612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5614 = 10'h112 == r_count_7_io_out ? io_r_274_b : _GEN_5613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5615 = 10'h113 == r_count_7_io_out ? io_r_275_b : _GEN_5614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5616 = 10'h114 == r_count_7_io_out ? io_r_276_b : _GEN_5615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5617 = 10'h115 == r_count_7_io_out ? io_r_277_b : _GEN_5616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5618 = 10'h116 == r_count_7_io_out ? io_r_278_b : _GEN_5617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5619 = 10'h117 == r_count_7_io_out ? io_r_279_b : _GEN_5618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5620 = 10'h118 == r_count_7_io_out ? io_r_280_b : _GEN_5619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5621 = 10'h119 == r_count_7_io_out ? io_r_281_b : _GEN_5620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5622 = 10'h11a == r_count_7_io_out ? io_r_282_b : _GEN_5621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5623 = 10'h11b == r_count_7_io_out ? io_r_283_b : _GEN_5622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5624 = 10'h11c == r_count_7_io_out ? io_r_284_b : _GEN_5623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5625 = 10'h11d == r_count_7_io_out ? io_r_285_b : _GEN_5624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5626 = 10'h11e == r_count_7_io_out ? io_r_286_b : _GEN_5625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5627 = 10'h11f == r_count_7_io_out ? io_r_287_b : _GEN_5626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5628 = 10'h120 == r_count_7_io_out ? io_r_288_b : _GEN_5627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5629 = 10'h121 == r_count_7_io_out ? io_r_289_b : _GEN_5628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5630 = 10'h122 == r_count_7_io_out ? io_r_290_b : _GEN_5629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5631 = 10'h123 == r_count_7_io_out ? io_r_291_b : _GEN_5630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5632 = 10'h124 == r_count_7_io_out ? io_r_292_b : _GEN_5631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5633 = 10'h125 == r_count_7_io_out ? io_r_293_b : _GEN_5632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5634 = 10'h126 == r_count_7_io_out ? io_r_294_b : _GEN_5633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5635 = 10'h127 == r_count_7_io_out ? io_r_295_b : _GEN_5634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5636 = 10'h128 == r_count_7_io_out ? io_r_296_b : _GEN_5635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5637 = 10'h129 == r_count_7_io_out ? io_r_297_b : _GEN_5636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5638 = 10'h12a == r_count_7_io_out ? io_r_298_b : _GEN_5637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5639 = 10'h12b == r_count_7_io_out ? io_r_299_b : _GEN_5638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5640 = 10'h12c == r_count_7_io_out ? io_r_300_b : _GEN_5639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5641 = 10'h12d == r_count_7_io_out ? io_r_301_b : _GEN_5640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5642 = 10'h12e == r_count_7_io_out ? io_r_302_b : _GEN_5641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5643 = 10'h12f == r_count_7_io_out ? io_r_303_b : _GEN_5642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5644 = 10'h130 == r_count_7_io_out ? io_r_304_b : _GEN_5643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5645 = 10'h131 == r_count_7_io_out ? io_r_305_b : _GEN_5644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5646 = 10'h132 == r_count_7_io_out ? io_r_306_b : _GEN_5645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5647 = 10'h133 == r_count_7_io_out ? io_r_307_b : _GEN_5646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5648 = 10'h134 == r_count_7_io_out ? io_r_308_b : _GEN_5647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5649 = 10'h135 == r_count_7_io_out ? io_r_309_b : _GEN_5648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5650 = 10'h136 == r_count_7_io_out ? io_r_310_b : _GEN_5649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5651 = 10'h137 == r_count_7_io_out ? io_r_311_b : _GEN_5650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5652 = 10'h138 == r_count_7_io_out ? io_r_312_b : _GEN_5651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5653 = 10'h139 == r_count_7_io_out ? io_r_313_b : _GEN_5652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5654 = 10'h13a == r_count_7_io_out ? io_r_314_b : _GEN_5653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5655 = 10'h13b == r_count_7_io_out ? io_r_315_b : _GEN_5654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5656 = 10'h13c == r_count_7_io_out ? io_r_316_b : _GEN_5655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5657 = 10'h13d == r_count_7_io_out ? io_r_317_b : _GEN_5656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5658 = 10'h13e == r_count_7_io_out ? io_r_318_b : _GEN_5657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5659 = 10'h13f == r_count_7_io_out ? io_r_319_b : _GEN_5658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5660 = 10'h140 == r_count_7_io_out ? io_r_320_b : _GEN_5659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5661 = 10'h141 == r_count_7_io_out ? io_r_321_b : _GEN_5660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5662 = 10'h142 == r_count_7_io_out ? io_r_322_b : _GEN_5661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5663 = 10'h143 == r_count_7_io_out ? io_r_323_b : _GEN_5662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5664 = 10'h144 == r_count_7_io_out ? io_r_324_b : _GEN_5663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5665 = 10'h145 == r_count_7_io_out ? io_r_325_b : _GEN_5664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5666 = 10'h146 == r_count_7_io_out ? io_r_326_b : _GEN_5665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5667 = 10'h147 == r_count_7_io_out ? io_r_327_b : _GEN_5666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5668 = 10'h148 == r_count_7_io_out ? io_r_328_b : _GEN_5667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5669 = 10'h149 == r_count_7_io_out ? io_r_329_b : _GEN_5668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5670 = 10'h14a == r_count_7_io_out ? io_r_330_b : _GEN_5669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5671 = 10'h14b == r_count_7_io_out ? io_r_331_b : _GEN_5670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5672 = 10'h14c == r_count_7_io_out ? io_r_332_b : _GEN_5671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5673 = 10'h14d == r_count_7_io_out ? io_r_333_b : _GEN_5672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5674 = 10'h14e == r_count_7_io_out ? io_r_334_b : _GEN_5673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5675 = 10'h14f == r_count_7_io_out ? io_r_335_b : _GEN_5674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5676 = 10'h150 == r_count_7_io_out ? io_r_336_b : _GEN_5675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5677 = 10'h151 == r_count_7_io_out ? io_r_337_b : _GEN_5676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5678 = 10'h152 == r_count_7_io_out ? io_r_338_b : _GEN_5677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5679 = 10'h153 == r_count_7_io_out ? io_r_339_b : _GEN_5678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5680 = 10'h154 == r_count_7_io_out ? io_r_340_b : _GEN_5679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5681 = 10'h155 == r_count_7_io_out ? io_r_341_b : _GEN_5680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5682 = 10'h156 == r_count_7_io_out ? io_r_342_b : _GEN_5681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5683 = 10'h157 == r_count_7_io_out ? io_r_343_b : _GEN_5682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5684 = 10'h158 == r_count_7_io_out ? io_r_344_b : _GEN_5683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5685 = 10'h159 == r_count_7_io_out ? io_r_345_b : _GEN_5684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5686 = 10'h15a == r_count_7_io_out ? io_r_346_b : _GEN_5685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5687 = 10'h15b == r_count_7_io_out ? io_r_347_b : _GEN_5686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5688 = 10'h15c == r_count_7_io_out ? io_r_348_b : _GEN_5687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5689 = 10'h15d == r_count_7_io_out ? io_r_349_b : _GEN_5688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5690 = 10'h15e == r_count_7_io_out ? io_r_350_b : _GEN_5689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5691 = 10'h15f == r_count_7_io_out ? io_r_351_b : _GEN_5690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5692 = 10'h160 == r_count_7_io_out ? io_r_352_b : _GEN_5691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5693 = 10'h161 == r_count_7_io_out ? io_r_353_b : _GEN_5692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5694 = 10'h162 == r_count_7_io_out ? io_r_354_b : _GEN_5693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5695 = 10'h163 == r_count_7_io_out ? io_r_355_b : _GEN_5694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5696 = 10'h164 == r_count_7_io_out ? io_r_356_b : _GEN_5695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5697 = 10'h165 == r_count_7_io_out ? io_r_357_b : _GEN_5696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5698 = 10'h166 == r_count_7_io_out ? io_r_358_b : _GEN_5697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5699 = 10'h167 == r_count_7_io_out ? io_r_359_b : _GEN_5698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5700 = 10'h168 == r_count_7_io_out ? io_r_360_b : _GEN_5699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5701 = 10'h169 == r_count_7_io_out ? io_r_361_b : _GEN_5700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5702 = 10'h16a == r_count_7_io_out ? io_r_362_b : _GEN_5701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5703 = 10'h16b == r_count_7_io_out ? io_r_363_b : _GEN_5702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5704 = 10'h16c == r_count_7_io_out ? io_r_364_b : _GEN_5703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5705 = 10'h16d == r_count_7_io_out ? io_r_365_b : _GEN_5704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5706 = 10'h16e == r_count_7_io_out ? io_r_366_b : _GEN_5705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5707 = 10'h16f == r_count_7_io_out ? io_r_367_b : _GEN_5706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5708 = 10'h170 == r_count_7_io_out ? io_r_368_b : _GEN_5707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5709 = 10'h171 == r_count_7_io_out ? io_r_369_b : _GEN_5708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5710 = 10'h172 == r_count_7_io_out ? io_r_370_b : _GEN_5709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5711 = 10'h173 == r_count_7_io_out ? io_r_371_b : _GEN_5710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5712 = 10'h174 == r_count_7_io_out ? io_r_372_b : _GEN_5711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5713 = 10'h175 == r_count_7_io_out ? io_r_373_b : _GEN_5712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5714 = 10'h176 == r_count_7_io_out ? io_r_374_b : _GEN_5713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5715 = 10'h177 == r_count_7_io_out ? io_r_375_b : _GEN_5714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5716 = 10'h178 == r_count_7_io_out ? io_r_376_b : _GEN_5715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5717 = 10'h179 == r_count_7_io_out ? io_r_377_b : _GEN_5716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5718 = 10'h17a == r_count_7_io_out ? io_r_378_b : _GEN_5717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5719 = 10'h17b == r_count_7_io_out ? io_r_379_b : _GEN_5718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5720 = 10'h17c == r_count_7_io_out ? io_r_380_b : _GEN_5719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5721 = 10'h17d == r_count_7_io_out ? io_r_381_b : _GEN_5720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5722 = 10'h17e == r_count_7_io_out ? io_r_382_b : _GEN_5721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5723 = 10'h17f == r_count_7_io_out ? io_r_383_b : _GEN_5722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5724 = 10'h180 == r_count_7_io_out ? io_r_384_b : _GEN_5723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5725 = 10'h181 == r_count_7_io_out ? io_r_385_b : _GEN_5724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5726 = 10'h182 == r_count_7_io_out ? io_r_386_b : _GEN_5725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5727 = 10'h183 == r_count_7_io_out ? io_r_387_b : _GEN_5726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5728 = 10'h184 == r_count_7_io_out ? io_r_388_b : _GEN_5727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5729 = 10'h185 == r_count_7_io_out ? io_r_389_b : _GEN_5728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5730 = 10'h186 == r_count_7_io_out ? io_r_390_b : _GEN_5729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5731 = 10'h187 == r_count_7_io_out ? io_r_391_b : _GEN_5730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5732 = 10'h188 == r_count_7_io_out ? io_r_392_b : _GEN_5731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5733 = 10'h189 == r_count_7_io_out ? io_r_393_b : _GEN_5732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5734 = 10'h18a == r_count_7_io_out ? io_r_394_b : _GEN_5733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5735 = 10'h18b == r_count_7_io_out ? io_r_395_b : _GEN_5734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5736 = 10'h18c == r_count_7_io_out ? io_r_396_b : _GEN_5735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5737 = 10'h18d == r_count_7_io_out ? io_r_397_b : _GEN_5736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5738 = 10'h18e == r_count_7_io_out ? io_r_398_b : _GEN_5737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5739 = 10'h18f == r_count_7_io_out ? io_r_399_b : _GEN_5738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5740 = 10'h190 == r_count_7_io_out ? io_r_400_b : _GEN_5739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5741 = 10'h191 == r_count_7_io_out ? io_r_401_b : _GEN_5740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5742 = 10'h192 == r_count_7_io_out ? io_r_402_b : _GEN_5741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5743 = 10'h193 == r_count_7_io_out ? io_r_403_b : _GEN_5742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5744 = 10'h194 == r_count_7_io_out ? io_r_404_b : _GEN_5743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5745 = 10'h195 == r_count_7_io_out ? io_r_405_b : _GEN_5744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5746 = 10'h196 == r_count_7_io_out ? io_r_406_b : _GEN_5745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5747 = 10'h197 == r_count_7_io_out ? io_r_407_b : _GEN_5746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5748 = 10'h198 == r_count_7_io_out ? io_r_408_b : _GEN_5747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5749 = 10'h199 == r_count_7_io_out ? io_r_409_b : _GEN_5748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5750 = 10'h19a == r_count_7_io_out ? io_r_410_b : _GEN_5749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5751 = 10'h19b == r_count_7_io_out ? io_r_411_b : _GEN_5750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5752 = 10'h19c == r_count_7_io_out ? io_r_412_b : _GEN_5751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5753 = 10'h19d == r_count_7_io_out ? io_r_413_b : _GEN_5752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5754 = 10'h19e == r_count_7_io_out ? io_r_414_b : _GEN_5753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5755 = 10'h19f == r_count_7_io_out ? io_r_415_b : _GEN_5754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5756 = 10'h1a0 == r_count_7_io_out ? io_r_416_b : _GEN_5755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5757 = 10'h1a1 == r_count_7_io_out ? io_r_417_b : _GEN_5756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5758 = 10'h1a2 == r_count_7_io_out ? io_r_418_b : _GEN_5757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5759 = 10'h1a3 == r_count_7_io_out ? io_r_419_b : _GEN_5758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5760 = 10'h1a4 == r_count_7_io_out ? io_r_420_b : _GEN_5759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5761 = 10'h1a5 == r_count_7_io_out ? io_r_421_b : _GEN_5760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5762 = 10'h1a6 == r_count_7_io_out ? io_r_422_b : _GEN_5761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5763 = 10'h1a7 == r_count_7_io_out ? io_r_423_b : _GEN_5762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5764 = 10'h1a8 == r_count_7_io_out ? io_r_424_b : _GEN_5763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5765 = 10'h1a9 == r_count_7_io_out ? io_r_425_b : _GEN_5764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5766 = 10'h1aa == r_count_7_io_out ? io_r_426_b : _GEN_5765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5767 = 10'h1ab == r_count_7_io_out ? io_r_427_b : _GEN_5766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5768 = 10'h1ac == r_count_7_io_out ? io_r_428_b : _GEN_5767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5769 = 10'h1ad == r_count_7_io_out ? io_r_429_b : _GEN_5768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5770 = 10'h1ae == r_count_7_io_out ? io_r_430_b : _GEN_5769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5771 = 10'h1af == r_count_7_io_out ? io_r_431_b : _GEN_5770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5772 = 10'h1b0 == r_count_7_io_out ? io_r_432_b : _GEN_5771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5773 = 10'h1b1 == r_count_7_io_out ? io_r_433_b : _GEN_5772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5774 = 10'h1b2 == r_count_7_io_out ? io_r_434_b : _GEN_5773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5775 = 10'h1b3 == r_count_7_io_out ? io_r_435_b : _GEN_5774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5776 = 10'h1b4 == r_count_7_io_out ? io_r_436_b : _GEN_5775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5777 = 10'h1b5 == r_count_7_io_out ? io_r_437_b : _GEN_5776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5778 = 10'h1b6 == r_count_7_io_out ? io_r_438_b : _GEN_5777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5779 = 10'h1b7 == r_count_7_io_out ? io_r_439_b : _GEN_5778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5780 = 10'h1b8 == r_count_7_io_out ? io_r_440_b : _GEN_5779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5781 = 10'h1b9 == r_count_7_io_out ? io_r_441_b : _GEN_5780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5782 = 10'h1ba == r_count_7_io_out ? io_r_442_b : _GEN_5781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5783 = 10'h1bb == r_count_7_io_out ? io_r_443_b : _GEN_5782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5784 = 10'h1bc == r_count_7_io_out ? io_r_444_b : _GEN_5783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5785 = 10'h1bd == r_count_7_io_out ? io_r_445_b : _GEN_5784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5786 = 10'h1be == r_count_7_io_out ? io_r_446_b : _GEN_5785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5787 = 10'h1bf == r_count_7_io_out ? io_r_447_b : _GEN_5786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5788 = 10'h1c0 == r_count_7_io_out ? io_r_448_b : _GEN_5787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5789 = 10'h1c1 == r_count_7_io_out ? io_r_449_b : _GEN_5788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5790 = 10'h1c2 == r_count_7_io_out ? io_r_450_b : _GEN_5789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5791 = 10'h1c3 == r_count_7_io_out ? io_r_451_b : _GEN_5790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5792 = 10'h1c4 == r_count_7_io_out ? io_r_452_b : _GEN_5791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5793 = 10'h1c5 == r_count_7_io_out ? io_r_453_b : _GEN_5792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5794 = 10'h1c6 == r_count_7_io_out ? io_r_454_b : _GEN_5793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5795 = 10'h1c7 == r_count_7_io_out ? io_r_455_b : _GEN_5794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5796 = 10'h1c8 == r_count_7_io_out ? io_r_456_b : _GEN_5795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5797 = 10'h1c9 == r_count_7_io_out ? io_r_457_b : _GEN_5796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5798 = 10'h1ca == r_count_7_io_out ? io_r_458_b : _GEN_5797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5799 = 10'h1cb == r_count_7_io_out ? io_r_459_b : _GEN_5798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5800 = 10'h1cc == r_count_7_io_out ? io_r_460_b : _GEN_5799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5801 = 10'h1cd == r_count_7_io_out ? io_r_461_b : _GEN_5800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5802 = 10'h1ce == r_count_7_io_out ? io_r_462_b : _GEN_5801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5803 = 10'h1cf == r_count_7_io_out ? io_r_463_b : _GEN_5802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5804 = 10'h1d0 == r_count_7_io_out ? io_r_464_b : _GEN_5803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5805 = 10'h1d1 == r_count_7_io_out ? io_r_465_b : _GEN_5804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5806 = 10'h1d2 == r_count_7_io_out ? io_r_466_b : _GEN_5805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5807 = 10'h1d3 == r_count_7_io_out ? io_r_467_b : _GEN_5806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5808 = 10'h1d4 == r_count_7_io_out ? io_r_468_b : _GEN_5807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5809 = 10'h1d5 == r_count_7_io_out ? io_r_469_b : _GEN_5808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5810 = 10'h1d6 == r_count_7_io_out ? io_r_470_b : _GEN_5809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5811 = 10'h1d7 == r_count_7_io_out ? io_r_471_b : _GEN_5810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5812 = 10'h1d8 == r_count_7_io_out ? io_r_472_b : _GEN_5811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5813 = 10'h1d9 == r_count_7_io_out ? io_r_473_b : _GEN_5812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5814 = 10'h1da == r_count_7_io_out ? io_r_474_b : _GEN_5813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5815 = 10'h1db == r_count_7_io_out ? io_r_475_b : _GEN_5814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5816 = 10'h1dc == r_count_7_io_out ? io_r_476_b : _GEN_5815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5817 = 10'h1dd == r_count_7_io_out ? io_r_477_b : _GEN_5816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5818 = 10'h1de == r_count_7_io_out ? io_r_478_b : _GEN_5817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5819 = 10'h1df == r_count_7_io_out ? io_r_479_b : _GEN_5818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5820 = 10'h1e0 == r_count_7_io_out ? io_r_480_b : _GEN_5819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5821 = 10'h1e1 == r_count_7_io_out ? io_r_481_b : _GEN_5820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5822 = 10'h1e2 == r_count_7_io_out ? io_r_482_b : _GEN_5821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5823 = 10'h1e3 == r_count_7_io_out ? io_r_483_b : _GEN_5822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5824 = 10'h1e4 == r_count_7_io_out ? io_r_484_b : _GEN_5823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5825 = 10'h1e5 == r_count_7_io_out ? io_r_485_b : _GEN_5824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5826 = 10'h1e6 == r_count_7_io_out ? io_r_486_b : _GEN_5825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5827 = 10'h1e7 == r_count_7_io_out ? io_r_487_b : _GEN_5826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5828 = 10'h1e8 == r_count_7_io_out ? io_r_488_b : _GEN_5827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5829 = 10'h1e9 == r_count_7_io_out ? io_r_489_b : _GEN_5828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5830 = 10'h1ea == r_count_7_io_out ? io_r_490_b : _GEN_5829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5831 = 10'h1eb == r_count_7_io_out ? io_r_491_b : _GEN_5830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5832 = 10'h1ec == r_count_7_io_out ? io_r_492_b : _GEN_5831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5833 = 10'h1ed == r_count_7_io_out ? io_r_493_b : _GEN_5832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5834 = 10'h1ee == r_count_7_io_out ? io_r_494_b : _GEN_5833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5835 = 10'h1ef == r_count_7_io_out ? io_r_495_b : _GEN_5834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5836 = 10'h1f0 == r_count_7_io_out ? io_r_496_b : _GEN_5835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5837 = 10'h1f1 == r_count_7_io_out ? io_r_497_b : _GEN_5836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5838 = 10'h1f2 == r_count_7_io_out ? io_r_498_b : _GEN_5837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5839 = 10'h1f3 == r_count_7_io_out ? io_r_499_b : _GEN_5838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5840 = 10'h1f4 == r_count_7_io_out ? io_r_500_b : _GEN_5839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5841 = 10'h1f5 == r_count_7_io_out ? io_r_501_b : _GEN_5840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5842 = 10'h1f6 == r_count_7_io_out ? io_r_502_b : _GEN_5841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5843 = 10'h1f7 == r_count_7_io_out ? io_r_503_b : _GEN_5842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5844 = 10'h1f8 == r_count_7_io_out ? io_r_504_b : _GEN_5843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5845 = 10'h1f9 == r_count_7_io_out ? io_r_505_b : _GEN_5844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5846 = 10'h1fa == r_count_7_io_out ? io_r_506_b : _GEN_5845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5847 = 10'h1fb == r_count_7_io_out ? io_r_507_b : _GEN_5846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5848 = 10'h1fc == r_count_7_io_out ? io_r_508_b : _GEN_5847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5849 = 10'h1fd == r_count_7_io_out ? io_r_509_b : _GEN_5848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5850 = 10'h1fe == r_count_7_io_out ? io_r_510_b : _GEN_5849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5851 = 10'h1ff == r_count_7_io_out ? io_r_511_b : _GEN_5850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5852 = 10'h200 == r_count_7_io_out ? io_r_512_b : _GEN_5851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5853 = 10'h201 == r_count_7_io_out ? io_r_513_b : _GEN_5852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5854 = 10'h202 == r_count_7_io_out ? io_r_514_b : _GEN_5853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5855 = 10'h203 == r_count_7_io_out ? io_r_515_b : _GEN_5854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5856 = 10'h204 == r_count_7_io_out ? io_r_516_b : _GEN_5855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5857 = 10'h205 == r_count_7_io_out ? io_r_517_b : _GEN_5856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5858 = 10'h206 == r_count_7_io_out ? io_r_518_b : _GEN_5857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5859 = 10'h207 == r_count_7_io_out ? io_r_519_b : _GEN_5858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5860 = 10'h208 == r_count_7_io_out ? io_r_520_b : _GEN_5859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5861 = 10'h209 == r_count_7_io_out ? io_r_521_b : _GEN_5860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5862 = 10'h20a == r_count_7_io_out ? io_r_522_b : _GEN_5861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5863 = 10'h20b == r_count_7_io_out ? io_r_523_b : _GEN_5862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5864 = 10'h20c == r_count_7_io_out ? io_r_524_b : _GEN_5863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5865 = 10'h20d == r_count_7_io_out ? io_r_525_b : _GEN_5864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5866 = 10'h20e == r_count_7_io_out ? io_r_526_b : _GEN_5865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5867 = 10'h20f == r_count_7_io_out ? io_r_527_b : _GEN_5866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5868 = 10'h210 == r_count_7_io_out ? io_r_528_b : _GEN_5867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5869 = 10'h211 == r_count_7_io_out ? io_r_529_b : _GEN_5868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5870 = 10'h212 == r_count_7_io_out ? io_r_530_b : _GEN_5869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5871 = 10'h213 == r_count_7_io_out ? io_r_531_b : _GEN_5870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5872 = 10'h214 == r_count_7_io_out ? io_r_532_b : _GEN_5871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5873 = 10'h215 == r_count_7_io_out ? io_r_533_b : _GEN_5872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5874 = 10'h216 == r_count_7_io_out ? io_r_534_b : _GEN_5873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5875 = 10'h217 == r_count_7_io_out ? io_r_535_b : _GEN_5874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5876 = 10'h218 == r_count_7_io_out ? io_r_536_b : _GEN_5875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5877 = 10'h219 == r_count_7_io_out ? io_r_537_b : _GEN_5876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5878 = 10'h21a == r_count_7_io_out ? io_r_538_b : _GEN_5877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5879 = 10'h21b == r_count_7_io_out ? io_r_539_b : _GEN_5878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5880 = 10'h21c == r_count_7_io_out ? io_r_540_b : _GEN_5879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5881 = 10'h21d == r_count_7_io_out ? io_r_541_b : _GEN_5880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5882 = 10'h21e == r_count_7_io_out ? io_r_542_b : _GEN_5881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5883 = 10'h21f == r_count_7_io_out ? io_r_543_b : _GEN_5882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5884 = 10'h220 == r_count_7_io_out ? io_r_544_b : _GEN_5883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5885 = 10'h221 == r_count_7_io_out ? io_r_545_b : _GEN_5884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5886 = 10'h222 == r_count_7_io_out ? io_r_546_b : _GEN_5885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5887 = 10'h223 == r_count_7_io_out ? io_r_547_b : _GEN_5886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5888 = 10'h224 == r_count_7_io_out ? io_r_548_b : _GEN_5887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5889 = 10'h225 == r_count_7_io_out ? io_r_549_b : _GEN_5888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5890 = 10'h226 == r_count_7_io_out ? io_r_550_b : _GEN_5889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5891 = 10'h227 == r_count_7_io_out ? io_r_551_b : _GEN_5890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5892 = 10'h228 == r_count_7_io_out ? io_r_552_b : _GEN_5891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5893 = 10'h229 == r_count_7_io_out ? io_r_553_b : _GEN_5892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5894 = 10'h22a == r_count_7_io_out ? io_r_554_b : _GEN_5893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5895 = 10'h22b == r_count_7_io_out ? io_r_555_b : _GEN_5894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5896 = 10'h22c == r_count_7_io_out ? io_r_556_b : _GEN_5895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5897 = 10'h22d == r_count_7_io_out ? io_r_557_b : _GEN_5896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5898 = 10'h22e == r_count_7_io_out ? io_r_558_b : _GEN_5897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5899 = 10'h22f == r_count_7_io_out ? io_r_559_b : _GEN_5898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5900 = 10'h230 == r_count_7_io_out ? io_r_560_b : _GEN_5899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5901 = 10'h231 == r_count_7_io_out ? io_r_561_b : _GEN_5900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5902 = 10'h232 == r_count_7_io_out ? io_r_562_b : _GEN_5901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5903 = 10'h233 == r_count_7_io_out ? io_r_563_b : _GEN_5902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5904 = 10'h234 == r_count_7_io_out ? io_r_564_b : _GEN_5903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5905 = 10'h235 == r_count_7_io_out ? io_r_565_b : _GEN_5904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5906 = 10'h236 == r_count_7_io_out ? io_r_566_b : _GEN_5905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5907 = 10'h237 == r_count_7_io_out ? io_r_567_b : _GEN_5906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5908 = 10'h238 == r_count_7_io_out ? io_r_568_b : _GEN_5907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5909 = 10'h239 == r_count_7_io_out ? io_r_569_b : _GEN_5908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5910 = 10'h23a == r_count_7_io_out ? io_r_570_b : _GEN_5909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5911 = 10'h23b == r_count_7_io_out ? io_r_571_b : _GEN_5910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5912 = 10'h23c == r_count_7_io_out ? io_r_572_b : _GEN_5911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5913 = 10'h23d == r_count_7_io_out ? io_r_573_b : _GEN_5912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5914 = 10'h23e == r_count_7_io_out ? io_r_574_b : _GEN_5913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5915 = 10'h23f == r_count_7_io_out ? io_r_575_b : _GEN_5914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5916 = 10'h240 == r_count_7_io_out ? io_r_576_b : _GEN_5915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5917 = 10'h241 == r_count_7_io_out ? io_r_577_b : _GEN_5916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5918 = 10'h242 == r_count_7_io_out ? io_r_578_b : _GEN_5917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5919 = 10'h243 == r_count_7_io_out ? io_r_579_b : _GEN_5918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5920 = 10'h244 == r_count_7_io_out ? io_r_580_b : _GEN_5919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5921 = 10'h245 == r_count_7_io_out ? io_r_581_b : _GEN_5920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5922 = 10'h246 == r_count_7_io_out ? io_r_582_b : _GEN_5921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5923 = 10'h247 == r_count_7_io_out ? io_r_583_b : _GEN_5922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5924 = 10'h248 == r_count_7_io_out ? io_r_584_b : _GEN_5923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5925 = 10'h249 == r_count_7_io_out ? io_r_585_b : _GEN_5924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5926 = 10'h24a == r_count_7_io_out ? io_r_586_b : _GEN_5925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5927 = 10'h24b == r_count_7_io_out ? io_r_587_b : _GEN_5926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5928 = 10'h24c == r_count_7_io_out ? io_r_588_b : _GEN_5927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5929 = 10'h24d == r_count_7_io_out ? io_r_589_b : _GEN_5928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5930 = 10'h24e == r_count_7_io_out ? io_r_590_b : _GEN_5929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5931 = 10'h24f == r_count_7_io_out ? io_r_591_b : _GEN_5930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5932 = 10'h250 == r_count_7_io_out ? io_r_592_b : _GEN_5931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5933 = 10'h251 == r_count_7_io_out ? io_r_593_b : _GEN_5932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5934 = 10'h252 == r_count_7_io_out ? io_r_594_b : _GEN_5933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5935 = 10'h253 == r_count_7_io_out ? io_r_595_b : _GEN_5934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5936 = 10'h254 == r_count_7_io_out ? io_r_596_b : _GEN_5935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5937 = 10'h255 == r_count_7_io_out ? io_r_597_b : _GEN_5936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5938 = 10'h256 == r_count_7_io_out ? io_r_598_b : _GEN_5937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5939 = 10'h257 == r_count_7_io_out ? io_r_599_b : _GEN_5938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5940 = 10'h258 == r_count_7_io_out ? io_r_600_b : _GEN_5939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5941 = 10'h259 == r_count_7_io_out ? io_r_601_b : _GEN_5940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5942 = 10'h25a == r_count_7_io_out ? io_r_602_b : _GEN_5941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5943 = 10'h25b == r_count_7_io_out ? io_r_603_b : _GEN_5942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5944 = 10'h25c == r_count_7_io_out ? io_r_604_b : _GEN_5943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5945 = 10'h25d == r_count_7_io_out ? io_r_605_b : _GEN_5944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5946 = 10'h25e == r_count_7_io_out ? io_r_606_b : _GEN_5945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5947 = 10'h25f == r_count_7_io_out ? io_r_607_b : _GEN_5946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5948 = 10'h260 == r_count_7_io_out ? io_r_608_b : _GEN_5947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5949 = 10'h261 == r_count_7_io_out ? io_r_609_b : _GEN_5948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5950 = 10'h262 == r_count_7_io_out ? io_r_610_b : _GEN_5949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5951 = 10'h263 == r_count_7_io_out ? io_r_611_b : _GEN_5950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5952 = 10'h264 == r_count_7_io_out ? io_r_612_b : _GEN_5951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5953 = 10'h265 == r_count_7_io_out ? io_r_613_b : _GEN_5952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5954 = 10'h266 == r_count_7_io_out ? io_r_614_b : _GEN_5953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5955 = 10'h267 == r_count_7_io_out ? io_r_615_b : _GEN_5954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5956 = 10'h268 == r_count_7_io_out ? io_r_616_b : _GEN_5955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5957 = 10'h269 == r_count_7_io_out ? io_r_617_b : _GEN_5956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5958 = 10'h26a == r_count_7_io_out ? io_r_618_b : _GEN_5957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5959 = 10'h26b == r_count_7_io_out ? io_r_619_b : _GEN_5958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5960 = 10'h26c == r_count_7_io_out ? io_r_620_b : _GEN_5959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5961 = 10'h26d == r_count_7_io_out ? io_r_621_b : _GEN_5960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5962 = 10'h26e == r_count_7_io_out ? io_r_622_b : _GEN_5961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5963 = 10'h26f == r_count_7_io_out ? io_r_623_b : _GEN_5962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5964 = 10'h270 == r_count_7_io_out ? io_r_624_b : _GEN_5963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5965 = 10'h271 == r_count_7_io_out ? io_r_625_b : _GEN_5964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5966 = 10'h272 == r_count_7_io_out ? io_r_626_b : _GEN_5965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5967 = 10'h273 == r_count_7_io_out ? io_r_627_b : _GEN_5966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5968 = 10'h274 == r_count_7_io_out ? io_r_628_b : _GEN_5967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5969 = 10'h275 == r_count_7_io_out ? io_r_629_b : _GEN_5968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5970 = 10'h276 == r_count_7_io_out ? io_r_630_b : _GEN_5969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5971 = 10'h277 == r_count_7_io_out ? io_r_631_b : _GEN_5970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5972 = 10'h278 == r_count_7_io_out ? io_r_632_b : _GEN_5971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5973 = 10'h279 == r_count_7_io_out ? io_r_633_b : _GEN_5972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5974 = 10'h27a == r_count_7_io_out ? io_r_634_b : _GEN_5973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5975 = 10'h27b == r_count_7_io_out ? io_r_635_b : _GEN_5974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5976 = 10'h27c == r_count_7_io_out ? io_r_636_b : _GEN_5975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5977 = 10'h27d == r_count_7_io_out ? io_r_637_b : _GEN_5976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5978 = 10'h27e == r_count_7_io_out ? io_r_638_b : _GEN_5977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5979 = 10'h27f == r_count_7_io_out ? io_r_639_b : _GEN_5978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5980 = 10'h280 == r_count_7_io_out ? io_r_640_b : _GEN_5979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5981 = 10'h281 == r_count_7_io_out ? io_r_641_b : _GEN_5980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5982 = 10'h282 == r_count_7_io_out ? io_r_642_b : _GEN_5981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5983 = 10'h283 == r_count_7_io_out ? io_r_643_b : _GEN_5982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5984 = 10'h284 == r_count_7_io_out ? io_r_644_b : _GEN_5983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5985 = 10'h285 == r_count_7_io_out ? io_r_645_b : _GEN_5984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5986 = 10'h286 == r_count_7_io_out ? io_r_646_b : _GEN_5985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5987 = 10'h287 == r_count_7_io_out ? io_r_647_b : _GEN_5986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5988 = 10'h288 == r_count_7_io_out ? io_r_648_b : _GEN_5987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5989 = 10'h289 == r_count_7_io_out ? io_r_649_b : _GEN_5988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5990 = 10'h28a == r_count_7_io_out ? io_r_650_b : _GEN_5989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5991 = 10'h28b == r_count_7_io_out ? io_r_651_b : _GEN_5990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5992 = 10'h28c == r_count_7_io_out ? io_r_652_b : _GEN_5991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5993 = 10'h28d == r_count_7_io_out ? io_r_653_b : _GEN_5992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5994 = 10'h28e == r_count_7_io_out ? io_r_654_b : _GEN_5993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5995 = 10'h28f == r_count_7_io_out ? io_r_655_b : _GEN_5994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5996 = 10'h290 == r_count_7_io_out ? io_r_656_b : _GEN_5995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5997 = 10'h291 == r_count_7_io_out ? io_r_657_b : _GEN_5996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5998 = 10'h292 == r_count_7_io_out ? io_r_658_b : _GEN_5997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5999 = 10'h293 == r_count_7_io_out ? io_r_659_b : _GEN_5998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6000 = 10'h294 == r_count_7_io_out ? io_r_660_b : _GEN_5999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6001 = 10'h295 == r_count_7_io_out ? io_r_661_b : _GEN_6000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6002 = 10'h296 == r_count_7_io_out ? io_r_662_b : _GEN_6001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6003 = 10'h297 == r_count_7_io_out ? io_r_663_b : _GEN_6002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6004 = 10'h298 == r_count_7_io_out ? io_r_664_b : _GEN_6003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6005 = 10'h299 == r_count_7_io_out ? io_r_665_b : _GEN_6004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6006 = 10'h29a == r_count_7_io_out ? io_r_666_b : _GEN_6005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6007 = 10'h29b == r_count_7_io_out ? io_r_667_b : _GEN_6006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6008 = 10'h29c == r_count_7_io_out ? io_r_668_b : _GEN_6007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6009 = 10'h29d == r_count_7_io_out ? io_r_669_b : _GEN_6008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6010 = 10'h29e == r_count_7_io_out ? io_r_670_b : _GEN_6009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6011 = 10'h29f == r_count_7_io_out ? io_r_671_b : _GEN_6010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6012 = 10'h2a0 == r_count_7_io_out ? io_r_672_b : _GEN_6011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6013 = 10'h2a1 == r_count_7_io_out ? io_r_673_b : _GEN_6012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6014 = 10'h2a2 == r_count_7_io_out ? io_r_674_b : _GEN_6013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6015 = 10'h2a3 == r_count_7_io_out ? io_r_675_b : _GEN_6014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6016 = 10'h2a4 == r_count_7_io_out ? io_r_676_b : _GEN_6015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6017 = 10'h2a5 == r_count_7_io_out ? io_r_677_b : _GEN_6016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6018 = 10'h2a6 == r_count_7_io_out ? io_r_678_b : _GEN_6017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6019 = 10'h2a7 == r_count_7_io_out ? io_r_679_b : _GEN_6018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6020 = 10'h2a8 == r_count_7_io_out ? io_r_680_b : _GEN_6019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6021 = 10'h2a9 == r_count_7_io_out ? io_r_681_b : _GEN_6020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6022 = 10'h2aa == r_count_7_io_out ? io_r_682_b : _GEN_6021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6023 = 10'h2ab == r_count_7_io_out ? io_r_683_b : _GEN_6022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6024 = 10'h2ac == r_count_7_io_out ? io_r_684_b : _GEN_6023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6025 = 10'h2ad == r_count_7_io_out ? io_r_685_b : _GEN_6024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6026 = 10'h2ae == r_count_7_io_out ? io_r_686_b : _GEN_6025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6027 = 10'h2af == r_count_7_io_out ? io_r_687_b : _GEN_6026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6028 = 10'h2b0 == r_count_7_io_out ? io_r_688_b : _GEN_6027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6029 = 10'h2b1 == r_count_7_io_out ? io_r_689_b : _GEN_6028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6030 = 10'h2b2 == r_count_7_io_out ? io_r_690_b : _GEN_6029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6031 = 10'h2b3 == r_count_7_io_out ? io_r_691_b : _GEN_6030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6032 = 10'h2b4 == r_count_7_io_out ? io_r_692_b : _GEN_6031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6033 = 10'h2b5 == r_count_7_io_out ? io_r_693_b : _GEN_6032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6034 = 10'h2b6 == r_count_7_io_out ? io_r_694_b : _GEN_6033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6035 = 10'h2b7 == r_count_7_io_out ? io_r_695_b : _GEN_6034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6036 = 10'h2b8 == r_count_7_io_out ? io_r_696_b : _GEN_6035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6037 = 10'h2b9 == r_count_7_io_out ? io_r_697_b : _GEN_6036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6038 = 10'h2ba == r_count_7_io_out ? io_r_698_b : _GEN_6037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6039 = 10'h2bb == r_count_7_io_out ? io_r_699_b : _GEN_6038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6040 = 10'h2bc == r_count_7_io_out ? io_r_700_b : _GEN_6039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6041 = 10'h2bd == r_count_7_io_out ? io_r_701_b : _GEN_6040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6042 = 10'h2be == r_count_7_io_out ? io_r_702_b : _GEN_6041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6043 = 10'h2bf == r_count_7_io_out ? io_r_703_b : _GEN_6042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6044 = 10'h2c0 == r_count_7_io_out ? io_r_704_b : _GEN_6043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6045 = 10'h2c1 == r_count_7_io_out ? io_r_705_b : _GEN_6044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6046 = 10'h2c2 == r_count_7_io_out ? io_r_706_b : _GEN_6045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6047 = 10'h2c3 == r_count_7_io_out ? io_r_707_b : _GEN_6046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6048 = 10'h2c4 == r_count_7_io_out ? io_r_708_b : _GEN_6047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6049 = 10'h2c5 == r_count_7_io_out ? io_r_709_b : _GEN_6048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6050 = 10'h2c6 == r_count_7_io_out ? io_r_710_b : _GEN_6049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6051 = 10'h2c7 == r_count_7_io_out ? io_r_711_b : _GEN_6050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6052 = 10'h2c8 == r_count_7_io_out ? io_r_712_b : _GEN_6051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6053 = 10'h2c9 == r_count_7_io_out ? io_r_713_b : _GEN_6052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6054 = 10'h2ca == r_count_7_io_out ? io_r_714_b : _GEN_6053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6055 = 10'h2cb == r_count_7_io_out ? io_r_715_b : _GEN_6054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6056 = 10'h2cc == r_count_7_io_out ? io_r_716_b : _GEN_6055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6057 = 10'h2cd == r_count_7_io_out ? io_r_717_b : _GEN_6056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6058 = 10'h2ce == r_count_7_io_out ? io_r_718_b : _GEN_6057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6059 = 10'h2cf == r_count_7_io_out ? io_r_719_b : _GEN_6058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6060 = 10'h2d0 == r_count_7_io_out ? io_r_720_b : _GEN_6059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6061 = 10'h2d1 == r_count_7_io_out ? io_r_721_b : _GEN_6060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6062 = 10'h2d2 == r_count_7_io_out ? io_r_722_b : _GEN_6061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6063 = 10'h2d3 == r_count_7_io_out ? io_r_723_b : _GEN_6062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6064 = 10'h2d4 == r_count_7_io_out ? io_r_724_b : _GEN_6063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6065 = 10'h2d5 == r_count_7_io_out ? io_r_725_b : _GEN_6064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6066 = 10'h2d6 == r_count_7_io_out ? io_r_726_b : _GEN_6065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6067 = 10'h2d7 == r_count_7_io_out ? io_r_727_b : _GEN_6066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6068 = 10'h2d8 == r_count_7_io_out ? io_r_728_b : _GEN_6067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6069 = 10'h2d9 == r_count_7_io_out ? io_r_729_b : _GEN_6068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6070 = 10'h2da == r_count_7_io_out ? io_r_730_b : _GEN_6069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6071 = 10'h2db == r_count_7_io_out ? io_r_731_b : _GEN_6070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6072 = 10'h2dc == r_count_7_io_out ? io_r_732_b : _GEN_6071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6073 = 10'h2dd == r_count_7_io_out ? io_r_733_b : _GEN_6072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6074 = 10'h2de == r_count_7_io_out ? io_r_734_b : _GEN_6073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6075 = 10'h2df == r_count_7_io_out ? io_r_735_b : _GEN_6074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6076 = 10'h2e0 == r_count_7_io_out ? io_r_736_b : _GEN_6075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6077 = 10'h2e1 == r_count_7_io_out ? io_r_737_b : _GEN_6076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6078 = 10'h2e2 == r_count_7_io_out ? io_r_738_b : _GEN_6077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6079 = 10'h2e3 == r_count_7_io_out ? io_r_739_b : _GEN_6078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6080 = 10'h2e4 == r_count_7_io_out ? io_r_740_b : _GEN_6079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6081 = 10'h2e5 == r_count_7_io_out ? io_r_741_b : _GEN_6080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6082 = 10'h2e6 == r_count_7_io_out ? io_r_742_b : _GEN_6081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6083 = 10'h2e7 == r_count_7_io_out ? io_r_743_b : _GEN_6082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6084 = 10'h2e8 == r_count_7_io_out ? io_r_744_b : _GEN_6083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6085 = 10'h2e9 == r_count_7_io_out ? io_r_745_b : _GEN_6084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6086 = 10'h2ea == r_count_7_io_out ? io_r_746_b : _GEN_6085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6087 = 10'h2eb == r_count_7_io_out ? io_r_747_b : _GEN_6086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6088 = 10'h2ec == r_count_7_io_out ? io_r_748_b : _GEN_6087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6091 = 10'h1 == r_count_8_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6092 = 10'h2 == r_count_8_io_out ? io_r_2_b : _GEN_6091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6093 = 10'h3 == r_count_8_io_out ? io_r_3_b : _GEN_6092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6094 = 10'h4 == r_count_8_io_out ? io_r_4_b : _GEN_6093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6095 = 10'h5 == r_count_8_io_out ? io_r_5_b : _GEN_6094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6096 = 10'h6 == r_count_8_io_out ? io_r_6_b : _GEN_6095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6097 = 10'h7 == r_count_8_io_out ? io_r_7_b : _GEN_6096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6098 = 10'h8 == r_count_8_io_out ? io_r_8_b : _GEN_6097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6099 = 10'h9 == r_count_8_io_out ? io_r_9_b : _GEN_6098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6100 = 10'ha == r_count_8_io_out ? io_r_10_b : _GEN_6099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6101 = 10'hb == r_count_8_io_out ? io_r_11_b : _GEN_6100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6102 = 10'hc == r_count_8_io_out ? io_r_12_b : _GEN_6101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6103 = 10'hd == r_count_8_io_out ? io_r_13_b : _GEN_6102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6104 = 10'he == r_count_8_io_out ? io_r_14_b : _GEN_6103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6105 = 10'hf == r_count_8_io_out ? io_r_15_b : _GEN_6104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6106 = 10'h10 == r_count_8_io_out ? io_r_16_b : _GEN_6105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6107 = 10'h11 == r_count_8_io_out ? io_r_17_b : _GEN_6106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6108 = 10'h12 == r_count_8_io_out ? io_r_18_b : _GEN_6107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6109 = 10'h13 == r_count_8_io_out ? io_r_19_b : _GEN_6108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6110 = 10'h14 == r_count_8_io_out ? io_r_20_b : _GEN_6109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6111 = 10'h15 == r_count_8_io_out ? io_r_21_b : _GEN_6110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6112 = 10'h16 == r_count_8_io_out ? io_r_22_b : _GEN_6111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6113 = 10'h17 == r_count_8_io_out ? io_r_23_b : _GEN_6112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6114 = 10'h18 == r_count_8_io_out ? io_r_24_b : _GEN_6113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6115 = 10'h19 == r_count_8_io_out ? io_r_25_b : _GEN_6114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6116 = 10'h1a == r_count_8_io_out ? io_r_26_b : _GEN_6115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6117 = 10'h1b == r_count_8_io_out ? io_r_27_b : _GEN_6116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6118 = 10'h1c == r_count_8_io_out ? io_r_28_b : _GEN_6117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6119 = 10'h1d == r_count_8_io_out ? io_r_29_b : _GEN_6118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6120 = 10'h1e == r_count_8_io_out ? io_r_30_b : _GEN_6119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6121 = 10'h1f == r_count_8_io_out ? io_r_31_b : _GEN_6120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6122 = 10'h20 == r_count_8_io_out ? io_r_32_b : _GEN_6121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6123 = 10'h21 == r_count_8_io_out ? io_r_33_b : _GEN_6122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6124 = 10'h22 == r_count_8_io_out ? io_r_34_b : _GEN_6123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6125 = 10'h23 == r_count_8_io_out ? io_r_35_b : _GEN_6124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6126 = 10'h24 == r_count_8_io_out ? io_r_36_b : _GEN_6125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6127 = 10'h25 == r_count_8_io_out ? io_r_37_b : _GEN_6126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6128 = 10'h26 == r_count_8_io_out ? io_r_38_b : _GEN_6127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6129 = 10'h27 == r_count_8_io_out ? io_r_39_b : _GEN_6128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6130 = 10'h28 == r_count_8_io_out ? io_r_40_b : _GEN_6129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6131 = 10'h29 == r_count_8_io_out ? io_r_41_b : _GEN_6130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6132 = 10'h2a == r_count_8_io_out ? io_r_42_b : _GEN_6131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6133 = 10'h2b == r_count_8_io_out ? io_r_43_b : _GEN_6132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6134 = 10'h2c == r_count_8_io_out ? io_r_44_b : _GEN_6133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6135 = 10'h2d == r_count_8_io_out ? io_r_45_b : _GEN_6134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6136 = 10'h2e == r_count_8_io_out ? io_r_46_b : _GEN_6135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6137 = 10'h2f == r_count_8_io_out ? io_r_47_b : _GEN_6136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6138 = 10'h30 == r_count_8_io_out ? io_r_48_b : _GEN_6137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6139 = 10'h31 == r_count_8_io_out ? io_r_49_b : _GEN_6138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6140 = 10'h32 == r_count_8_io_out ? io_r_50_b : _GEN_6139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6141 = 10'h33 == r_count_8_io_out ? io_r_51_b : _GEN_6140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6142 = 10'h34 == r_count_8_io_out ? io_r_52_b : _GEN_6141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6143 = 10'h35 == r_count_8_io_out ? io_r_53_b : _GEN_6142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6144 = 10'h36 == r_count_8_io_out ? io_r_54_b : _GEN_6143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6145 = 10'h37 == r_count_8_io_out ? io_r_55_b : _GEN_6144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6146 = 10'h38 == r_count_8_io_out ? io_r_56_b : _GEN_6145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6147 = 10'h39 == r_count_8_io_out ? io_r_57_b : _GEN_6146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6148 = 10'h3a == r_count_8_io_out ? io_r_58_b : _GEN_6147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6149 = 10'h3b == r_count_8_io_out ? io_r_59_b : _GEN_6148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6150 = 10'h3c == r_count_8_io_out ? io_r_60_b : _GEN_6149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6151 = 10'h3d == r_count_8_io_out ? io_r_61_b : _GEN_6150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6152 = 10'h3e == r_count_8_io_out ? io_r_62_b : _GEN_6151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6153 = 10'h3f == r_count_8_io_out ? io_r_63_b : _GEN_6152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6154 = 10'h40 == r_count_8_io_out ? io_r_64_b : _GEN_6153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6155 = 10'h41 == r_count_8_io_out ? io_r_65_b : _GEN_6154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6156 = 10'h42 == r_count_8_io_out ? io_r_66_b : _GEN_6155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6157 = 10'h43 == r_count_8_io_out ? io_r_67_b : _GEN_6156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6158 = 10'h44 == r_count_8_io_out ? io_r_68_b : _GEN_6157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6159 = 10'h45 == r_count_8_io_out ? io_r_69_b : _GEN_6158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6160 = 10'h46 == r_count_8_io_out ? io_r_70_b : _GEN_6159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6161 = 10'h47 == r_count_8_io_out ? io_r_71_b : _GEN_6160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6162 = 10'h48 == r_count_8_io_out ? io_r_72_b : _GEN_6161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6163 = 10'h49 == r_count_8_io_out ? io_r_73_b : _GEN_6162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6164 = 10'h4a == r_count_8_io_out ? io_r_74_b : _GEN_6163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6165 = 10'h4b == r_count_8_io_out ? io_r_75_b : _GEN_6164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6166 = 10'h4c == r_count_8_io_out ? io_r_76_b : _GEN_6165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6167 = 10'h4d == r_count_8_io_out ? io_r_77_b : _GEN_6166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6168 = 10'h4e == r_count_8_io_out ? io_r_78_b : _GEN_6167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6169 = 10'h4f == r_count_8_io_out ? io_r_79_b : _GEN_6168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6170 = 10'h50 == r_count_8_io_out ? io_r_80_b : _GEN_6169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6171 = 10'h51 == r_count_8_io_out ? io_r_81_b : _GEN_6170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6172 = 10'h52 == r_count_8_io_out ? io_r_82_b : _GEN_6171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6173 = 10'h53 == r_count_8_io_out ? io_r_83_b : _GEN_6172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6174 = 10'h54 == r_count_8_io_out ? io_r_84_b : _GEN_6173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6175 = 10'h55 == r_count_8_io_out ? io_r_85_b : _GEN_6174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6176 = 10'h56 == r_count_8_io_out ? io_r_86_b : _GEN_6175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6177 = 10'h57 == r_count_8_io_out ? io_r_87_b : _GEN_6176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6178 = 10'h58 == r_count_8_io_out ? io_r_88_b : _GEN_6177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6179 = 10'h59 == r_count_8_io_out ? io_r_89_b : _GEN_6178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6180 = 10'h5a == r_count_8_io_out ? io_r_90_b : _GEN_6179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6181 = 10'h5b == r_count_8_io_out ? io_r_91_b : _GEN_6180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6182 = 10'h5c == r_count_8_io_out ? io_r_92_b : _GEN_6181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6183 = 10'h5d == r_count_8_io_out ? io_r_93_b : _GEN_6182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6184 = 10'h5e == r_count_8_io_out ? io_r_94_b : _GEN_6183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6185 = 10'h5f == r_count_8_io_out ? io_r_95_b : _GEN_6184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6186 = 10'h60 == r_count_8_io_out ? io_r_96_b : _GEN_6185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6187 = 10'h61 == r_count_8_io_out ? io_r_97_b : _GEN_6186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6188 = 10'h62 == r_count_8_io_out ? io_r_98_b : _GEN_6187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6189 = 10'h63 == r_count_8_io_out ? io_r_99_b : _GEN_6188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6190 = 10'h64 == r_count_8_io_out ? io_r_100_b : _GEN_6189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6191 = 10'h65 == r_count_8_io_out ? io_r_101_b : _GEN_6190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6192 = 10'h66 == r_count_8_io_out ? io_r_102_b : _GEN_6191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6193 = 10'h67 == r_count_8_io_out ? io_r_103_b : _GEN_6192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6194 = 10'h68 == r_count_8_io_out ? io_r_104_b : _GEN_6193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6195 = 10'h69 == r_count_8_io_out ? io_r_105_b : _GEN_6194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6196 = 10'h6a == r_count_8_io_out ? io_r_106_b : _GEN_6195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6197 = 10'h6b == r_count_8_io_out ? io_r_107_b : _GEN_6196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6198 = 10'h6c == r_count_8_io_out ? io_r_108_b : _GEN_6197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6199 = 10'h6d == r_count_8_io_out ? io_r_109_b : _GEN_6198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6200 = 10'h6e == r_count_8_io_out ? io_r_110_b : _GEN_6199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6201 = 10'h6f == r_count_8_io_out ? io_r_111_b : _GEN_6200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6202 = 10'h70 == r_count_8_io_out ? io_r_112_b : _GEN_6201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6203 = 10'h71 == r_count_8_io_out ? io_r_113_b : _GEN_6202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6204 = 10'h72 == r_count_8_io_out ? io_r_114_b : _GEN_6203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6205 = 10'h73 == r_count_8_io_out ? io_r_115_b : _GEN_6204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6206 = 10'h74 == r_count_8_io_out ? io_r_116_b : _GEN_6205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6207 = 10'h75 == r_count_8_io_out ? io_r_117_b : _GEN_6206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6208 = 10'h76 == r_count_8_io_out ? io_r_118_b : _GEN_6207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6209 = 10'h77 == r_count_8_io_out ? io_r_119_b : _GEN_6208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6210 = 10'h78 == r_count_8_io_out ? io_r_120_b : _GEN_6209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6211 = 10'h79 == r_count_8_io_out ? io_r_121_b : _GEN_6210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6212 = 10'h7a == r_count_8_io_out ? io_r_122_b : _GEN_6211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6213 = 10'h7b == r_count_8_io_out ? io_r_123_b : _GEN_6212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6214 = 10'h7c == r_count_8_io_out ? io_r_124_b : _GEN_6213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6215 = 10'h7d == r_count_8_io_out ? io_r_125_b : _GEN_6214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6216 = 10'h7e == r_count_8_io_out ? io_r_126_b : _GEN_6215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6217 = 10'h7f == r_count_8_io_out ? io_r_127_b : _GEN_6216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6218 = 10'h80 == r_count_8_io_out ? io_r_128_b : _GEN_6217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6219 = 10'h81 == r_count_8_io_out ? io_r_129_b : _GEN_6218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6220 = 10'h82 == r_count_8_io_out ? io_r_130_b : _GEN_6219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6221 = 10'h83 == r_count_8_io_out ? io_r_131_b : _GEN_6220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6222 = 10'h84 == r_count_8_io_out ? io_r_132_b : _GEN_6221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6223 = 10'h85 == r_count_8_io_out ? io_r_133_b : _GEN_6222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6224 = 10'h86 == r_count_8_io_out ? io_r_134_b : _GEN_6223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6225 = 10'h87 == r_count_8_io_out ? io_r_135_b : _GEN_6224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6226 = 10'h88 == r_count_8_io_out ? io_r_136_b : _GEN_6225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6227 = 10'h89 == r_count_8_io_out ? io_r_137_b : _GEN_6226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6228 = 10'h8a == r_count_8_io_out ? io_r_138_b : _GEN_6227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6229 = 10'h8b == r_count_8_io_out ? io_r_139_b : _GEN_6228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6230 = 10'h8c == r_count_8_io_out ? io_r_140_b : _GEN_6229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6231 = 10'h8d == r_count_8_io_out ? io_r_141_b : _GEN_6230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6232 = 10'h8e == r_count_8_io_out ? io_r_142_b : _GEN_6231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6233 = 10'h8f == r_count_8_io_out ? io_r_143_b : _GEN_6232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6234 = 10'h90 == r_count_8_io_out ? io_r_144_b : _GEN_6233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6235 = 10'h91 == r_count_8_io_out ? io_r_145_b : _GEN_6234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6236 = 10'h92 == r_count_8_io_out ? io_r_146_b : _GEN_6235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6237 = 10'h93 == r_count_8_io_out ? io_r_147_b : _GEN_6236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6238 = 10'h94 == r_count_8_io_out ? io_r_148_b : _GEN_6237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6239 = 10'h95 == r_count_8_io_out ? io_r_149_b : _GEN_6238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6240 = 10'h96 == r_count_8_io_out ? io_r_150_b : _GEN_6239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6241 = 10'h97 == r_count_8_io_out ? io_r_151_b : _GEN_6240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6242 = 10'h98 == r_count_8_io_out ? io_r_152_b : _GEN_6241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6243 = 10'h99 == r_count_8_io_out ? io_r_153_b : _GEN_6242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6244 = 10'h9a == r_count_8_io_out ? io_r_154_b : _GEN_6243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6245 = 10'h9b == r_count_8_io_out ? io_r_155_b : _GEN_6244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6246 = 10'h9c == r_count_8_io_out ? io_r_156_b : _GEN_6245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6247 = 10'h9d == r_count_8_io_out ? io_r_157_b : _GEN_6246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6248 = 10'h9e == r_count_8_io_out ? io_r_158_b : _GEN_6247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6249 = 10'h9f == r_count_8_io_out ? io_r_159_b : _GEN_6248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6250 = 10'ha0 == r_count_8_io_out ? io_r_160_b : _GEN_6249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6251 = 10'ha1 == r_count_8_io_out ? io_r_161_b : _GEN_6250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6252 = 10'ha2 == r_count_8_io_out ? io_r_162_b : _GEN_6251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6253 = 10'ha3 == r_count_8_io_out ? io_r_163_b : _GEN_6252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6254 = 10'ha4 == r_count_8_io_out ? io_r_164_b : _GEN_6253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6255 = 10'ha5 == r_count_8_io_out ? io_r_165_b : _GEN_6254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6256 = 10'ha6 == r_count_8_io_out ? io_r_166_b : _GEN_6255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6257 = 10'ha7 == r_count_8_io_out ? io_r_167_b : _GEN_6256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6258 = 10'ha8 == r_count_8_io_out ? io_r_168_b : _GEN_6257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6259 = 10'ha9 == r_count_8_io_out ? io_r_169_b : _GEN_6258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6260 = 10'haa == r_count_8_io_out ? io_r_170_b : _GEN_6259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6261 = 10'hab == r_count_8_io_out ? io_r_171_b : _GEN_6260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6262 = 10'hac == r_count_8_io_out ? io_r_172_b : _GEN_6261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6263 = 10'had == r_count_8_io_out ? io_r_173_b : _GEN_6262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6264 = 10'hae == r_count_8_io_out ? io_r_174_b : _GEN_6263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6265 = 10'haf == r_count_8_io_out ? io_r_175_b : _GEN_6264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6266 = 10'hb0 == r_count_8_io_out ? io_r_176_b : _GEN_6265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6267 = 10'hb1 == r_count_8_io_out ? io_r_177_b : _GEN_6266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6268 = 10'hb2 == r_count_8_io_out ? io_r_178_b : _GEN_6267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6269 = 10'hb3 == r_count_8_io_out ? io_r_179_b : _GEN_6268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6270 = 10'hb4 == r_count_8_io_out ? io_r_180_b : _GEN_6269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6271 = 10'hb5 == r_count_8_io_out ? io_r_181_b : _GEN_6270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6272 = 10'hb6 == r_count_8_io_out ? io_r_182_b : _GEN_6271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6273 = 10'hb7 == r_count_8_io_out ? io_r_183_b : _GEN_6272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6274 = 10'hb8 == r_count_8_io_out ? io_r_184_b : _GEN_6273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6275 = 10'hb9 == r_count_8_io_out ? io_r_185_b : _GEN_6274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6276 = 10'hba == r_count_8_io_out ? io_r_186_b : _GEN_6275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6277 = 10'hbb == r_count_8_io_out ? io_r_187_b : _GEN_6276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6278 = 10'hbc == r_count_8_io_out ? io_r_188_b : _GEN_6277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6279 = 10'hbd == r_count_8_io_out ? io_r_189_b : _GEN_6278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6280 = 10'hbe == r_count_8_io_out ? io_r_190_b : _GEN_6279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6281 = 10'hbf == r_count_8_io_out ? io_r_191_b : _GEN_6280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6282 = 10'hc0 == r_count_8_io_out ? io_r_192_b : _GEN_6281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6283 = 10'hc1 == r_count_8_io_out ? io_r_193_b : _GEN_6282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6284 = 10'hc2 == r_count_8_io_out ? io_r_194_b : _GEN_6283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6285 = 10'hc3 == r_count_8_io_out ? io_r_195_b : _GEN_6284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6286 = 10'hc4 == r_count_8_io_out ? io_r_196_b : _GEN_6285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6287 = 10'hc5 == r_count_8_io_out ? io_r_197_b : _GEN_6286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6288 = 10'hc6 == r_count_8_io_out ? io_r_198_b : _GEN_6287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6289 = 10'hc7 == r_count_8_io_out ? io_r_199_b : _GEN_6288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6290 = 10'hc8 == r_count_8_io_out ? io_r_200_b : _GEN_6289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6291 = 10'hc9 == r_count_8_io_out ? io_r_201_b : _GEN_6290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6292 = 10'hca == r_count_8_io_out ? io_r_202_b : _GEN_6291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6293 = 10'hcb == r_count_8_io_out ? io_r_203_b : _GEN_6292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6294 = 10'hcc == r_count_8_io_out ? io_r_204_b : _GEN_6293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6295 = 10'hcd == r_count_8_io_out ? io_r_205_b : _GEN_6294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6296 = 10'hce == r_count_8_io_out ? io_r_206_b : _GEN_6295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6297 = 10'hcf == r_count_8_io_out ? io_r_207_b : _GEN_6296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6298 = 10'hd0 == r_count_8_io_out ? io_r_208_b : _GEN_6297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6299 = 10'hd1 == r_count_8_io_out ? io_r_209_b : _GEN_6298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6300 = 10'hd2 == r_count_8_io_out ? io_r_210_b : _GEN_6299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6301 = 10'hd3 == r_count_8_io_out ? io_r_211_b : _GEN_6300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6302 = 10'hd4 == r_count_8_io_out ? io_r_212_b : _GEN_6301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6303 = 10'hd5 == r_count_8_io_out ? io_r_213_b : _GEN_6302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6304 = 10'hd6 == r_count_8_io_out ? io_r_214_b : _GEN_6303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6305 = 10'hd7 == r_count_8_io_out ? io_r_215_b : _GEN_6304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6306 = 10'hd8 == r_count_8_io_out ? io_r_216_b : _GEN_6305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6307 = 10'hd9 == r_count_8_io_out ? io_r_217_b : _GEN_6306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6308 = 10'hda == r_count_8_io_out ? io_r_218_b : _GEN_6307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6309 = 10'hdb == r_count_8_io_out ? io_r_219_b : _GEN_6308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6310 = 10'hdc == r_count_8_io_out ? io_r_220_b : _GEN_6309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6311 = 10'hdd == r_count_8_io_out ? io_r_221_b : _GEN_6310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6312 = 10'hde == r_count_8_io_out ? io_r_222_b : _GEN_6311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6313 = 10'hdf == r_count_8_io_out ? io_r_223_b : _GEN_6312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6314 = 10'he0 == r_count_8_io_out ? io_r_224_b : _GEN_6313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6315 = 10'he1 == r_count_8_io_out ? io_r_225_b : _GEN_6314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6316 = 10'he2 == r_count_8_io_out ? io_r_226_b : _GEN_6315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6317 = 10'he3 == r_count_8_io_out ? io_r_227_b : _GEN_6316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6318 = 10'he4 == r_count_8_io_out ? io_r_228_b : _GEN_6317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6319 = 10'he5 == r_count_8_io_out ? io_r_229_b : _GEN_6318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6320 = 10'he6 == r_count_8_io_out ? io_r_230_b : _GEN_6319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6321 = 10'he7 == r_count_8_io_out ? io_r_231_b : _GEN_6320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6322 = 10'he8 == r_count_8_io_out ? io_r_232_b : _GEN_6321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6323 = 10'he9 == r_count_8_io_out ? io_r_233_b : _GEN_6322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6324 = 10'hea == r_count_8_io_out ? io_r_234_b : _GEN_6323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6325 = 10'heb == r_count_8_io_out ? io_r_235_b : _GEN_6324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6326 = 10'hec == r_count_8_io_out ? io_r_236_b : _GEN_6325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6327 = 10'hed == r_count_8_io_out ? io_r_237_b : _GEN_6326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6328 = 10'hee == r_count_8_io_out ? io_r_238_b : _GEN_6327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6329 = 10'hef == r_count_8_io_out ? io_r_239_b : _GEN_6328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6330 = 10'hf0 == r_count_8_io_out ? io_r_240_b : _GEN_6329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6331 = 10'hf1 == r_count_8_io_out ? io_r_241_b : _GEN_6330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6332 = 10'hf2 == r_count_8_io_out ? io_r_242_b : _GEN_6331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6333 = 10'hf3 == r_count_8_io_out ? io_r_243_b : _GEN_6332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6334 = 10'hf4 == r_count_8_io_out ? io_r_244_b : _GEN_6333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6335 = 10'hf5 == r_count_8_io_out ? io_r_245_b : _GEN_6334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6336 = 10'hf6 == r_count_8_io_out ? io_r_246_b : _GEN_6335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6337 = 10'hf7 == r_count_8_io_out ? io_r_247_b : _GEN_6336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6338 = 10'hf8 == r_count_8_io_out ? io_r_248_b : _GEN_6337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6339 = 10'hf9 == r_count_8_io_out ? io_r_249_b : _GEN_6338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6340 = 10'hfa == r_count_8_io_out ? io_r_250_b : _GEN_6339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6341 = 10'hfb == r_count_8_io_out ? io_r_251_b : _GEN_6340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6342 = 10'hfc == r_count_8_io_out ? io_r_252_b : _GEN_6341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6343 = 10'hfd == r_count_8_io_out ? io_r_253_b : _GEN_6342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6344 = 10'hfe == r_count_8_io_out ? io_r_254_b : _GEN_6343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6345 = 10'hff == r_count_8_io_out ? io_r_255_b : _GEN_6344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6346 = 10'h100 == r_count_8_io_out ? io_r_256_b : _GEN_6345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6347 = 10'h101 == r_count_8_io_out ? io_r_257_b : _GEN_6346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6348 = 10'h102 == r_count_8_io_out ? io_r_258_b : _GEN_6347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6349 = 10'h103 == r_count_8_io_out ? io_r_259_b : _GEN_6348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6350 = 10'h104 == r_count_8_io_out ? io_r_260_b : _GEN_6349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6351 = 10'h105 == r_count_8_io_out ? io_r_261_b : _GEN_6350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6352 = 10'h106 == r_count_8_io_out ? io_r_262_b : _GEN_6351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6353 = 10'h107 == r_count_8_io_out ? io_r_263_b : _GEN_6352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6354 = 10'h108 == r_count_8_io_out ? io_r_264_b : _GEN_6353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6355 = 10'h109 == r_count_8_io_out ? io_r_265_b : _GEN_6354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6356 = 10'h10a == r_count_8_io_out ? io_r_266_b : _GEN_6355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6357 = 10'h10b == r_count_8_io_out ? io_r_267_b : _GEN_6356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6358 = 10'h10c == r_count_8_io_out ? io_r_268_b : _GEN_6357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6359 = 10'h10d == r_count_8_io_out ? io_r_269_b : _GEN_6358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6360 = 10'h10e == r_count_8_io_out ? io_r_270_b : _GEN_6359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6361 = 10'h10f == r_count_8_io_out ? io_r_271_b : _GEN_6360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6362 = 10'h110 == r_count_8_io_out ? io_r_272_b : _GEN_6361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6363 = 10'h111 == r_count_8_io_out ? io_r_273_b : _GEN_6362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6364 = 10'h112 == r_count_8_io_out ? io_r_274_b : _GEN_6363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6365 = 10'h113 == r_count_8_io_out ? io_r_275_b : _GEN_6364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6366 = 10'h114 == r_count_8_io_out ? io_r_276_b : _GEN_6365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6367 = 10'h115 == r_count_8_io_out ? io_r_277_b : _GEN_6366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6368 = 10'h116 == r_count_8_io_out ? io_r_278_b : _GEN_6367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6369 = 10'h117 == r_count_8_io_out ? io_r_279_b : _GEN_6368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6370 = 10'h118 == r_count_8_io_out ? io_r_280_b : _GEN_6369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6371 = 10'h119 == r_count_8_io_out ? io_r_281_b : _GEN_6370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6372 = 10'h11a == r_count_8_io_out ? io_r_282_b : _GEN_6371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6373 = 10'h11b == r_count_8_io_out ? io_r_283_b : _GEN_6372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6374 = 10'h11c == r_count_8_io_out ? io_r_284_b : _GEN_6373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6375 = 10'h11d == r_count_8_io_out ? io_r_285_b : _GEN_6374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6376 = 10'h11e == r_count_8_io_out ? io_r_286_b : _GEN_6375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6377 = 10'h11f == r_count_8_io_out ? io_r_287_b : _GEN_6376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6378 = 10'h120 == r_count_8_io_out ? io_r_288_b : _GEN_6377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6379 = 10'h121 == r_count_8_io_out ? io_r_289_b : _GEN_6378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6380 = 10'h122 == r_count_8_io_out ? io_r_290_b : _GEN_6379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6381 = 10'h123 == r_count_8_io_out ? io_r_291_b : _GEN_6380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6382 = 10'h124 == r_count_8_io_out ? io_r_292_b : _GEN_6381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6383 = 10'h125 == r_count_8_io_out ? io_r_293_b : _GEN_6382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6384 = 10'h126 == r_count_8_io_out ? io_r_294_b : _GEN_6383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6385 = 10'h127 == r_count_8_io_out ? io_r_295_b : _GEN_6384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6386 = 10'h128 == r_count_8_io_out ? io_r_296_b : _GEN_6385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6387 = 10'h129 == r_count_8_io_out ? io_r_297_b : _GEN_6386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6388 = 10'h12a == r_count_8_io_out ? io_r_298_b : _GEN_6387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6389 = 10'h12b == r_count_8_io_out ? io_r_299_b : _GEN_6388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6390 = 10'h12c == r_count_8_io_out ? io_r_300_b : _GEN_6389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6391 = 10'h12d == r_count_8_io_out ? io_r_301_b : _GEN_6390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6392 = 10'h12e == r_count_8_io_out ? io_r_302_b : _GEN_6391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6393 = 10'h12f == r_count_8_io_out ? io_r_303_b : _GEN_6392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6394 = 10'h130 == r_count_8_io_out ? io_r_304_b : _GEN_6393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6395 = 10'h131 == r_count_8_io_out ? io_r_305_b : _GEN_6394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6396 = 10'h132 == r_count_8_io_out ? io_r_306_b : _GEN_6395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6397 = 10'h133 == r_count_8_io_out ? io_r_307_b : _GEN_6396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6398 = 10'h134 == r_count_8_io_out ? io_r_308_b : _GEN_6397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6399 = 10'h135 == r_count_8_io_out ? io_r_309_b : _GEN_6398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6400 = 10'h136 == r_count_8_io_out ? io_r_310_b : _GEN_6399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6401 = 10'h137 == r_count_8_io_out ? io_r_311_b : _GEN_6400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6402 = 10'h138 == r_count_8_io_out ? io_r_312_b : _GEN_6401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6403 = 10'h139 == r_count_8_io_out ? io_r_313_b : _GEN_6402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6404 = 10'h13a == r_count_8_io_out ? io_r_314_b : _GEN_6403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6405 = 10'h13b == r_count_8_io_out ? io_r_315_b : _GEN_6404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6406 = 10'h13c == r_count_8_io_out ? io_r_316_b : _GEN_6405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6407 = 10'h13d == r_count_8_io_out ? io_r_317_b : _GEN_6406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6408 = 10'h13e == r_count_8_io_out ? io_r_318_b : _GEN_6407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6409 = 10'h13f == r_count_8_io_out ? io_r_319_b : _GEN_6408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6410 = 10'h140 == r_count_8_io_out ? io_r_320_b : _GEN_6409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6411 = 10'h141 == r_count_8_io_out ? io_r_321_b : _GEN_6410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6412 = 10'h142 == r_count_8_io_out ? io_r_322_b : _GEN_6411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6413 = 10'h143 == r_count_8_io_out ? io_r_323_b : _GEN_6412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6414 = 10'h144 == r_count_8_io_out ? io_r_324_b : _GEN_6413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6415 = 10'h145 == r_count_8_io_out ? io_r_325_b : _GEN_6414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6416 = 10'h146 == r_count_8_io_out ? io_r_326_b : _GEN_6415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6417 = 10'h147 == r_count_8_io_out ? io_r_327_b : _GEN_6416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6418 = 10'h148 == r_count_8_io_out ? io_r_328_b : _GEN_6417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6419 = 10'h149 == r_count_8_io_out ? io_r_329_b : _GEN_6418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6420 = 10'h14a == r_count_8_io_out ? io_r_330_b : _GEN_6419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6421 = 10'h14b == r_count_8_io_out ? io_r_331_b : _GEN_6420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6422 = 10'h14c == r_count_8_io_out ? io_r_332_b : _GEN_6421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6423 = 10'h14d == r_count_8_io_out ? io_r_333_b : _GEN_6422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6424 = 10'h14e == r_count_8_io_out ? io_r_334_b : _GEN_6423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6425 = 10'h14f == r_count_8_io_out ? io_r_335_b : _GEN_6424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6426 = 10'h150 == r_count_8_io_out ? io_r_336_b : _GEN_6425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6427 = 10'h151 == r_count_8_io_out ? io_r_337_b : _GEN_6426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6428 = 10'h152 == r_count_8_io_out ? io_r_338_b : _GEN_6427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6429 = 10'h153 == r_count_8_io_out ? io_r_339_b : _GEN_6428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6430 = 10'h154 == r_count_8_io_out ? io_r_340_b : _GEN_6429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6431 = 10'h155 == r_count_8_io_out ? io_r_341_b : _GEN_6430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6432 = 10'h156 == r_count_8_io_out ? io_r_342_b : _GEN_6431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6433 = 10'h157 == r_count_8_io_out ? io_r_343_b : _GEN_6432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6434 = 10'h158 == r_count_8_io_out ? io_r_344_b : _GEN_6433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6435 = 10'h159 == r_count_8_io_out ? io_r_345_b : _GEN_6434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6436 = 10'h15a == r_count_8_io_out ? io_r_346_b : _GEN_6435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6437 = 10'h15b == r_count_8_io_out ? io_r_347_b : _GEN_6436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6438 = 10'h15c == r_count_8_io_out ? io_r_348_b : _GEN_6437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6439 = 10'h15d == r_count_8_io_out ? io_r_349_b : _GEN_6438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6440 = 10'h15e == r_count_8_io_out ? io_r_350_b : _GEN_6439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6441 = 10'h15f == r_count_8_io_out ? io_r_351_b : _GEN_6440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6442 = 10'h160 == r_count_8_io_out ? io_r_352_b : _GEN_6441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6443 = 10'h161 == r_count_8_io_out ? io_r_353_b : _GEN_6442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6444 = 10'h162 == r_count_8_io_out ? io_r_354_b : _GEN_6443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6445 = 10'h163 == r_count_8_io_out ? io_r_355_b : _GEN_6444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6446 = 10'h164 == r_count_8_io_out ? io_r_356_b : _GEN_6445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6447 = 10'h165 == r_count_8_io_out ? io_r_357_b : _GEN_6446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6448 = 10'h166 == r_count_8_io_out ? io_r_358_b : _GEN_6447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6449 = 10'h167 == r_count_8_io_out ? io_r_359_b : _GEN_6448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6450 = 10'h168 == r_count_8_io_out ? io_r_360_b : _GEN_6449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6451 = 10'h169 == r_count_8_io_out ? io_r_361_b : _GEN_6450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6452 = 10'h16a == r_count_8_io_out ? io_r_362_b : _GEN_6451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6453 = 10'h16b == r_count_8_io_out ? io_r_363_b : _GEN_6452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6454 = 10'h16c == r_count_8_io_out ? io_r_364_b : _GEN_6453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6455 = 10'h16d == r_count_8_io_out ? io_r_365_b : _GEN_6454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6456 = 10'h16e == r_count_8_io_out ? io_r_366_b : _GEN_6455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6457 = 10'h16f == r_count_8_io_out ? io_r_367_b : _GEN_6456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6458 = 10'h170 == r_count_8_io_out ? io_r_368_b : _GEN_6457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6459 = 10'h171 == r_count_8_io_out ? io_r_369_b : _GEN_6458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6460 = 10'h172 == r_count_8_io_out ? io_r_370_b : _GEN_6459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6461 = 10'h173 == r_count_8_io_out ? io_r_371_b : _GEN_6460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6462 = 10'h174 == r_count_8_io_out ? io_r_372_b : _GEN_6461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6463 = 10'h175 == r_count_8_io_out ? io_r_373_b : _GEN_6462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6464 = 10'h176 == r_count_8_io_out ? io_r_374_b : _GEN_6463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6465 = 10'h177 == r_count_8_io_out ? io_r_375_b : _GEN_6464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6466 = 10'h178 == r_count_8_io_out ? io_r_376_b : _GEN_6465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6467 = 10'h179 == r_count_8_io_out ? io_r_377_b : _GEN_6466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6468 = 10'h17a == r_count_8_io_out ? io_r_378_b : _GEN_6467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6469 = 10'h17b == r_count_8_io_out ? io_r_379_b : _GEN_6468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6470 = 10'h17c == r_count_8_io_out ? io_r_380_b : _GEN_6469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6471 = 10'h17d == r_count_8_io_out ? io_r_381_b : _GEN_6470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6472 = 10'h17e == r_count_8_io_out ? io_r_382_b : _GEN_6471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6473 = 10'h17f == r_count_8_io_out ? io_r_383_b : _GEN_6472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6474 = 10'h180 == r_count_8_io_out ? io_r_384_b : _GEN_6473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6475 = 10'h181 == r_count_8_io_out ? io_r_385_b : _GEN_6474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6476 = 10'h182 == r_count_8_io_out ? io_r_386_b : _GEN_6475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6477 = 10'h183 == r_count_8_io_out ? io_r_387_b : _GEN_6476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6478 = 10'h184 == r_count_8_io_out ? io_r_388_b : _GEN_6477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6479 = 10'h185 == r_count_8_io_out ? io_r_389_b : _GEN_6478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6480 = 10'h186 == r_count_8_io_out ? io_r_390_b : _GEN_6479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6481 = 10'h187 == r_count_8_io_out ? io_r_391_b : _GEN_6480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6482 = 10'h188 == r_count_8_io_out ? io_r_392_b : _GEN_6481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6483 = 10'h189 == r_count_8_io_out ? io_r_393_b : _GEN_6482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6484 = 10'h18a == r_count_8_io_out ? io_r_394_b : _GEN_6483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6485 = 10'h18b == r_count_8_io_out ? io_r_395_b : _GEN_6484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6486 = 10'h18c == r_count_8_io_out ? io_r_396_b : _GEN_6485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6487 = 10'h18d == r_count_8_io_out ? io_r_397_b : _GEN_6486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6488 = 10'h18e == r_count_8_io_out ? io_r_398_b : _GEN_6487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6489 = 10'h18f == r_count_8_io_out ? io_r_399_b : _GEN_6488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6490 = 10'h190 == r_count_8_io_out ? io_r_400_b : _GEN_6489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6491 = 10'h191 == r_count_8_io_out ? io_r_401_b : _GEN_6490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6492 = 10'h192 == r_count_8_io_out ? io_r_402_b : _GEN_6491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6493 = 10'h193 == r_count_8_io_out ? io_r_403_b : _GEN_6492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6494 = 10'h194 == r_count_8_io_out ? io_r_404_b : _GEN_6493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6495 = 10'h195 == r_count_8_io_out ? io_r_405_b : _GEN_6494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6496 = 10'h196 == r_count_8_io_out ? io_r_406_b : _GEN_6495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6497 = 10'h197 == r_count_8_io_out ? io_r_407_b : _GEN_6496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6498 = 10'h198 == r_count_8_io_out ? io_r_408_b : _GEN_6497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6499 = 10'h199 == r_count_8_io_out ? io_r_409_b : _GEN_6498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6500 = 10'h19a == r_count_8_io_out ? io_r_410_b : _GEN_6499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6501 = 10'h19b == r_count_8_io_out ? io_r_411_b : _GEN_6500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6502 = 10'h19c == r_count_8_io_out ? io_r_412_b : _GEN_6501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6503 = 10'h19d == r_count_8_io_out ? io_r_413_b : _GEN_6502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6504 = 10'h19e == r_count_8_io_out ? io_r_414_b : _GEN_6503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6505 = 10'h19f == r_count_8_io_out ? io_r_415_b : _GEN_6504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6506 = 10'h1a0 == r_count_8_io_out ? io_r_416_b : _GEN_6505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6507 = 10'h1a1 == r_count_8_io_out ? io_r_417_b : _GEN_6506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6508 = 10'h1a2 == r_count_8_io_out ? io_r_418_b : _GEN_6507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6509 = 10'h1a3 == r_count_8_io_out ? io_r_419_b : _GEN_6508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6510 = 10'h1a4 == r_count_8_io_out ? io_r_420_b : _GEN_6509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6511 = 10'h1a5 == r_count_8_io_out ? io_r_421_b : _GEN_6510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6512 = 10'h1a6 == r_count_8_io_out ? io_r_422_b : _GEN_6511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6513 = 10'h1a7 == r_count_8_io_out ? io_r_423_b : _GEN_6512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6514 = 10'h1a8 == r_count_8_io_out ? io_r_424_b : _GEN_6513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6515 = 10'h1a9 == r_count_8_io_out ? io_r_425_b : _GEN_6514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6516 = 10'h1aa == r_count_8_io_out ? io_r_426_b : _GEN_6515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6517 = 10'h1ab == r_count_8_io_out ? io_r_427_b : _GEN_6516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6518 = 10'h1ac == r_count_8_io_out ? io_r_428_b : _GEN_6517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6519 = 10'h1ad == r_count_8_io_out ? io_r_429_b : _GEN_6518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6520 = 10'h1ae == r_count_8_io_out ? io_r_430_b : _GEN_6519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6521 = 10'h1af == r_count_8_io_out ? io_r_431_b : _GEN_6520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6522 = 10'h1b0 == r_count_8_io_out ? io_r_432_b : _GEN_6521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6523 = 10'h1b1 == r_count_8_io_out ? io_r_433_b : _GEN_6522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6524 = 10'h1b2 == r_count_8_io_out ? io_r_434_b : _GEN_6523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6525 = 10'h1b3 == r_count_8_io_out ? io_r_435_b : _GEN_6524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6526 = 10'h1b4 == r_count_8_io_out ? io_r_436_b : _GEN_6525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6527 = 10'h1b5 == r_count_8_io_out ? io_r_437_b : _GEN_6526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6528 = 10'h1b6 == r_count_8_io_out ? io_r_438_b : _GEN_6527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6529 = 10'h1b7 == r_count_8_io_out ? io_r_439_b : _GEN_6528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6530 = 10'h1b8 == r_count_8_io_out ? io_r_440_b : _GEN_6529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6531 = 10'h1b9 == r_count_8_io_out ? io_r_441_b : _GEN_6530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6532 = 10'h1ba == r_count_8_io_out ? io_r_442_b : _GEN_6531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6533 = 10'h1bb == r_count_8_io_out ? io_r_443_b : _GEN_6532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6534 = 10'h1bc == r_count_8_io_out ? io_r_444_b : _GEN_6533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6535 = 10'h1bd == r_count_8_io_out ? io_r_445_b : _GEN_6534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6536 = 10'h1be == r_count_8_io_out ? io_r_446_b : _GEN_6535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6537 = 10'h1bf == r_count_8_io_out ? io_r_447_b : _GEN_6536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6538 = 10'h1c0 == r_count_8_io_out ? io_r_448_b : _GEN_6537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6539 = 10'h1c1 == r_count_8_io_out ? io_r_449_b : _GEN_6538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6540 = 10'h1c2 == r_count_8_io_out ? io_r_450_b : _GEN_6539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6541 = 10'h1c3 == r_count_8_io_out ? io_r_451_b : _GEN_6540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6542 = 10'h1c4 == r_count_8_io_out ? io_r_452_b : _GEN_6541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6543 = 10'h1c5 == r_count_8_io_out ? io_r_453_b : _GEN_6542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6544 = 10'h1c6 == r_count_8_io_out ? io_r_454_b : _GEN_6543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6545 = 10'h1c7 == r_count_8_io_out ? io_r_455_b : _GEN_6544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6546 = 10'h1c8 == r_count_8_io_out ? io_r_456_b : _GEN_6545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6547 = 10'h1c9 == r_count_8_io_out ? io_r_457_b : _GEN_6546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6548 = 10'h1ca == r_count_8_io_out ? io_r_458_b : _GEN_6547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6549 = 10'h1cb == r_count_8_io_out ? io_r_459_b : _GEN_6548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6550 = 10'h1cc == r_count_8_io_out ? io_r_460_b : _GEN_6549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6551 = 10'h1cd == r_count_8_io_out ? io_r_461_b : _GEN_6550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6552 = 10'h1ce == r_count_8_io_out ? io_r_462_b : _GEN_6551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6553 = 10'h1cf == r_count_8_io_out ? io_r_463_b : _GEN_6552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6554 = 10'h1d0 == r_count_8_io_out ? io_r_464_b : _GEN_6553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6555 = 10'h1d1 == r_count_8_io_out ? io_r_465_b : _GEN_6554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6556 = 10'h1d2 == r_count_8_io_out ? io_r_466_b : _GEN_6555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6557 = 10'h1d3 == r_count_8_io_out ? io_r_467_b : _GEN_6556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6558 = 10'h1d4 == r_count_8_io_out ? io_r_468_b : _GEN_6557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6559 = 10'h1d5 == r_count_8_io_out ? io_r_469_b : _GEN_6558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6560 = 10'h1d6 == r_count_8_io_out ? io_r_470_b : _GEN_6559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6561 = 10'h1d7 == r_count_8_io_out ? io_r_471_b : _GEN_6560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6562 = 10'h1d8 == r_count_8_io_out ? io_r_472_b : _GEN_6561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6563 = 10'h1d9 == r_count_8_io_out ? io_r_473_b : _GEN_6562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6564 = 10'h1da == r_count_8_io_out ? io_r_474_b : _GEN_6563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6565 = 10'h1db == r_count_8_io_out ? io_r_475_b : _GEN_6564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6566 = 10'h1dc == r_count_8_io_out ? io_r_476_b : _GEN_6565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6567 = 10'h1dd == r_count_8_io_out ? io_r_477_b : _GEN_6566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6568 = 10'h1de == r_count_8_io_out ? io_r_478_b : _GEN_6567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6569 = 10'h1df == r_count_8_io_out ? io_r_479_b : _GEN_6568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6570 = 10'h1e0 == r_count_8_io_out ? io_r_480_b : _GEN_6569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6571 = 10'h1e1 == r_count_8_io_out ? io_r_481_b : _GEN_6570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6572 = 10'h1e2 == r_count_8_io_out ? io_r_482_b : _GEN_6571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6573 = 10'h1e3 == r_count_8_io_out ? io_r_483_b : _GEN_6572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6574 = 10'h1e4 == r_count_8_io_out ? io_r_484_b : _GEN_6573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6575 = 10'h1e5 == r_count_8_io_out ? io_r_485_b : _GEN_6574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6576 = 10'h1e6 == r_count_8_io_out ? io_r_486_b : _GEN_6575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6577 = 10'h1e7 == r_count_8_io_out ? io_r_487_b : _GEN_6576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6578 = 10'h1e8 == r_count_8_io_out ? io_r_488_b : _GEN_6577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6579 = 10'h1e9 == r_count_8_io_out ? io_r_489_b : _GEN_6578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6580 = 10'h1ea == r_count_8_io_out ? io_r_490_b : _GEN_6579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6581 = 10'h1eb == r_count_8_io_out ? io_r_491_b : _GEN_6580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6582 = 10'h1ec == r_count_8_io_out ? io_r_492_b : _GEN_6581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6583 = 10'h1ed == r_count_8_io_out ? io_r_493_b : _GEN_6582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6584 = 10'h1ee == r_count_8_io_out ? io_r_494_b : _GEN_6583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6585 = 10'h1ef == r_count_8_io_out ? io_r_495_b : _GEN_6584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6586 = 10'h1f0 == r_count_8_io_out ? io_r_496_b : _GEN_6585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6587 = 10'h1f1 == r_count_8_io_out ? io_r_497_b : _GEN_6586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6588 = 10'h1f2 == r_count_8_io_out ? io_r_498_b : _GEN_6587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6589 = 10'h1f3 == r_count_8_io_out ? io_r_499_b : _GEN_6588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6590 = 10'h1f4 == r_count_8_io_out ? io_r_500_b : _GEN_6589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6591 = 10'h1f5 == r_count_8_io_out ? io_r_501_b : _GEN_6590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6592 = 10'h1f6 == r_count_8_io_out ? io_r_502_b : _GEN_6591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6593 = 10'h1f7 == r_count_8_io_out ? io_r_503_b : _GEN_6592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6594 = 10'h1f8 == r_count_8_io_out ? io_r_504_b : _GEN_6593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6595 = 10'h1f9 == r_count_8_io_out ? io_r_505_b : _GEN_6594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6596 = 10'h1fa == r_count_8_io_out ? io_r_506_b : _GEN_6595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6597 = 10'h1fb == r_count_8_io_out ? io_r_507_b : _GEN_6596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6598 = 10'h1fc == r_count_8_io_out ? io_r_508_b : _GEN_6597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6599 = 10'h1fd == r_count_8_io_out ? io_r_509_b : _GEN_6598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6600 = 10'h1fe == r_count_8_io_out ? io_r_510_b : _GEN_6599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6601 = 10'h1ff == r_count_8_io_out ? io_r_511_b : _GEN_6600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6602 = 10'h200 == r_count_8_io_out ? io_r_512_b : _GEN_6601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6603 = 10'h201 == r_count_8_io_out ? io_r_513_b : _GEN_6602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6604 = 10'h202 == r_count_8_io_out ? io_r_514_b : _GEN_6603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6605 = 10'h203 == r_count_8_io_out ? io_r_515_b : _GEN_6604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6606 = 10'h204 == r_count_8_io_out ? io_r_516_b : _GEN_6605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6607 = 10'h205 == r_count_8_io_out ? io_r_517_b : _GEN_6606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6608 = 10'h206 == r_count_8_io_out ? io_r_518_b : _GEN_6607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6609 = 10'h207 == r_count_8_io_out ? io_r_519_b : _GEN_6608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6610 = 10'h208 == r_count_8_io_out ? io_r_520_b : _GEN_6609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6611 = 10'h209 == r_count_8_io_out ? io_r_521_b : _GEN_6610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6612 = 10'h20a == r_count_8_io_out ? io_r_522_b : _GEN_6611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6613 = 10'h20b == r_count_8_io_out ? io_r_523_b : _GEN_6612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6614 = 10'h20c == r_count_8_io_out ? io_r_524_b : _GEN_6613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6615 = 10'h20d == r_count_8_io_out ? io_r_525_b : _GEN_6614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6616 = 10'h20e == r_count_8_io_out ? io_r_526_b : _GEN_6615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6617 = 10'h20f == r_count_8_io_out ? io_r_527_b : _GEN_6616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6618 = 10'h210 == r_count_8_io_out ? io_r_528_b : _GEN_6617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6619 = 10'h211 == r_count_8_io_out ? io_r_529_b : _GEN_6618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6620 = 10'h212 == r_count_8_io_out ? io_r_530_b : _GEN_6619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6621 = 10'h213 == r_count_8_io_out ? io_r_531_b : _GEN_6620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6622 = 10'h214 == r_count_8_io_out ? io_r_532_b : _GEN_6621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6623 = 10'h215 == r_count_8_io_out ? io_r_533_b : _GEN_6622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6624 = 10'h216 == r_count_8_io_out ? io_r_534_b : _GEN_6623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6625 = 10'h217 == r_count_8_io_out ? io_r_535_b : _GEN_6624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6626 = 10'h218 == r_count_8_io_out ? io_r_536_b : _GEN_6625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6627 = 10'h219 == r_count_8_io_out ? io_r_537_b : _GEN_6626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6628 = 10'h21a == r_count_8_io_out ? io_r_538_b : _GEN_6627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6629 = 10'h21b == r_count_8_io_out ? io_r_539_b : _GEN_6628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6630 = 10'h21c == r_count_8_io_out ? io_r_540_b : _GEN_6629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6631 = 10'h21d == r_count_8_io_out ? io_r_541_b : _GEN_6630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6632 = 10'h21e == r_count_8_io_out ? io_r_542_b : _GEN_6631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6633 = 10'h21f == r_count_8_io_out ? io_r_543_b : _GEN_6632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6634 = 10'h220 == r_count_8_io_out ? io_r_544_b : _GEN_6633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6635 = 10'h221 == r_count_8_io_out ? io_r_545_b : _GEN_6634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6636 = 10'h222 == r_count_8_io_out ? io_r_546_b : _GEN_6635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6637 = 10'h223 == r_count_8_io_out ? io_r_547_b : _GEN_6636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6638 = 10'h224 == r_count_8_io_out ? io_r_548_b : _GEN_6637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6639 = 10'h225 == r_count_8_io_out ? io_r_549_b : _GEN_6638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6640 = 10'h226 == r_count_8_io_out ? io_r_550_b : _GEN_6639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6641 = 10'h227 == r_count_8_io_out ? io_r_551_b : _GEN_6640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6642 = 10'h228 == r_count_8_io_out ? io_r_552_b : _GEN_6641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6643 = 10'h229 == r_count_8_io_out ? io_r_553_b : _GEN_6642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6644 = 10'h22a == r_count_8_io_out ? io_r_554_b : _GEN_6643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6645 = 10'h22b == r_count_8_io_out ? io_r_555_b : _GEN_6644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6646 = 10'h22c == r_count_8_io_out ? io_r_556_b : _GEN_6645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6647 = 10'h22d == r_count_8_io_out ? io_r_557_b : _GEN_6646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6648 = 10'h22e == r_count_8_io_out ? io_r_558_b : _GEN_6647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6649 = 10'h22f == r_count_8_io_out ? io_r_559_b : _GEN_6648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6650 = 10'h230 == r_count_8_io_out ? io_r_560_b : _GEN_6649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6651 = 10'h231 == r_count_8_io_out ? io_r_561_b : _GEN_6650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6652 = 10'h232 == r_count_8_io_out ? io_r_562_b : _GEN_6651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6653 = 10'h233 == r_count_8_io_out ? io_r_563_b : _GEN_6652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6654 = 10'h234 == r_count_8_io_out ? io_r_564_b : _GEN_6653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6655 = 10'h235 == r_count_8_io_out ? io_r_565_b : _GEN_6654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6656 = 10'h236 == r_count_8_io_out ? io_r_566_b : _GEN_6655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6657 = 10'h237 == r_count_8_io_out ? io_r_567_b : _GEN_6656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6658 = 10'h238 == r_count_8_io_out ? io_r_568_b : _GEN_6657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6659 = 10'h239 == r_count_8_io_out ? io_r_569_b : _GEN_6658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6660 = 10'h23a == r_count_8_io_out ? io_r_570_b : _GEN_6659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6661 = 10'h23b == r_count_8_io_out ? io_r_571_b : _GEN_6660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6662 = 10'h23c == r_count_8_io_out ? io_r_572_b : _GEN_6661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6663 = 10'h23d == r_count_8_io_out ? io_r_573_b : _GEN_6662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6664 = 10'h23e == r_count_8_io_out ? io_r_574_b : _GEN_6663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6665 = 10'h23f == r_count_8_io_out ? io_r_575_b : _GEN_6664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6666 = 10'h240 == r_count_8_io_out ? io_r_576_b : _GEN_6665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6667 = 10'h241 == r_count_8_io_out ? io_r_577_b : _GEN_6666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6668 = 10'h242 == r_count_8_io_out ? io_r_578_b : _GEN_6667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6669 = 10'h243 == r_count_8_io_out ? io_r_579_b : _GEN_6668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6670 = 10'h244 == r_count_8_io_out ? io_r_580_b : _GEN_6669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6671 = 10'h245 == r_count_8_io_out ? io_r_581_b : _GEN_6670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6672 = 10'h246 == r_count_8_io_out ? io_r_582_b : _GEN_6671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6673 = 10'h247 == r_count_8_io_out ? io_r_583_b : _GEN_6672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6674 = 10'h248 == r_count_8_io_out ? io_r_584_b : _GEN_6673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6675 = 10'h249 == r_count_8_io_out ? io_r_585_b : _GEN_6674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6676 = 10'h24a == r_count_8_io_out ? io_r_586_b : _GEN_6675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6677 = 10'h24b == r_count_8_io_out ? io_r_587_b : _GEN_6676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6678 = 10'h24c == r_count_8_io_out ? io_r_588_b : _GEN_6677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6679 = 10'h24d == r_count_8_io_out ? io_r_589_b : _GEN_6678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6680 = 10'h24e == r_count_8_io_out ? io_r_590_b : _GEN_6679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6681 = 10'h24f == r_count_8_io_out ? io_r_591_b : _GEN_6680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6682 = 10'h250 == r_count_8_io_out ? io_r_592_b : _GEN_6681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6683 = 10'h251 == r_count_8_io_out ? io_r_593_b : _GEN_6682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6684 = 10'h252 == r_count_8_io_out ? io_r_594_b : _GEN_6683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6685 = 10'h253 == r_count_8_io_out ? io_r_595_b : _GEN_6684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6686 = 10'h254 == r_count_8_io_out ? io_r_596_b : _GEN_6685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6687 = 10'h255 == r_count_8_io_out ? io_r_597_b : _GEN_6686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6688 = 10'h256 == r_count_8_io_out ? io_r_598_b : _GEN_6687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6689 = 10'h257 == r_count_8_io_out ? io_r_599_b : _GEN_6688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6690 = 10'h258 == r_count_8_io_out ? io_r_600_b : _GEN_6689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6691 = 10'h259 == r_count_8_io_out ? io_r_601_b : _GEN_6690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6692 = 10'h25a == r_count_8_io_out ? io_r_602_b : _GEN_6691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6693 = 10'h25b == r_count_8_io_out ? io_r_603_b : _GEN_6692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6694 = 10'h25c == r_count_8_io_out ? io_r_604_b : _GEN_6693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6695 = 10'h25d == r_count_8_io_out ? io_r_605_b : _GEN_6694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6696 = 10'h25e == r_count_8_io_out ? io_r_606_b : _GEN_6695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6697 = 10'h25f == r_count_8_io_out ? io_r_607_b : _GEN_6696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6698 = 10'h260 == r_count_8_io_out ? io_r_608_b : _GEN_6697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6699 = 10'h261 == r_count_8_io_out ? io_r_609_b : _GEN_6698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6700 = 10'h262 == r_count_8_io_out ? io_r_610_b : _GEN_6699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6701 = 10'h263 == r_count_8_io_out ? io_r_611_b : _GEN_6700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6702 = 10'h264 == r_count_8_io_out ? io_r_612_b : _GEN_6701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6703 = 10'h265 == r_count_8_io_out ? io_r_613_b : _GEN_6702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6704 = 10'h266 == r_count_8_io_out ? io_r_614_b : _GEN_6703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6705 = 10'h267 == r_count_8_io_out ? io_r_615_b : _GEN_6704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6706 = 10'h268 == r_count_8_io_out ? io_r_616_b : _GEN_6705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6707 = 10'h269 == r_count_8_io_out ? io_r_617_b : _GEN_6706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6708 = 10'h26a == r_count_8_io_out ? io_r_618_b : _GEN_6707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6709 = 10'h26b == r_count_8_io_out ? io_r_619_b : _GEN_6708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6710 = 10'h26c == r_count_8_io_out ? io_r_620_b : _GEN_6709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6711 = 10'h26d == r_count_8_io_out ? io_r_621_b : _GEN_6710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6712 = 10'h26e == r_count_8_io_out ? io_r_622_b : _GEN_6711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6713 = 10'h26f == r_count_8_io_out ? io_r_623_b : _GEN_6712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6714 = 10'h270 == r_count_8_io_out ? io_r_624_b : _GEN_6713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6715 = 10'h271 == r_count_8_io_out ? io_r_625_b : _GEN_6714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6716 = 10'h272 == r_count_8_io_out ? io_r_626_b : _GEN_6715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6717 = 10'h273 == r_count_8_io_out ? io_r_627_b : _GEN_6716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6718 = 10'h274 == r_count_8_io_out ? io_r_628_b : _GEN_6717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6719 = 10'h275 == r_count_8_io_out ? io_r_629_b : _GEN_6718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6720 = 10'h276 == r_count_8_io_out ? io_r_630_b : _GEN_6719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6721 = 10'h277 == r_count_8_io_out ? io_r_631_b : _GEN_6720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6722 = 10'h278 == r_count_8_io_out ? io_r_632_b : _GEN_6721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6723 = 10'h279 == r_count_8_io_out ? io_r_633_b : _GEN_6722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6724 = 10'h27a == r_count_8_io_out ? io_r_634_b : _GEN_6723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6725 = 10'h27b == r_count_8_io_out ? io_r_635_b : _GEN_6724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6726 = 10'h27c == r_count_8_io_out ? io_r_636_b : _GEN_6725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6727 = 10'h27d == r_count_8_io_out ? io_r_637_b : _GEN_6726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6728 = 10'h27e == r_count_8_io_out ? io_r_638_b : _GEN_6727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6729 = 10'h27f == r_count_8_io_out ? io_r_639_b : _GEN_6728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6730 = 10'h280 == r_count_8_io_out ? io_r_640_b : _GEN_6729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6731 = 10'h281 == r_count_8_io_out ? io_r_641_b : _GEN_6730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6732 = 10'h282 == r_count_8_io_out ? io_r_642_b : _GEN_6731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6733 = 10'h283 == r_count_8_io_out ? io_r_643_b : _GEN_6732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6734 = 10'h284 == r_count_8_io_out ? io_r_644_b : _GEN_6733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6735 = 10'h285 == r_count_8_io_out ? io_r_645_b : _GEN_6734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6736 = 10'h286 == r_count_8_io_out ? io_r_646_b : _GEN_6735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6737 = 10'h287 == r_count_8_io_out ? io_r_647_b : _GEN_6736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6738 = 10'h288 == r_count_8_io_out ? io_r_648_b : _GEN_6737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6739 = 10'h289 == r_count_8_io_out ? io_r_649_b : _GEN_6738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6740 = 10'h28a == r_count_8_io_out ? io_r_650_b : _GEN_6739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6741 = 10'h28b == r_count_8_io_out ? io_r_651_b : _GEN_6740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6742 = 10'h28c == r_count_8_io_out ? io_r_652_b : _GEN_6741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6743 = 10'h28d == r_count_8_io_out ? io_r_653_b : _GEN_6742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6744 = 10'h28e == r_count_8_io_out ? io_r_654_b : _GEN_6743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6745 = 10'h28f == r_count_8_io_out ? io_r_655_b : _GEN_6744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6746 = 10'h290 == r_count_8_io_out ? io_r_656_b : _GEN_6745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6747 = 10'h291 == r_count_8_io_out ? io_r_657_b : _GEN_6746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6748 = 10'h292 == r_count_8_io_out ? io_r_658_b : _GEN_6747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6749 = 10'h293 == r_count_8_io_out ? io_r_659_b : _GEN_6748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6750 = 10'h294 == r_count_8_io_out ? io_r_660_b : _GEN_6749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6751 = 10'h295 == r_count_8_io_out ? io_r_661_b : _GEN_6750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6752 = 10'h296 == r_count_8_io_out ? io_r_662_b : _GEN_6751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6753 = 10'h297 == r_count_8_io_out ? io_r_663_b : _GEN_6752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6754 = 10'h298 == r_count_8_io_out ? io_r_664_b : _GEN_6753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6755 = 10'h299 == r_count_8_io_out ? io_r_665_b : _GEN_6754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6756 = 10'h29a == r_count_8_io_out ? io_r_666_b : _GEN_6755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6757 = 10'h29b == r_count_8_io_out ? io_r_667_b : _GEN_6756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6758 = 10'h29c == r_count_8_io_out ? io_r_668_b : _GEN_6757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6759 = 10'h29d == r_count_8_io_out ? io_r_669_b : _GEN_6758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6760 = 10'h29e == r_count_8_io_out ? io_r_670_b : _GEN_6759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6761 = 10'h29f == r_count_8_io_out ? io_r_671_b : _GEN_6760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6762 = 10'h2a0 == r_count_8_io_out ? io_r_672_b : _GEN_6761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6763 = 10'h2a1 == r_count_8_io_out ? io_r_673_b : _GEN_6762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6764 = 10'h2a2 == r_count_8_io_out ? io_r_674_b : _GEN_6763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6765 = 10'h2a3 == r_count_8_io_out ? io_r_675_b : _GEN_6764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6766 = 10'h2a4 == r_count_8_io_out ? io_r_676_b : _GEN_6765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6767 = 10'h2a5 == r_count_8_io_out ? io_r_677_b : _GEN_6766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6768 = 10'h2a6 == r_count_8_io_out ? io_r_678_b : _GEN_6767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6769 = 10'h2a7 == r_count_8_io_out ? io_r_679_b : _GEN_6768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6770 = 10'h2a8 == r_count_8_io_out ? io_r_680_b : _GEN_6769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6771 = 10'h2a9 == r_count_8_io_out ? io_r_681_b : _GEN_6770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6772 = 10'h2aa == r_count_8_io_out ? io_r_682_b : _GEN_6771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6773 = 10'h2ab == r_count_8_io_out ? io_r_683_b : _GEN_6772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6774 = 10'h2ac == r_count_8_io_out ? io_r_684_b : _GEN_6773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6775 = 10'h2ad == r_count_8_io_out ? io_r_685_b : _GEN_6774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6776 = 10'h2ae == r_count_8_io_out ? io_r_686_b : _GEN_6775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6777 = 10'h2af == r_count_8_io_out ? io_r_687_b : _GEN_6776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6778 = 10'h2b0 == r_count_8_io_out ? io_r_688_b : _GEN_6777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6779 = 10'h2b1 == r_count_8_io_out ? io_r_689_b : _GEN_6778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6780 = 10'h2b2 == r_count_8_io_out ? io_r_690_b : _GEN_6779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6781 = 10'h2b3 == r_count_8_io_out ? io_r_691_b : _GEN_6780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6782 = 10'h2b4 == r_count_8_io_out ? io_r_692_b : _GEN_6781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6783 = 10'h2b5 == r_count_8_io_out ? io_r_693_b : _GEN_6782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6784 = 10'h2b6 == r_count_8_io_out ? io_r_694_b : _GEN_6783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6785 = 10'h2b7 == r_count_8_io_out ? io_r_695_b : _GEN_6784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6786 = 10'h2b8 == r_count_8_io_out ? io_r_696_b : _GEN_6785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6787 = 10'h2b9 == r_count_8_io_out ? io_r_697_b : _GEN_6786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6788 = 10'h2ba == r_count_8_io_out ? io_r_698_b : _GEN_6787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6789 = 10'h2bb == r_count_8_io_out ? io_r_699_b : _GEN_6788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6790 = 10'h2bc == r_count_8_io_out ? io_r_700_b : _GEN_6789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6791 = 10'h2bd == r_count_8_io_out ? io_r_701_b : _GEN_6790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6792 = 10'h2be == r_count_8_io_out ? io_r_702_b : _GEN_6791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6793 = 10'h2bf == r_count_8_io_out ? io_r_703_b : _GEN_6792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6794 = 10'h2c0 == r_count_8_io_out ? io_r_704_b : _GEN_6793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6795 = 10'h2c1 == r_count_8_io_out ? io_r_705_b : _GEN_6794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6796 = 10'h2c2 == r_count_8_io_out ? io_r_706_b : _GEN_6795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6797 = 10'h2c3 == r_count_8_io_out ? io_r_707_b : _GEN_6796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6798 = 10'h2c4 == r_count_8_io_out ? io_r_708_b : _GEN_6797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6799 = 10'h2c5 == r_count_8_io_out ? io_r_709_b : _GEN_6798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6800 = 10'h2c6 == r_count_8_io_out ? io_r_710_b : _GEN_6799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6801 = 10'h2c7 == r_count_8_io_out ? io_r_711_b : _GEN_6800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6802 = 10'h2c8 == r_count_8_io_out ? io_r_712_b : _GEN_6801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6803 = 10'h2c9 == r_count_8_io_out ? io_r_713_b : _GEN_6802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6804 = 10'h2ca == r_count_8_io_out ? io_r_714_b : _GEN_6803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6805 = 10'h2cb == r_count_8_io_out ? io_r_715_b : _GEN_6804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6806 = 10'h2cc == r_count_8_io_out ? io_r_716_b : _GEN_6805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6807 = 10'h2cd == r_count_8_io_out ? io_r_717_b : _GEN_6806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6808 = 10'h2ce == r_count_8_io_out ? io_r_718_b : _GEN_6807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6809 = 10'h2cf == r_count_8_io_out ? io_r_719_b : _GEN_6808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6810 = 10'h2d0 == r_count_8_io_out ? io_r_720_b : _GEN_6809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6811 = 10'h2d1 == r_count_8_io_out ? io_r_721_b : _GEN_6810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6812 = 10'h2d2 == r_count_8_io_out ? io_r_722_b : _GEN_6811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6813 = 10'h2d3 == r_count_8_io_out ? io_r_723_b : _GEN_6812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6814 = 10'h2d4 == r_count_8_io_out ? io_r_724_b : _GEN_6813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6815 = 10'h2d5 == r_count_8_io_out ? io_r_725_b : _GEN_6814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6816 = 10'h2d6 == r_count_8_io_out ? io_r_726_b : _GEN_6815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6817 = 10'h2d7 == r_count_8_io_out ? io_r_727_b : _GEN_6816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6818 = 10'h2d8 == r_count_8_io_out ? io_r_728_b : _GEN_6817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6819 = 10'h2d9 == r_count_8_io_out ? io_r_729_b : _GEN_6818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6820 = 10'h2da == r_count_8_io_out ? io_r_730_b : _GEN_6819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6821 = 10'h2db == r_count_8_io_out ? io_r_731_b : _GEN_6820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6822 = 10'h2dc == r_count_8_io_out ? io_r_732_b : _GEN_6821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6823 = 10'h2dd == r_count_8_io_out ? io_r_733_b : _GEN_6822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6824 = 10'h2de == r_count_8_io_out ? io_r_734_b : _GEN_6823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6825 = 10'h2df == r_count_8_io_out ? io_r_735_b : _GEN_6824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6826 = 10'h2e0 == r_count_8_io_out ? io_r_736_b : _GEN_6825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6827 = 10'h2e1 == r_count_8_io_out ? io_r_737_b : _GEN_6826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6828 = 10'h2e2 == r_count_8_io_out ? io_r_738_b : _GEN_6827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6829 = 10'h2e3 == r_count_8_io_out ? io_r_739_b : _GEN_6828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6830 = 10'h2e4 == r_count_8_io_out ? io_r_740_b : _GEN_6829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6831 = 10'h2e5 == r_count_8_io_out ? io_r_741_b : _GEN_6830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6832 = 10'h2e6 == r_count_8_io_out ? io_r_742_b : _GEN_6831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6833 = 10'h2e7 == r_count_8_io_out ? io_r_743_b : _GEN_6832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6834 = 10'h2e8 == r_count_8_io_out ? io_r_744_b : _GEN_6833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6835 = 10'h2e9 == r_count_8_io_out ? io_r_745_b : _GEN_6834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6836 = 10'h2ea == r_count_8_io_out ? io_r_746_b : _GEN_6835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6837 = 10'h2eb == r_count_8_io_out ? io_r_747_b : _GEN_6836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6838 = 10'h2ec == r_count_8_io_out ? io_r_748_b : _GEN_6837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6841 = 10'h1 == r_count_9_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6842 = 10'h2 == r_count_9_io_out ? io_r_2_b : _GEN_6841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6843 = 10'h3 == r_count_9_io_out ? io_r_3_b : _GEN_6842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6844 = 10'h4 == r_count_9_io_out ? io_r_4_b : _GEN_6843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6845 = 10'h5 == r_count_9_io_out ? io_r_5_b : _GEN_6844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6846 = 10'h6 == r_count_9_io_out ? io_r_6_b : _GEN_6845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6847 = 10'h7 == r_count_9_io_out ? io_r_7_b : _GEN_6846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6848 = 10'h8 == r_count_9_io_out ? io_r_8_b : _GEN_6847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6849 = 10'h9 == r_count_9_io_out ? io_r_9_b : _GEN_6848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6850 = 10'ha == r_count_9_io_out ? io_r_10_b : _GEN_6849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6851 = 10'hb == r_count_9_io_out ? io_r_11_b : _GEN_6850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6852 = 10'hc == r_count_9_io_out ? io_r_12_b : _GEN_6851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6853 = 10'hd == r_count_9_io_out ? io_r_13_b : _GEN_6852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6854 = 10'he == r_count_9_io_out ? io_r_14_b : _GEN_6853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6855 = 10'hf == r_count_9_io_out ? io_r_15_b : _GEN_6854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6856 = 10'h10 == r_count_9_io_out ? io_r_16_b : _GEN_6855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6857 = 10'h11 == r_count_9_io_out ? io_r_17_b : _GEN_6856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6858 = 10'h12 == r_count_9_io_out ? io_r_18_b : _GEN_6857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6859 = 10'h13 == r_count_9_io_out ? io_r_19_b : _GEN_6858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6860 = 10'h14 == r_count_9_io_out ? io_r_20_b : _GEN_6859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6861 = 10'h15 == r_count_9_io_out ? io_r_21_b : _GEN_6860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6862 = 10'h16 == r_count_9_io_out ? io_r_22_b : _GEN_6861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6863 = 10'h17 == r_count_9_io_out ? io_r_23_b : _GEN_6862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6864 = 10'h18 == r_count_9_io_out ? io_r_24_b : _GEN_6863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6865 = 10'h19 == r_count_9_io_out ? io_r_25_b : _GEN_6864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6866 = 10'h1a == r_count_9_io_out ? io_r_26_b : _GEN_6865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6867 = 10'h1b == r_count_9_io_out ? io_r_27_b : _GEN_6866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6868 = 10'h1c == r_count_9_io_out ? io_r_28_b : _GEN_6867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6869 = 10'h1d == r_count_9_io_out ? io_r_29_b : _GEN_6868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6870 = 10'h1e == r_count_9_io_out ? io_r_30_b : _GEN_6869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6871 = 10'h1f == r_count_9_io_out ? io_r_31_b : _GEN_6870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6872 = 10'h20 == r_count_9_io_out ? io_r_32_b : _GEN_6871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6873 = 10'h21 == r_count_9_io_out ? io_r_33_b : _GEN_6872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6874 = 10'h22 == r_count_9_io_out ? io_r_34_b : _GEN_6873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6875 = 10'h23 == r_count_9_io_out ? io_r_35_b : _GEN_6874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6876 = 10'h24 == r_count_9_io_out ? io_r_36_b : _GEN_6875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6877 = 10'h25 == r_count_9_io_out ? io_r_37_b : _GEN_6876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6878 = 10'h26 == r_count_9_io_out ? io_r_38_b : _GEN_6877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6879 = 10'h27 == r_count_9_io_out ? io_r_39_b : _GEN_6878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6880 = 10'h28 == r_count_9_io_out ? io_r_40_b : _GEN_6879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6881 = 10'h29 == r_count_9_io_out ? io_r_41_b : _GEN_6880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6882 = 10'h2a == r_count_9_io_out ? io_r_42_b : _GEN_6881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6883 = 10'h2b == r_count_9_io_out ? io_r_43_b : _GEN_6882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6884 = 10'h2c == r_count_9_io_out ? io_r_44_b : _GEN_6883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6885 = 10'h2d == r_count_9_io_out ? io_r_45_b : _GEN_6884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6886 = 10'h2e == r_count_9_io_out ? io_r_46_b : _GEN_6885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6887 = 10'h2f == r_count_9_io_out ? io_r_47_b : _GEN_6886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6888 = 10'h30 == r_count_9_io_out ? io_r_48_b : _GEN_6887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6889 = 10'h31 == r_count_9_io_out ? io_r_49_b : _GEN_6888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6890 = 10'h32 == r_count_9_io_out ? io_r_50_b : _GEN_6889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6891 = 10'h33 == r_count_9_io_out ? io_r_51_b : _GEN_6890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6892 = 10'h34 == r_count_9_io_out ? io_r_52_b : _GEN_6891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6893 = 10'h35 == r_count_9_io_out ? io_r_53_b : _GEN_6892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6894 = 10'h36 == r_count_9_io_out ? io_r_54_b : _GEN_6893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6895 = 10'h37 == r_count_9_io_out ? io_r_55_b : _GEN_6894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6896 = 10'h38 == r_count_9_io_out ? io_r_56_b : _GEN_6895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6897 = 10'h39 == r_count_9_io_out ? io_r_57_b : _GEN_6896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6898 = 10'h3a == r_count_9_io_out ? io_r_58_b : _GEN_6897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6899 = 10'h3b == r_count_9_io_out ? io_r_59_b : _GEN_6898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6900 = 10'h3c == r_count_9_io_out ? io_r_60_b : _GEN_6899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6901 = 10'h3d == r_count_9_io_out ? io_r_61_b : _GEN_6900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6902 = 10'h3e == r_count_9_io_out ? io_r_62_b : _GEN_6901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6903 = 10'h3f == r_count_9_io_out ? io_r_63_b : _GEN_6902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6904 = 10'h40 == r_count_9_io_out ? io_r_64_b : _GEN_6903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6905 = 10'h41 == r_count_9_io_out ? io_r_65_b : _GEN_6904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6906 = 10'h42 == r_count_9_io_out ? io_r_66_b : _GEN_6905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6907 = 10'h43 == r_count_9_io_out ? io_r_67_b : _GEN_6906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6908 = 10'h44 == r_count_9_io_out ? io_r_68_b : _GEN_6907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6909 = 10'h45 == r_count_9_io_out ? io_r_69_b : _GEN_6908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6910 = 10'h46 == r_count_9_io_out ? io_r_70_b : _GEN_6909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6911 = 10'h47 == r_count_9_io_out ? io_r_71_b : _GEN_6910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6912 = 10'h48 == r_count_9_io_out ? io_r_72_b : _GEN_6911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6913 = 10'h49 == r_count_9_io_out ? io_r_73_b : _GEN_6912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6914 = 10'h4a == r_count_9_io_out ? io_r_74_b : _GEN_6913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6915 = 10'h4b == r_count_9_io_out ? io_r_75_b : _GEN_6914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6916 = 10'h4c == r_count_9_io_out ? io_r_76_b : _GEN_6915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6917 = 10'h4d == r_count_9_io_out ? io_r_77_b : _GEN_6916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6918 = 10'h4e == r_count_9_io_out ? io_r_78_b : _GEN_6917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6919 = 10'h4f == r_count_9_io_out ? io_r_79_b : _GEN_6918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6920 = 10'h50 == r_count_9_io_out ? io_r_80_b : _GEN_6919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6921 = 10'h51 == r_count_9_io_out ? io_r_81_b : _GEN_6920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6922 = 10'h52 == r_count_9_io_out ? io_r_82_b : _GEN_6921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6923 = 10'h53 == r_count_9_io_out ? io_r_83_b : _GEN_6922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6924 = 10'h54 == r_count_9_io_out ? io_r_84_b : _GEN_6923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6925 = 10'h55 == r_count_9_io_out ? io_r_85_b : _GEN_6924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6926 = 10'h56 == r_count_9_io_out ? io_r_86_b : _GEN_6925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6927 = 10'h57 == r_count_9_io_out ? io_r_87_b : _GEN_6926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6928 = 10'h58 == r_count_9_io_out ? io_r_88_b : _GEN_6927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6929 = 10'h59 == r_count_9_io_out ? io_r_89_b : _GEN_6928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6930 = 10'h5a == r_count_9_io_out ? io_r_90_b : _GEN_6929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6931 = 10'h5b == r_count_9_io_out ? io_r_91_b : _GEN_6930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6932 = 10'h5c == r_count_9_io_out ? io_r_92_b : _GEN_6931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6933 = 10'h5d == r_count_9_io_out ? io_r_93_b : _GEN_6932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6934 = 10'h5e == r_count_9_io_out ? io_r_94_b : _GEN_6933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6935 = 10'h5f == r_count_9_io_out ? io_r_95_b : _GEN_6934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6936 = 10'h60 == r_count_9_io_out ? io_r_96_b : _GEN_6935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6937 = 10'h61 == r_count_9_io_out ? io_r_97_b : _GEN_6936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6938 = 10'h62 == r_count_9_io_out ? io_r_98_b : _GEN_6937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6939 = 10'h63 == r_count_9_io_out ? io_r_99_b : _GEN_6938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6940 = 10'h64 == r_count_9_io_out ? io_r_100_b : _GEN_6939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6941 = 10'h65 == r_count_9_io_out ? io_r_101_b : _GEN_6940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6942 = 10'h66 == r_count_9_io_out ? io_r_102_b : _GEN_6941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6943 = 10'h67 == r_count_9_io_out ? io_r_103_b : _GEN_6942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6944 = 10'h68 == r_count_9_io_out ? io_r_104_b : _GEN_6943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6945 = 10'h69 == r_count_9_io_out ? io_r_105_b : _GEN_6944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6946 = 10'h6a == r_count_9_io_out ? io_r_106_b : _GEN_6945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6947 = 10'h6b == r_count_9_io_out ? io_r_107_b : _GEN_6946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6948 = 10'h6c == r_count_9_io_out ? io_r_108_b : _GEN_6947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6949 = 10'h6d == r_count_9_io_out ? io_r_109_b : _GEN_6948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6950 = 10'h6e == r_count_9_io_out ? io_r_110_b : _GEN_6949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6951 = 10'h6f == r_count_9_io_out ? io_r_111_b : _GEN_6950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6952 = 10'h70 == r_count_9_io_out ? io_r_112_b : _GEN_6951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6953 = 10'h71 == r_count_9_io_out ? io_r_113_b : _GEN_6952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6954 = 10'h72 == r_count_9_io_out ? io_r_114_b : _GEN_6953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6955 = 10'h73 == r_count_9_io_out ? io_r_115_b : _GEN_6954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6956 = 10'h74 == r_count_9_io_out ? io_r_116_b : _GEN_6955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6957 = 10'h75 == r_count_9_io_out ? io_r_117_b : _GEN_6956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6958 = 10'h76 == r_count_9_io_out ? io_r_118_b : _GEN_6957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6959 = 10'h77 == r_count_9_io_out ? io_r_119_b : _GEN_6958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6960 = 10'h78 == r_count_9_io_out ? io_r_120_b : _GEN_6959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6961 = 10'h79 == r_count_9_io_out ? io_r_121_b : _GEN_6960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6962 = 10'h7a == r_count_9_io_out ? io_r_122_b : _GEN_6961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6963 = 10'h7b == r_count_9_io_out ? io_r_123_b : _GEN_6962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6964 = 10'h7c == r_count_9_io_out ? io_r_124_b : _GEN_6963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6965 = 10'h7d == r_count_9_io_out ? io_r_125_b : _GEN_6964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6966 = 10'h7e == r_count_9_io_out ? io_r_126_b : _GEN_6965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6967 = 10'h7f == r_count_9_io_out ? io_r_127_b : _GEN_6966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6968 = 10'h80 == r_count_9_io_out ? io_r_128_b : _GEN_6967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6969 = 10'h81 == r_count_9_io_out ? io_r_129_b : _GEN_6968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6970 = 10'h82 == r_count_9_io_out ? io_r_130_b : _GEN_6969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6971 = 10'h83 == r_count_9_io_out ? io_r_131_b : _GEN_6970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6972 = 10'h84 == r_count_9_io_out ? io_r_132_b : _GEN_6971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6973 = 10'h85 == r_count_9_io_out ? io_r_133_b : _GEN_6972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6974 = 10'h86 == r_count_9_io_out ? io_r_134_b : _GEN_6973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6975 = 10'h87 == r_count_9_io_out ? io_r_135_b : _GEN_6974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6976 = 10'h88 == r_count_9_io_out ? io_r_136_b : _GEN_6975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6977 = 10'h89 == r_count_9_io_out ? io_r_137_b : _GEN_6976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6978 = 10'h8a == r_count_9_io_out ? io_r_138_b : _GEN_6977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6979 = 10'h8b == r_count_9_io_out ? io_r_139_b : _GEN_6978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6980 = 10'h8c == r_count_9_io_out ? io_r_140_b : _GEN_6979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6981 = 10'h8d == r_count_9_io_out ? io_r_141_b : _GEN_6980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6982 = 10'h8e == r_count_9_io_out ? io_r_142_b : _GEN_6981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6983 = 10'h8f == r_count_9_io_out ? io_r_143_b : _GEN_6982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6984 = 10'h90 == r_count_9_io_out ? io_r_144_b : _GEN_6983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6985 = 10'h91 == r_count_9_io_out ? io_r_145_b : _GEN_6984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6986 = 10'h92 == r_count_9_io_out ? io_r_146_b : _GEN_6985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6987 = 10'h93 == r_count_9_io_out ? io_r_147_b : _GEN_6986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6988 = 10'h94 == r_count_9_io_out ? io_r_148_b : _GEN_6987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6989 = 10'h95 == r_count_9_io_out ? io_r_149_b : _GEN_6988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6990 = 10'h96 == r_count_9_io_out ? io_r_150_b : _GEN_6989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6991 = 10'h97 == r_count_9_io_out ? io_r_151_b : _GEN_6990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6992 = 10'h98 == r_count_9_io_out ? io_r_152_b : _GEN_6991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6993 = 10'h99 == r_count_9_io_out ? io_r_153_b : _GEN_6992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6994 = 10'h9a == r_count_9_io_out ? io_r_154_b : _GEN_6993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6995 = 10'h9b == r_count_9_io_out ? io_r_155_b : _GEN_6994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6996 = 10'h9c == r_count_9_io_out ? io_r_156_b : _GEN_6995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6997 = 10'h9d == r_count_9_io_out ? io_r_157_b : _GEN_6996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6998 = 10'h9e == r_count_9_io_out ? io_r_158_b : _GEN_6997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6999 = 10'h9f == r_count_9_io_out ? io_r_159_b : _GEN_6998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7000 = 10'ha0 == r_count_9_io_out ? io_r_160_b : _GEN_6999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7001 = 10'ha1 == r_count_9_io_out ? io_r_161_b : _GEN_7000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7002 = 10'ha2 == r_count_9_io_out ? io_r_162_b : _GEN_7001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7003 = 10'ha3 == r_count_9_io_out ? io_r_163_b : _GEN_7002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7004 = 10'ha4 == r_count_9_io_out ? io_r_164_b : _GEN_7003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7005 = 10'ha5 == r_count_9_io_out ? io_r_165_b : _GEN_7004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7006 = 10'ha6 == r_count_9_io_out ? io_r_166_b : _GEN_7005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7007 = 10'ha7 == r_count_9_io_out ? io_r_167_b : _GEN_7006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7008 = 10'ha8 == r_count_9_io_out ? io_r_168_b : _GEN_7007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7009 = 10'ha9 == r_count_9_io_out ? io_r_169_b : _GEN_7008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7010 = 10'haa == r_count_9_io_out ? io_r_170_b : _GEN_7009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7011 = 10'hab == r_count_9_io_out ? io_r_171_b : _GEN_7010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7012 = 10'hac == r_count_9_io_out ? io_r_172_b : _GEN_7011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7013 = 10'had == r_count_9_io_out ? io_r_173_b : _GEN_7012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7014 = 10'hae == r_count_9_io_out ? io_r_174_b : _GEN_7013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7015 = 10'haf == r_count_9_io_out ? io_r_175_b : _GEN_7014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7016 = 10'hb0 == r_count_9_io_out ? io_r_176_b : _GEN_7015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7017 = 10'hb1 == r_count_9_io_out ? io_r_177_b : _GEN_7016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7018 = 10'hb2 == r_count_9_io_out ? io_r_178_b : _GEN_7017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7019 = 10'hb3 == r_count_9_io_out ? io_r_179_b : _GEN_7018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7020 = 10'hb4 == r_count_9_io_out ? io_r_180_b : _GEN_7019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7021 = 10'hb5 == r_count_9_io_out ? io_r_181_b : _GEN_7020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7022 = 10'hb6 == r_count_9_io_out ? io_r_182_b : _GEN_7021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7023 = 10'hb7 == r_count_9_io_out ? io_r_183_b : _GEN_7022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7024 = 10'hb8 == r_count_9_io_out ? io_r_184_b : _GEN_7023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7025 = 10'hb9 == r_count_9_io_out ? io_r_185_b : _GEN_7024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7026 = 10'hba == r_count_9_io_out ? io_r_186_b : _GEN_7025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7027 = 10'hbb == r_count_9_io_out ? io_r_187_b : _GEN_7026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7028 = 10'hbc == r_count_9_io_out ? io_r_188_b : _GEN_7027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7029 = 10'hbd == r_count_9_io_out ? io_r_189_b : _GEN_7028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7030 = 10'hbe == r_count_9_io_out ? io_r_190_b : _GEN_7029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7031 = 10'hbf == r_count_9_io_out ? io_r_191_b : _GEN_7030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7032 = 10'hc0 == r_count_9_io_out ? io_r_192_b : _GEN_7031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7033 = 10'hc1 == r_count_9_io_out ? io_r_193_b : _GEN_7032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7034 = 10'hc2 == r_count_9_io_out ? io_r_194_b : _GEN_7033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7035 = 10'hc3 == r_count_9_io_out ? io_r_195_b : _GEN_7034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7036 = 10'hc4 == r_count_9_io_out ? io_r_196_b : _GEN_7035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7037 = 10'hc5 == r_count_9_io_out ? io_r_197_b : _GEN_7036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7038 = 10'hc6 == r_count_9_io_out ? io_r_198_b : _GEN_7037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7039 = 10'hc7 == r_count_9_io_out ? io_r_199_b : _GEN_7038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7040 = 10'hc8 == r_count_9_io_out ? io_r_200_b : _GEN_7039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7041 = 10'hc9 == r_count_9_io_out ? io_r_201_b : _GEN_7040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7042 = 10'hca == r_count_9_io_out ? io_r_202_b : _GEN_7041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7043 = 10'hcb == r_count_9_io_out ? io_r_203_b : _GEN_7042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7044 = 10'hcc == r_count_9_io_out ? io_r_204_b : _GEN_7043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7045 = 10'hcd == r_count_9_io_out ? io_r_205_b : _GEN_7044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7046 = 10'hce == r_count_9_io_out ? io_r_206_b : _GEN_7045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7047 = 10'hcf == r_count_9_io_out ? io_r_207_b : _GEN_7046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7048 = 10'hd0 == r_count_9_io_out ? io_r_208_b : _GEN_7047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7049 = 10'hd1 == r_count_9_io_out ? io_r_209_b : _GEN_7048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7050 = 10'hd2 == r_count_9_io_out ? io_r_210_b : _GEN_7049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7051 = 10'hd3 == r_count_9_io_out ? io_r_211_b : _GEN_7050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7052 = 10'hd4 == r_count_9_io_out ? io_r_212_b : _GEN_7051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7053 = 10'hd5 == r_count_9_io_out ? io_r_213_b : _GEN_7052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7054 = 10'hd6 == r_count_9_io_out ? io_r_214_b : _GEN_7053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7055 = 10'hd7 == r_count_9_io_out ? io_r_215_b : _GEN_7054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7056 = 10'hd8 == r_count_9_io_out ? io_r_216_b : _GEN_7055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7057 = 10'hd9 == r_count_9_io_out ? io_r_217_b : _GEN_7056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7058 = 10'hda == r_count_9_io_out ? io_r_218_b : _GEN_7057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7059 = 10'hdb == r_count_9_io_out ? io_r_219_b : _GEN_7058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7060 = 10'hdc == r_count_9_io_out ? io_r_220_b : _GEN_7059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7061 = 10'hdd == r_count_9_io_out ? io_r_221_b : _GEN_7060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7062 = 10'hde == r_count_9_io_out ? io_r_222_b : _GEN_7061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7063 = 10'hdf == r_count_9_io_out ? io_r_223_b : _GEN_7062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7064 = 10'he0 == r_count_9_io_out ? io_r_224_b : _GEN_7063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7065 = 10'he1 == r_count_9_io_out ? io_r_225_b : _GEN_7064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7066 = 10'he2 == r_count_9_io_out ? io_r_226_b : _GEN_7065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7067 = 10'he3 == r_count_9_io_out ? io_r_227_b : _GEN_7066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7068 = 10'he4 == r_count_9_io_out ? io_r_228_b : _GEN_7067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7069 = 10'he5 == r_count_9_io_out ? io_r_229_b : _GEN_7068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7070 = 10'he6 == r_count_9_io_out ? io_r_230_b : _GEN_7069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7071 = 10'he7 == r_count_9_io_out ? io_r_231_b : _GEN_7070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7072 = 10'he8 == r_count_9_io_out ? io_r_232_b : _GEN_7071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7073 = 10'he9 == r_count_9_io_out ? io_r_233_b : _GEN_7072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7074 = 10'hea == r_count_9_io_out ? io_r_234_b : _GEN_7073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7075 = 10'heb == r_count_9_io_out ? io_r_235_b : _GEN_7074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7076 = 10'hec == r_count_9_io_out ? io_r_236_b : _GEN_7075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7077 = 10'hed == r_count_9_io_out ? io_r_237_b : _GEN_7076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7078 = 10'hee == r_count_9_io_out ? io_r_238_b : _GEN_7077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7079 = 10'hef == r_count_9_io_out ? io_r_239_b : _GEN_7078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7080 = 10'hf0 == r_count_9_io_out ? io_r_240_b : _GEN_7079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7081 = 10'hf1 == r_count_9_io_out ? io_r_241_b : _GEN_7080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7082 = 10'hf2 == r_count_9_io_out ? io_r_242_b : _GEN_7081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7083 = 10'hf3 == r_count_9_io_out ? io_r_243_b : _GEN_7082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7084 = 10'hf4 == r_count_9_io_out ? io_r_244_b : _GEN_7083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7085 = 10'hf5 == r_count_9_io_out ? io_r_245_b : _GEN_7084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7086 = 10'hf6 == r_count_9_io_out ? io_r_246_b : _GEN_7085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7087 = 10'hf7 == r_count_9_io_out ? io_r_247_b : _GEN_7086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7088 = 10'hf8 == r_count_9_io_out ? io_r_248_b : _GEN_7087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7089 = 10'hf9 == r_count_9_io_out ? io_r_249_b : _GEN_7088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7090 = 10'hfa == r_count_9_io_out ? io_r_250_b : _GEN_7089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7091 = 10'hfb == r_count_9_io_out ? io_r_251_b : _GEN_7090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7092 = 10'hfc == r_count_9_io_out ? io_r_252_b : _GEN_7091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7093 = 10'hfd == r_count_9_io_out ? io_r_253_b : _GEN_7092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7094 = 10'hfe == r_count_9_io_out ? io_r_254_b : _GEN_7093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7095 = 10'hff == r_count_9_io_out ? io_r_255_b : _GEN_7094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7096 = 10'h100 == r_count_9_io_out ? io_r_256_b : _GEN_7095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7097 = 10'h101 == r_count_9_io_out ? io_r_257_b : _GEN_7096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7098 = 10'h102 == r_count_9_io_out ? io_r_258_b : _GEN_7097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7099 = 10'h103 == r_count_9_io_out ? io_r_259_b : _GEN_7098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7100 = 10'h104 == r_count_9_io_out ? io_r_260_b : _GEN_7099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7101 = 10'h105 == r_count_9_io_out ? io_r_261_b : _GEN_7100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7102 = 10'h106 == r_count_9_io_out ? io_r_262_b : _GEN_7101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7103 = 10'h107 == r_count_9_io_out ? io_r_263_b : _GEN_7102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7104 = 10'h108 == r_count_9_io_out ? io_r_264_b : _GEN_7103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7105 = 10'h109 == r_count_9_io_out ? io_r_265_b : _GEN_7104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7106 = 10'h10a == r_count_9_io_out ? io_r_266_b : _GEN_7105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7107 = 10'h10b == r_count_9_io_out ? io_r_267_b : _GEN_7106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7108 = 10'h10c == r_count_9_io_out ? io_r_268_b : _GEN_7107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7109 = 10'h10d == r_count_9_io_out ? io_r_269_b : _GEN_7108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7110 = 10'h10e == r_count_9_io_out ? io_r_270_b : _GEN_7109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7111 = 10'h10f == r_count_9_io_out ? io_r_271_b : _GEN_7110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7112 = 10'h110 == r_count_9_io_out ? io_r_272_b : _GEN_7111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7113 = 10'h111 == r_count_9_io_out ? io_r_273_b : _GEN_7112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7114 = 10'h112 == r_count_9_io_out ? io_r_274_b : _GEN_7113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7115 = 10'h113 == r_count_9_io_out ? io_r_275_b : _GEN_7114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7116 = 10'h114 == r_count_9_io_out ? io_r_276_b : _GEN_7115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7117 = 10'h115 == r_count_9_io_out ? io_r_277_b : _GEN_7116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7118 = 10'h116 == r_count_9_io_out ? io_r_278_b : _GEN_7117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7119 = 10'h117 == r_count_9_io_out ? io_r_279_b : _GEN_7118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7120 = 10'h118 == r_count_9_io_out ? io_r_280_b : _GEN_7119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7121 = 10'h119 == r_count_9_io_out ? io_r_281_b : _GEN_7120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7122 = 10'h11a == r_count_9_io_out ? io_r_282_b : _GEN_7121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7123 = 10'h11b == r_count_9_io_out ? io_r_283_b : _GEN_7122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7124 = 10'h11c == r_count_9_io_out ? io_r_284_b : _GEN_7123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7125 = 10'h11d == r_count_9_io_out ? io_r_285_b : _GEN_7124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7126 = 10'h11e == r_count_9_io_out ? io_r_286_b : _GEN_7125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7127 = 10'h11f == r_count_9_io_out ? io_r_287_b : _GEN_7126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7128 = 10'h120 == r_count_9_io_out ? io_r_288_b : _GEN_7127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7129 = 10'h121 == r_count_9_io_out ? io_r_289_b : _GEN_7128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7130 = 10'h122 == r_count_9_io_out ? io_r_290_b : _GEN_7129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7131 = 10'h123 == r_count_9_io_out ? io_r_291_b : _GEN_7130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7132 = 10'h124 == r_count_9_io_out ? io_r_292_b : _GEN_7131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7133 = 10'h125 == r_count_9_io_out ? io_r_293_b : _GEN_7132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7134 = 10'h126 == r_count_9_io_out ? io_r_294_b : _GEN_7133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7135 = 10'h127 == r_count_9_io_out ? io_r_295_b : _GEN_7134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7136 = 10'h128 == r_count_9_io_out ? io_r_296_b : _GEN_7135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7137 = 10'h129 == r_count_9_io_out ? io_r_297_b : _GEN_7136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7138 = 10'h12a == r_count_9_io_out ? io_r_298_b : _GEN_7137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7139 = 10'h12b == r_count_9_io_out ? io_r_299_b : _GEN_7138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7140 = 10'h12c == r_count_9_io_out ? io_r_300_b : _GEN_7139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7141 = 10'h12d == r_count_9_io_out ? io_r_301_b : _GEN_7140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7142 = 10'h12e == r_count_9_io_out ? io_r_302_b : _GEN_7141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7143 = 10'h12f == r_count_9_io_out ? io_r_303_b : _GEN_7142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7144 = 10'h130 == r_count_9_io_out ? io_r_304_b : _GEN_7143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7145 = 10'h131 == r_count_9_io_out ? io_r_305_b : _GEN_7144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7146 = 10'h132 == r_count_9_io_out ? io_r_306_b : _GEN_7145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7147 = 10'h133 == r_count_9_io_out ? io_r_307_b : _GEN_7146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7148 = 10'h134 == r_count_9_io_out ? io_r_308_b : _GEN_7147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7149 = 10'h135 == r_count_9_io_out ? io_r_309_b : _GEN_7148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7150 = 10'h136 == r_count_9_io_out ? io_r_310_b : _GEN_7149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7151 = 10'h137 == r_count_9_io_out ? io_r_311_b : _GEN_7150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7152 = 10'h138 == r_count_9_io_out ? io_r_312_b : _GEN_7151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7153 = 10'h139 == r_count_9_io_out ? io_r_313_b : _GEN_7152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7154 = 10'h13a == r_count_9_io_out ? io_r_314_b : _GEN_7153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7155 = 10'h13b == r_count_9_io_out ? io_r_315_b : _GEN_7154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7156 = 10'h13c == r_count_9_io_out ? io_r_316_b : _GEN_7155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7157 = 10'h13d == r_count_9_io_out ? io_r_317_b : _GEN_7156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7158 = 10'h13e == r_count_9_io_out ? io_r_318_b : _GEN_7157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7159 = 10'h13f == r_count_9_io_out ? io_r_319_b : _GEN_7158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7160 = 10'h140 == r_count_9_io_out ? io_r_320_b : _GEN_7159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7161 = 10'h141 == r_count_9_io_out ? io_r_321_b : _GEN_7160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7162 = 10'h142 == r_count_9_io_out ? io_r_322_b : _GEN_7161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7163 = 10'h143 == r_count_9_io_out ? io_r_323_b : _GEN_7162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7164 = 10'h144 == r_count_9_io_out ? io_r_324_b : _GEN_7163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7165 = 10'h145 == r_count_9_io_out ? io_r_325_b : _GEN_7164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7166 = 10'h146 == r_count_9_io_out ? io_r_326_b : _GEN_7165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7167 = 10'h147 == r_count_9_io_out ? io_r_327_b : _GEN_7166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7168 = 10'h148 == r_count_9_io_out ? io_r_328_b : _GEN_7167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7169 = 10'h149 == r_count_9_io_out ? io_r_329_b : _GEN_7168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7170 = 10'h14a == r_count_9_io_out ? io_r_330_b : _GEN_7169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7171 = 10'h14b == r_count_9_io_out ? io_r_331_b : _GEN_7170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7172 = 10'h14c == r_count_9_io_out ? io_r_332_b : _GEN_7171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7173 = 10'h14d == r_count_9_io_out ? io_r_333_b : _GEN_7172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7174 = 10'h14e == r_count_9_io_out ? io_r_334_b : _GEN_7173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7175 = 10'h14f == r_count_9_io_out ? io_r_335_b : _GEN_7174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7176 = 10'h150 == r_count_9_io_out ? io_r_336_b : _GEN_7175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7177 = 10'h151 == r_count_9_io_out ? io_r_337_b : _GEN_7176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7178 = 10'h152 == r_count_9_io_out ? io_r_338_b : _GEN_7177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7179 = 10'h153 == r_count_9_io_out ? io_r_339_b : _GEN_7178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7180 = 10'h154 == r_count_9_io_out ? io_r_340_b : _GEN_7179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7181 = 10'h155 == r_count_9_io_out ? io_r_341_b : _GEN_7180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7182 = 10'h156 == r_count_9_io_out ? io_r_342_b : _GEN_7181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7183 = 10'h157 == r_count_9_io_out ? io_r_343_b : _GEN_7182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7184 = 10'h158 == r_count_9_io_out ? io_r_344_b : _GEN_7183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7185 = 10'h159 == r_count_9_io_out ? io_r_345_b : _GEN_7184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7186 = 10'h15a == r_count_9_io_out ? io_r_346_b : _GEN_7185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7187 = 10'h15b == r_count_9_io_out ? io_r_347_b : _GEN_7186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7188 = 10'h15c == r_count_9_io_out ? io_r_348_b : _GEN_7187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7189 = 10'h15d == r_count_9_io_out ? io_r_349_b : _GEN_7188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7190 = 10'h15e == r_count_9_io_out ? io_r_350_b : _GEN_7189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7191 = 10'h15f == r_count_9_io_out ? io_r_351_b : _GEN_7190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7192 = 10'h160 == r_count_9_io_out ? io_r_352_b : _GEN_7191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7193 = 10'h161 == r_count_9_io_out ? io_r_353_b : _GEN_7192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7194 = 10'h162 == r_count_9_io_out ? io_r_354_b : _GEN_7193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7195 = 10'h163 == r_count_9_io_out ? io_r_355_b : _GEN_7194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7196 = 10'h164 == r_count_9_io_out ? io_r_356_b : _GEN_7195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7197 = 10'h165 == r_count_9_io_out ? io_r_357_b : _GEN_7196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7198 = 10'h166 == r_count_9_io_out ? io_r_358_b : _GEN_7197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7199 = 10'h167 == r_count_9_io_out ? io_r_359_b : _GEN_7198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7200 = 10'h168 == r_count_9_io_out ? io_r_360_b : _GEN_7199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7201 = 10'h169 == r_count_9_io_out ? io_r_361_b : _GEN_7200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7202 = 10'h16a == r_count_9_io_out ? io_r_362_b : _GEN_7201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7203 = 10'h16b == r_count_9_io_out ? io_r_363_b : _GEN_7202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7204 = 10'h16c == r_count_9_io_out ? io_r_364_b : _GEN_7203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7205 = 10'h16d == r_count_9_io_out ? io_r_365_b : _GEN_7204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7206 = 10'h16e == r_count_9_io_out ? io_r_366_b : _GEN_7205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7207 = 10'h16f == r_count_9_io_out ? io_r_367_b : _GEN_7206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7208 = 10'h170 == r_count_9_io_out ? io_r_368_b : _GEN_7207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7209 = 10'h171 == r_count_9_io_out ? io_r_369_b : _GEN_7208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7210 = 10'h172 == r_count_9_io_out ? io_r_370_b : _GEN_7209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7211 = 10'h173 == r_count_9_io_out ? io_r_371_b : _GEN_7210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7212 = 10'h174 == r_count_9_io_out ? io_r_372_b : _GEN_7211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7213 = 10'h175 == r_count_9_io_out ? io_r_373_b : _GEN_7212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7214 = 10'h176 == r_count_9_io_out ? io_r_374_b : _GEN_7213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7215 = 10'h177 == r_count_9_io_out ? io_r_375_b : _GEN_7214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7216 = 10'h178 == r_count_9_io_out ? io_r_376_b : _GEN_7215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7217 = 10'h179 == r_count_9_io_out ? io_r_377_b : _GEN_7216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7218 = 10'h17a == r_count_9_io_out ? io_r_378_b : _GEN_7217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7219 = 10'h17b == r_count_9_io_out ? io_r_379_b : _GEN_7218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7220 = 10'h17c == r_count_9_io_out ? io_r_380_b : _GEN_7219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7221 = 10'h17d == r_count_9_io_out ? io_r_381_b : _GEN_7220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7222 = 10'h17e == r_count_9_io_out ? io_r_382_b : _GEN_7221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7223 = 10'h17f == r_count_9_io_out ? io_r_383_b : _GEN_7222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7224 = 10'h180 == r_count_9_io_out ? io_r_384_b : _GEN_7223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7225 = 10'h181 == r_count_9_io_out ? io_r_385_b : _GEN_7224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7226 = 10'h182 == r_count_9_io_out ? io_r_386_b : _GEN_7225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7227 = 10'h183 == r_count_9_io_out ? io_r_387_b : _GEN_7226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7228 = 10'h184 == r_count_9_io_out ? io_r_388_b : _GEN_7227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7229 = 10'h185 == r_count_9_io_out ? io_r_389_b : _GEN_7228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7230 = 10'h186 == r_count_9_io_out ? io_r_390_b : _GEN_7229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7231 = 10'h187 == r_count_9_io_out ? io_r_391_b : _GEN_7230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7232 = 10'h188 == r_count_9_io_out ? io_r_392_b : _GEN_7231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7233 = 10'h189 == r_count_9_io_out ? io_r_393_b : _GEN_7232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7234 = 10'h18a == r_count_9_io_out ? io_r_394_b : _GEN_7233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7235 = 10'h18b == r_count_9_io_out ? io_r_395_b : _GEN_7234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7236 = 10'h18c == r_count_9_io_out ? io_r_396_b : _GEN_7235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7237 = 10'h18d == r_count_9_io_out ? io_r_397_b : _GEN_7236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7238 = 10'h18e == r_count_9_io_out ? io_r_398_b : _GEN_7237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7239 = 10'h18f == r_count_9_io_out ? io_r_399_b : _GEN_7238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7240 = 10'h190 == r_count_9_io_out ? io_r_400_b : _GEN_7239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7241 = 10'h191 == r_count_9_io_out ? io_r_401_b : _GEN_7240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7242 = 10'h192 == r_count_9_io_out ? io_r_402_b : _GEN_7241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7243 = 10'h193 == r_count_9_io_out ? io_r_403_b : _GEN_7242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7244 = 10'h194 == r_count_9_io_out ? io_r_404_b : _GEN_7243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7245 = 10'h195 == r_count_9_io_out ? io_r_405_b : _GEN_7244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7246 = 10'h196 == r_count_9_io_out ? io_r_406_b : _GEN_7245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7247 = 10'h197 == r_count_9_io_out ? io_r_407_b : _GEN_7246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7248 = 10'h198 == r_count_9_io_out ? io_r_408_b : _GEN_7247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7249 = 10'h199 == r_count_9_io_out ? io_r_409_b : _GEN_7248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7250 = 10'h19a == r_count_9_io_out ? io_r_410_b : _GEN_7249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7251 = 10'h19b == r_count_9_io_out ? io_r_411_b : _GEN_7250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7252 = 10'h19c == r_count_9_io_out ? io_r_412_b : _GEN_7251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7253 = 10'h19d == r_count_9_io_out ? io_r_413_b : _GEN_7252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7254 = 10'h19e == r_count_9_io_out ? io_r_414_b : _GEN_7253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7255 = 10'h19f == r_count_9_io_out ? io_r_415_b : _GEN_7254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7256 = 10'h1a0 == r_count_9_io_out ? io_r_416_b : _GEN_7255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7257 = 10'h1a1 == r_count_9_io_out ? io_r_417_b : _GEN_7256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7258 = 10'h1a2 == r_count_9_io_out ? io_r_418_b : _GEN_7257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7259 = 10'h1a3 == r_count_9_io_out ? io_r_419_b : _GEN_7258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7260 = 10'h1a4 == r_count_9_io_out ? io_r_420_b : _GEN_7259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7261 = 10'h1a5 == r_count_9_io_out ? io_r_421_b : _GEN_7260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7262 = 10'h1a6 == r_count_9_io_out ? io_r_422_b : _GEN_7261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7263 = 10'h1a7 == r_count_9_io_out ? io_r_423_b : _GEN_7262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7264 = 10'h1a8 == r_count_9_io_out ? io_r_424_b : _GEN_7263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7265 = 10'h1a9 == r_count_9_io_out ? io_r_425_b : _GEN_7264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7266 = 10'h1aa == r_count_9_io_out ? io_r_426_b : _GEN_7265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7267 = 10'h1ab == r_count_9_io_out ? io_r_427_b : _GEN_7266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7268 = 10'h1ac == r_count_9_io_out ? io_r_428_b : _GEN_7267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7269 = 10'h1ad == r_count_9_io_out ? io_r_429_b : _GEN_7268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7270 = 10'h1ae == r_count_9_io_out ? io_r_430_b : _GEN_7269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7271 = 10'h1af == r_count_9_io_out ? io_r_431_b : _GEN_7270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7272 = 10'h1b0 == r_count_9_io_out ? io_r_432_b : _GEN_7271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7273 = 10'h1b1 == r_count_9_io_out ? io_r_433_b : _GEN_7272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7274 = 10'h1b2 == r_count_9_io_out ? io_r_434_b : _GEN_7273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7275 = 10'h1b3 == r_count_9_io_out ? io_r_435_b : _GEN_7274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7276 = 10'h1b4 == r_count_9_io_out ? io_r_436_b : _GEN_7275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7277 = 10'h1b5 == r_count_9_io_out ? io_r_437_b : _GEN_7276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7278 = 10'h1b6 == r_count_9_io_out ? io_r_438_b : _GEN_7277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7279 = 10'h1b7 == r_count_9_io_out ? io_r_439_b : _GEN_7278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7280 = 10'h1b8 == r_count_9_io_out ? io_r_440_b : _GEN_7279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7281 = 10'h1b9 == r_count_9_io_out ? io_r_441_b : _GEN_7280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7282 = 10'h1ba == r_count_9_io_out ? io_r_442_b : _GEN_7281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7283 = 10'h1bb == r_count_9_io_out ? io_r_443_b : _GEN_7282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7284 = 10'h1bc == r_count_9_io_out ? io_r_444_b : _GEN_7283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7285 = 10'h1bd == r_count_9_io_out ? io_r_445_b : _GEN_7284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7286 = 10'h1be == r_count_9_io_out ? io_r_446_b : _GEN_7285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7287 = 10'h1bf == r_count_9_io_out ? io_r_447_b : _GEN_7286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7288 = 10'h1c0 == r_count_9_io_out ? io_r_448_b : _GEN_7287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7289 = 10'h1c1 == r_count_9_io_out ? io_r_449_b : _GEN_7288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7290 = 10'h1c2 == r_count_9_io_out ? io_r_450_b : _GEN_7289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7291 = 10'h1c3 == r_count_9_io_out ? io_r_451_b : _GEN_7290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7292 = 10'h1c4 == r_count_9_io_out ? io_r_452_b : _GEN_7291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7293 = 10'h1c5 == r_count_9_io_out ? io_r_453_b : _GEN_7292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7294 = 10'h1c6 == r_count_9_io_out ? io_r_454_b : _GEN_7293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7295 = 10'h1c7 == r_count_9_io_out ? io_r_455_b : _GEN_7294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7296 = 10'h1c8 == r_count_9_io_out ? io_r_456_b : _GEN_7295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7297 = 10'h1c9 == r_count_9_io_out ? io_r_457_b : _GEN_7296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7298 = 10'h1ca == r_count_9_io_out ? io_r_458_b : _GEN_7297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7299 = 10'h1cb == r_count_9_io_out ? io_r_459_b : _GEN_7298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7300 = 10'h1cc == r_count_9_io_out ? io_r_460_b : _GEN_7299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7301 = 10'h1cd == r_count_9_io_out ? io_r_461_b : _GEN_7300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7302 = 10'h1ce == r_count_9_io_out ? io_r_462_b : _GEN_7301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7303 = 10'h1cf == r_count_9_io_out ? io_r_463_b : _GEN_7302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7304 = 10'h1d0 == r_count_9_io_out ? io_r_464_b : _GEN_7303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7305 = 10'h1d1 == r_count_9_io_out ? io_r_465_b : _GEN_7304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7306 = 10'h1d2 == r_count_9_io_out ? io_r_466_b : _GEN_7305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7307 = 10'h1d3 == r_count_9_io_out ? io_r_467_b : _GEN_7306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7308 = 10'h1d4 == r_count_9_io_out ? io_r_468_b : _GEN_7307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7309 = 10'h1d5 == r_count_9_io_out ? io_r_469_b : _GEN_7308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7310 = 10'h1d6 == r_count_9_io_out ? io_r_470_b : _GEN_7309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7311 = 10'h1d7 == r_count_9_io_out ? io_r_471_b : _GEN_7310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7312 = 10'h1d8 == r_count_9_io_out ? io_r_472_b : _GEN_7311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7313 = 10'h1d9 == r_count_9_io_out ? io_r_473_b : _GEN_7312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7314 = 10'h1da == r_count_9_io_out ? io_r_474_b : _GEN_7313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7315 = 10'h1db == r_count_9_io_out ? io_r_475_b : _GEN_7314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7316 = 10'h1dc == r_count_9_io_out ? io_r_476_b : _GEN_7315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7317 = 10'h1dd == r_count_9_io_out ? io_r_477_b : _GEN_7316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7318 = 10'h1de == r_count_9_io_out ? io_r_478_b : _GEN_7317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7319 = 10'h1df == r_count_9_io_out ? io_r_479_b : _GEN_7318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7320 = 10'h1e0 == r_count_9_io_out ? io_r_480_b : _GEN_7319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7321 = 10'h1e1 == r_count_9_io_out ? io_r_481_b : _GEN_7320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7322 = 10'h1e2 == r_count_9_io_out ? io_r_482_b : _GEN_7321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7323 = 10'h1e3 == r_count_9_io_out ? io_r_483_b : _GEN_7322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7324 = 10'h1e4 == r_count_9_io_out ? io_r_484_b : _GEN_7323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7325 = 10'h1e5 == r_count_9_io_out ? io_r_485_b : _GEN_7324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7326 = 10'h1e6 == r_count_9_io_out ? io_r_486_b : _GEN_7325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7327 = 10'h1e7 == r_count_9_io_out ? io_r_487_b : _GEN_7326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7328 = 10'h1e8 == r_count_9_io_out ? io_r_488_b : _GEN_7327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7329 = 10'h1e9 == r_count_9_io_out ? io_r_489_b : _GEN_7328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7330 = 10'h1ea == r_count_9_io_out ? io_r_490_b : _GEN_7329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7331 = 10'h1eb == r_count_9_io_out ? io_r_491_b : _GEN_7330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7332 = 10'h1ec == r_count_9_io_out ? io_r_492_b : _GEN_7331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7333 = 10'h1ed == r_count_9_io_out ? io_r_493_b : _GEN_7332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7334 = 10'h1ee == r_count_9_io_out ? io_r_494_b : _GEN_7333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7335 = 10'h1ef == r_count_9_io_out ? io_r_495_b : _GEN_7334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7336 = 10'h1f0 == r_count_9_io_out ? io_r_496_b : _GEN_7335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7337 = 10'h1f1 == r_count_9_io_out ? io_r_497_b : _GEN_7336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7338 = 10'h1f2 == r_count_9_io_out ? io_r_498_b : _GEN_7337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7339 = 10'h1f3 == r_count_9_io_out ? io_r_499_b : _GEN_7338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7340 = 10'h1f4 == r_count_9_io_out ? io_r_500_b : _GEN_7339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7341 = 10'h1f5 == r_count_9_io_out ? io_r_501_b : _GEN_7340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7342 = 10'h1f6 == r_count_9_io_out ? io_r_502_b : _GEN_7341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7343 = 10'h1f7 == r_count_9_io_out ? io_r_503_b : _GEN_7342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7344 = 10'h1f8 == r_count_9_io_out ? io_r_504_b : _GEN_7343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7345 = 10'h1f9 == r_count_9_io_out ? io_r_505_b : _GEN_7344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7346 = 10'h1fa == r_count_9_io_out ? io_r_506_b : _GEN_7345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7347 = 10'h1fb == r_count_9_io_out ? io_r_507_b : _GEN_7346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7348 = 10'h1fc == r_count_9_io_out ? io_r_508_b : _GEN_7347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7349 = 10'h1fd == r_count_9_io_out ? io_r_509_b : _GEN_7348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7350 = 10'h1fe == r_count_9_io_out ? io_r_510_b : _GEN_7349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7351 = 10'h1ff == r_count_9_io_out ? io_r_511_b : _GEN_7350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7352 = 10'h200 == r_count_9_io_out ? io_r_512_b : _GEN_7351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7353 = 10'h201 == r_count_9_io_out ? io_r_513_b : _GEN_7352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7354 = 10'h202 == r_count_9_io_out ? io_r_514_b : _GEN_7353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7355 = 10'h203 == r_count_9_io_out ? io_r_515_b : _GEN_7354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7356 = 10'h204 == r_count_9_io_out ? io_r_516_b : _GEN_7355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7357 = 10'h205 == r_count_9_io_out ? io_r_517_b : _GEN_7356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7358 = 10'h206 == r_count_9_io_out ? io_r_518_b : _GEN_7357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7359 = 10'h207 == r_count_9_io_out ? io_r_519_b : _GEN_7358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7360 = 10'h208 == r_count_9_io_out ? io_r_520_b : _GEN_7359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7361 = 10'h209 == r_count_9_io_out ? io_r_521_b : _GEN_7360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7362 = 10'h20a == r_count_9_io_out ? io_r_522_b : _GEN_7361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7363 = 10'h20b == r_count_9_io_out ? io_r_523_b : _GEN_7362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7364 = 10'h20c == r_count_9_io_out ? io_r_524_b : _GEN_7363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7365 = 10'h20d == r_count_9_io_out ? io_r_525_b : _GEN_7364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7366 = 10'h20e == r_count_9_io_out ? io_r_526_b : _GEN_7365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7367 = 10'h20f == r_count_9_io_out ? io_r_527_b : _GEN_7366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7368 = 10'h210 == r_count_9_io_out ? io_r_528_b : _GEN_7367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7369 = 10'h211 == r_count_9_io_out ? io_r_529_b : _GEN_7368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7370 = 10'h212 == r_count_9_io_out ? io_r_530_b : _GEN_7369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7371 = 10'h213 == r_count_9_io_out ? io_r_531_b : _GEN_7370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7372 = 10'h214 == r_count_9_io_out ? io_r_532_b : _GEN_7371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7373 = 10'h215 == r_count_9_io_out ? io_r_533_b : _GEN_7372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7374 = 10'h216 == r_count_9_io_out ? io_r_534_b : _GEN_7373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7375 = 10'h217 == r_count_9_io_out ? io_r_535_b : _GEN_7374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7376 = 10'h218 == r_count_9_io_out ? io_r_536_b : _GEN_7375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7377 = 10'h219 == r_count_9_io_out ? io_r_537_b : _GEN_7376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7378 = 10'h21a == r_count_9_io_out ? io_r_538_b : _GEN_7377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7379 = 10'h21b == r_count_9_io_out ? io_r_539_b : _GEN_7378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7380 = 10'h21c == r_count_9_io_out ? io_r_540_b : _GEN_7379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7381 = 10'h21d == r_count_9_io_out ? io_r_541_b : _GEN_7380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7382 = 10'h21e == r_count_9_io_out ? io_r_542_b : _GEN_7381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7383 = 10'h21f == r_count_9_io_out ? io_r_543_b : _GEN_7382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7384 = 10'h220 == r_count_9_io_out ? io_r_544_b : _GEN_7383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7385 = 10'h221 == r_count_9_io_out ? io_r_545_b : _GEN_7384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7386 = 10'h222 == r_count_9_io_out ? io_r_546_b : _GEN_7385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7387 = 10'h223 == r_count_9_io_out ? io_r_547_b : _GEN_7386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7388 = 10'h224 == r_count_9_io_out ? io_r_548_b : _GEN_7387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7389 = 10'h225 == r_count_9_io_out ? io_r_549_b : _GEN_7388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7390 = 10'h226 == r_count_9_io_out ? io_r_550_b : _GEN_7389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7391 = 10'h227 == r_count_9_io_out ? io_r_551_b : _GEN_7390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7392 = 10'h228 == r_count_9_io_out ? io_r_552_b : _GEN_7391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7393 = 10'h229 == r_count_9_io_out ? io_r_553_b : _GEN_7392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7394 = 10'h22a == r_count_9_io_out ? io_r_554_b : _GEN_7393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7395 = 10'h22b == r_count_9_io_out ? io_r_555_b : _GEN_7394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7396 = 10'h22c == r_count_9_io_out ? io_r_556_b : _GEN_7395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7397 = 10'h22d == r_count_9_io_out ? io_r_557_b : _GEN_7396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7398 = 10'h22e == r_count_9_io_out ? io_r_558_b : _GEN_7397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7399 = 10'h22f == r_count_9_io_out ? io_r_559_b : _GEN_7398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7400 = 10'h230 == r_count_9_io_out ? io_r_560_b : _GEN_7399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7401 = 10'h231 == r_count_9_io_out ? io_r_561_b : _GEN_7400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7402 = 10'h232 == r_count_9_io_out ? io_r_562_b : _GEN_7401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7403 = 10'h233 == r_count_9_io_out ? io_r_563_b : _GEN_7402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7404 = 10'h234 == r_count_9_io_out ? io_r_564_b : _GEN_7403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7405 = 10'h235 == r_count_9_io_out ? io_r_565_b : _GEN_7404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7406 = 10'h236 == r_count_9_io_out ? io_r_566_b : _GEN_7405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7407 = 10'h237 == r_count_9_io_out ? io_r_567_b : _GEN_7406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7408 = 10'h238 == r_count_9_io_out ? io_r_568_b : _GEN_7407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7409 = 10'h239 == r_count_9_io_out ? io_r_569_b : _GEN_7408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7410 = 10'h23a == r_count_9_io_out ? io_r_570_b : _GEN_7409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7411 = 10'h23b == r_count_9_io_out ? io_r_571_b : _GEN_7410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7412 = 10'h23c == r_count_9_io_out ? io_r_572_b : _GEN_7411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7413 = 10'h23d == r_count_9_io_out ? io_r_573_b : _GEN_7412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7414 = 10'h23e == r_count_9_io_out ? io_r_574_b : _GEN_7413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7415 = 10'h23f == r_count_9_io_out ? io_r_575_b : _GEN_7414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7416 = 10'h240 == r_count_9_io_out ? io_r_576_b : _GEN_7415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7417 = 10'h241 == r_count_9_io_out ? io_r_577_b : _GEN_7416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7418 = 10'h242 == r_count_9_io_out ? io_r_578_b : _GEN_7417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7419 = 10'h243 == r_count_9_io_out ? io_r_579_b : _GEN_7418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7420 = 10'h244 == r_count_9_io_out ? io_r_580_b : _GEN_7419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7421 = 10'h245 == r_count_9_io_out ? io_r_581_b : _GEN_7420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7422 = 10'h246 == r_count_9_io_out ? io_r_582_b : _GEN_7421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7423 = 10'h247 == r_count_9_io_out ? io_r_583_b : _GEN_7422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7424 = 10'h248 == r_count_9_io_out ? io_r_584_b : _GEN_7423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7425 = 10'h249 == r_count_9_io_out ? io_r_585_b : _GEN_7424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7426 = 10'h24a == r_count_9_io_out ? io_r_586_b : _GEN_7425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7427 = 10'h24b == r_count_9_io_out ? io_r_587_b : _GEN_7426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7428 = 10'h24c == r_count_9_io_out ? io_r_588_b : _GEN_7427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7429 = 10'h24d == r_count_9_io_out ? io_r_589_b : _GEN_7428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7430 = 10'h24e == r_count_9_io_out ? io_r_590_b : _GEN_7429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7431 = 10'h24f == r_count_9_io_out ? io_r_591_b : _GEN_7430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7432 = 10'h250 == r_count_9_io_out ? io_r_592_b : _GEN_7431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7433 = 10'h251 == r_count_9_io_out ? io_r_593_b : _GEN_7432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7434 = 10'h252 == r_count_9_io_out ? io_r_594_b : _GEN_7433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7435 = 10'h253 == r_count_9_io_out ? io_r_595_b : _GEN_7434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7436 = 10'h254 == r_count_9_io_out ? io_r_596_b : _GEN_7435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7437 = 10'h255 == r_count_9_io_out ? io_r_597_b : _GEN_7436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7438 = 10'h256 == r_count_9_io_out ? io_r_598_b : _GEN_7437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7439 = 10'h257 == r_count_9_io_out ? io_r_599_b : _GEN_7438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7440 = 10'h258 == r_count_9_io_out ? io_r_600_b : _GEN_7439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7441 = 10'h259 == r_count_9_io_out ? io_r_601_b : _GEN_7440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7442 = 10'h25a == r_count_9_io_out ? io_r_602_b : _GEN_7441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7443 = 10'h25b == r_count_9_io_out ? io_r_603_b : _GEN_7442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7444 = 10'h25c == r_count_9_io_out ? io_r_604_b : _GEN_7443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7445 = 10'h25d == r_count_9_io_out ? io_r_605_b : _GEN_7444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7446 = 10'h25e == r_count_9_io_out ? io_r_606_b : _GEN_7445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7447 = 10'h25f == r_count_9_io_out ? io_r_607_b : _GEN_7446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7448 = 10'h260 == r_count_9_io_out ? io_r_608_b : _GEN_7447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7449 = 10'h261 == r_count_9_io_out ? io_r_609_b : _GEN_7448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7450 = 10'h262 == r_count_9_io_out ? io_r_610_b : _GEN_7449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7451 = 10'h263 == r_count_9_io_out ? io_r_611_b : _GEN_7450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7452 = 10'h264 == r_count_9_io_out ? io_r_612_b : _GEN_7451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7453 = 10'h265 == r_count_9_io_out ? io_r_613_b : _GEN_7452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7454 = 10'h266 == r_count_9_io_out ? io_r_614_b : _GEN_7453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7455 = 10'h267 == r_count_9_io_out ? io_r_615_b : _GEN_7454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7456 = 10'h268 == r_count_9_io_out ? io_r_616_b : _GEN_7455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7457 = 10'h269 == r_count_9_io_out ? io_r_617_b : _GEN_7456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7458 = 10'h26a == r_count_9_io_out ? io_r_618_b : _GEN_7457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7459 = 10'h26b == r_count_9_io_out ? io_r_619_b : _GEN_7458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7460 = 10'h26c == r_count_9_io_out ? io_r_620_b : _GEN_7459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7461 = 10'h26d == r_count_9_io_out ? io_r_621_b : _GEN_7460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7462 = 10'h26e == r_count_9_io_out ? io_r_622_b : _GEN_7461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7463 = 10'h26f == r_count_9_io_out ? io_r_623_b : _GEN_7462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7464 = 10'h270 == r_count_9_io_out ? io_r_624_b : _GEN_7463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7465 = 10'h271 == r_count_9_io_out ? io_r_625_b : _GEN_7464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7466 = 10'h272 == r_count_9_io_out ? io_r_626_b : _GEN_7465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7467 = 10'h273 == r_count_9_io_out ? io_r_627_b : _GEN_7466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7468 = 10'h274 == r_count_9_io_out ? io_r_628_b : _GEN_7467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7469 = 10'h275 == r_count_9_io_out ? io_r_629_b : _GEN_7468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7470 = 10'h276 == r_count_9_io_out ? io_r_630_b : _GEN_7469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7471 = 10'h277 == r_count_9_io_out ? io_r_631_b : _GEN_7470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7472 = 10'h278 == r_count_9_io_out ? io_r_632_b : _GEN_7471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7473 = 10'h279 == r_count_9_io_out ? io_r_633_b : _GEN_7472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7474 = 10'h27a == r_count_9_io_out ? io_r_634_b : _GEN_7473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7475 = 10'h27b == r_count_9_io_out ? io_r_635_b : _GEN_7474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7476 = 10'h27c == r_count_9_io_out ? io_r_636_b : _GEN_7475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7477 = 10'h27d == r_count_9_io_out ? io_r_637_b : _GEN_7476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7478 = 10'h27e == r_count_9_io_out ? io_r_638_b : _GEN_7477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7479 = 10'h27f == r_count_9_io_out ? io_r_639_b : _GEN_7478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7480 = 10'h280 == r_count_9_io_out ? io_r_640_b : _GEN_7479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7481 = 10'h281 == r_count_9_io_out ? io_r_641_b : _GEN_7480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7482 = 10'h282 == r_count_9_io_out ? io_r_642_b : _GEN_7481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7483 = 10'h283 == r_count_9_io_out ? io_r_643_b : _GEN_7482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7484 = 10'h284 == r_count_9_io_out ? io_r_644_b : _GEN_7483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7485 = 10'h285 == r_count_9_io_out ? io_r_645_b : _GEN_7484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7486 = 10'h286 == r_count_9_io_out ? io_r_646_b : _GEN_7485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7487 = 10'h287 == r_count_9_io_out ? io_r_647_b : _GEN_7486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7488 = 10'h288 == r_count_9_io_out ? io_r_648_b : _GEN_7487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7489 = 10'h289 == r_count_9_io_out ? io_r_649_b : _GEN_7488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7490 = 10'h28a == r_count_9_io_out ? io_r_650_b : _GEN_7489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7491 = 10'h28b == r_count_9_io_out ? io_r_651_b : _GEN_7490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7492 = 10'h28c == r_count_9_io_out ? io_r_652_b : _GEN_7491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7493 = 10'h28d == r_count_9_io_out ? io_r_653_b : _GEN_7492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7494 = 10'h28e == r_count_9_io_out ? io_r_654_b : _GEN_7493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7495 = 10'h28f == r_count_9_io_out ? io_r_655_b : _GEN_7494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7496 = 10'h290 == r_count_9_io_out ? io_r_656_b : _GEN_7495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7497 = 10'h291 == r_count_9_io_out ? io_r_657_b : _GEN_7496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7498 = 10'h292 == r_count_9_io_out ? io_r_658_b : _GEN_7497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7499 = 10'h293 == r_count_9_io_out ? io_r_659_b : _GEN_7498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7500 = 10'h294 == r_count_9_io_out ? io_r_660_b : _GEN_7499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7501 = 10'h295 == r_count_9_io_out ? io_r_661_b : _GEN_7500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7502 = 10'h296 == r_count_9_io_out ? io_r_662_b : _GEN_7501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7503 = 10'h297 == r_count_9_io_out ? io_r_663_b : _GEN_7502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7504 = 10'h298 == r_count_9_io_out ? io_r_664_b : _GEN_7503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7505 = 10'h299 == r_count_9_io_out ? io_r_665_b : _GEN_7504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7506 = 10'h29a == r_count_9_io_out ? io_r_666_b : _GEN_7505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7507 = 10'h29b == r_count_9_io_out ? io_r_667_b : _GEN_7506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7508 = 10'h29c == r_count_9_io_out ? io_r_668_b : _GEN_7507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7509 = 10'h29d == r_count_9_io_out ? io_r_669_b : _GEN_7508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7510 = 10'h29e == r_count_9_io_out ? io_r_670_b : _GEN_7509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7511 = 10'h29f == r_count_9_io_out ? io_r_671_b : _GEN_7510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7512 = 10'h2a0 == r_count_9_io_out ? io_r_672_b : _GEN_7511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7513 = 10'h2a1 == r_count_9_io_out ? io_r_673_b : _GEN_7512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7514 = 10'h2a2 == r_count_9_io_out ? io_r_674_b : _GEN_7513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7515 = 10'h2a3 == r_count_9_io_out ? io_r_675_b : _GEN_7514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7516 = 10'h2a4 == r_count_9_io_out ? io_r_676_b : _GEN_7515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7517 = 10'h2a5 == r_count_9_io_out ? io_r_677_b : _GEN_7516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7518 = 10'h2a6 == r_count_9_io_out ? io_r_678_b : _GEN_7517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7519 = 10'h2a7 == r_count_9_io_out ? io_r_679_b : _GEN_7518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7520 = 10'h2a8 == r_count_9_io_out ? io_r_680_b : _GEN_7519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7521 = 10'h2a9 == r_count_9_io_out ? io_r_681_b : _GEN_7520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7522 = 10'h2aa == r_count_9_io_out ? io_r_682_b : _GEN_7521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7523 = 10'h2ab == r_count_9_io_out ? io_r_683_b : _GEN_7522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7524 = 10'h2ac == r_count_9_io_out ? io_r_684_b : _GEN_7523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7525 = 10'h2ad == r_count_9_io_out ? io_r_685_b : _GEN_7524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7526 = 10'h2ae == r_count_9_io_out ? io_r_686_b : _GEN_7525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7527 = 10'h2af == r_count_9_io_out ? io_r_687_b : _GEN_7526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7528 = 10'h2b0 == r_count_9_io_out ? io_r_688_b : _GEN_7527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7529 = 10'h2b1 == r_count_9_io_out ? io_r_689_b : _GEN_7528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7530 = 10'h2b2 == r_count_9_io_out ? io_r_690_b : _GEN_7529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7531 = 10'h2b3 == r_count_9_io_out ? io_r_691_b : _GEN_7530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7532 = 10'h2b4 == r_count_9_io_out ? io_r_692_b : _GEN_7531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7533 = 10'h2b5 == r_count_9_io_out ? io_r_693_b : _GEN_7532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7534 = 10'h2b6 == r_count_9_io_out ? io_r_694_b : _GEN_7533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7535 = 10'h2b7 == r_count_9_io_out ? io_r_695_b : _GEN_7534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7536 = 10'h2b8 == r_count_9_io_out ? io_r_696_b : _GEN_7535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7537 = 10'h2b9 == r_count_9_io_out ? io_r_697_b : _GEN_7536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7538 = 10'h2ba == r_count_9_io_out ? io_r_698_b : _GEN_7537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7539 = 10'h2bb == r_count_9_io_out ? io_r_699_b : _GEN_7538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7540 = 10'h2bc == r_count_9_io_out ? io_r_700_b : _GEN_7539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7541 = 10'h2bd == r_count_9_io_out ? io_r_701_b : _GEN_7540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7542 = 10'h2be == r_count_9_io_out ? io_r_702_b : _GEN_7541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7543 = 10'h2bf == r_count_9_io_out ? io_r_703_b : _GEN_7542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7544 = 10'h2c0 == r_count_9_io_out ? io_r_704_b : _GEN_7543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7545 = 10'h2c1 == r_count_9_io_out ? io_r_705_b : _GEN_7544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7546 = 10'h2c2 == r_count_9_io_out ? io_r_706_b : _GEN_7545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7547 = 10'h2c3 == r_count_9_io_out ? io_r_707_b : _GEN_7546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7548 = 10'h2c4 == r_count_9_io_out ? io_r_708_b : _GEN_7547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7549 = 10'h2c5 == r_count_9_io_out ? io_r_709_b : _GEN_7548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7550 = 10'h2c6 == r_count_9_io_out ? io_r_710_b : _GEN_7549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7551 = 10'h2c7 == r_count_9_io_out ? io_r_711_b : _GEN_7550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7552 = 10'h2c8 == r_count_9_io_out ? io_r_712_b : _GEN_7551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7553 = 10'h2c9 == r_count_9_io_out ? io_r_713_b : _GEN_7552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7554 = 10'h2ca == r_count_9_io_out ? io_r_714_b : _GEN_7553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7555 = 10'h2cb == r_count_9_io_out ? io_r_715_b : _GEN_7554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7556 = 10'h2cc == r_count_9_io_out ? io_r_716_b : _GEN_7555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7557 = 10'h2cd == r_count_9_io_out ? io_r_717_b : _GEN_7556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7558 = 10'h2ce == r_count_9_io_out ? io_r_718_b : _GEN_7557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7559 = 10'h2cf == r_count_9_io_out ? io_r_719_b : _GEN_7558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7560 = 10'h2d0 == r_count_9_io_out ? io_r_720_b : _GEN_7559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7561 = 10'h2d1 == r_count_9_io_out ? io_r_721_b : _GEN_7560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7562 = 10'h2d2 == r_count_9_io_out ? io_r_722_b : _GEN_7561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7563 = 10'h2d3 == r_count_9_io_out ? io_r_723_b : _GEN_7562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7564 = 10'h2d4 == r_count_9_io_out ? io_r_724_b : _GEN_7563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7565 = 10'h2d5 == r_count_9_io_out ? io_r_725_b : _GEN_7564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7566 = 10'h2d6 == r_count_9_io_out ? io_r_726_b : _GEN_7565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7567 = 10'h2d7 == r_count_9_io_out ? io_r_727_b : _GEN_7566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7568 = 10'h2d8 == r_count_9_io_out ? io_r_728_b : _GEN_7567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7569 = 10'h2d9 == r_count_9_io_out ? io_r_729_b : _GEN_7568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7570 = 10'h2da == r_count_9_io_out ? io_r_730_b : _GEN_7569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7571 = 10'h2db == r_count_9_io_out ? io_r_731_b : _GEN_7570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7572 = 10'h2dc == r_count_9_io_out ? io_r_732_b : _GEN_7571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7573 = 10'h2dd == r_count_9_io_out ? io_r_733_b : _GEN_7572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7574 = 10'h2de == r_count_9_io_out ? io_r_734_b : _GEN_7573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7575 = 10'h2df == r_count_9_io_out ? io_r_735_b : _GEN_7574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7576 = 10'h2e0 == r_count_9_io_out ? io_r_736_b : _GEN_7575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7577 = 10'h2e1 == r_count_9_io_out ? io_r_737_b : _GEN_7576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7578 = 10'h2e2 == r_count_9_io_out ? io_r_738_b : _GEN_7577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7579 = 10'h2e3 == r_count_9_io_out ? io_r_739_b : _GEN_7578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7580 = 10'h2e4 == r_count_9_io_out ? io_r_740_b : _GEN_7579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7581 = 10'h2e5 == r_count_9_io_out ? io_r_741_b : _GEN_7580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7582 = 10'h2e6 == r_count_9_io_out ? io_r_742_b : _GEN_7581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7583 = 10'h2e7 == r_count_9_io_out ? io_r_743_b : _GEN_7582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7584 = 10'h2e8 == r_count_9_io_out ? io_r_744_b : _GEN_7583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7585 = 10'h2e9 == r_count_9_io_out ? io_r_745_b : _GEN_7584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7586 = 10'h2ea == r_count_9_io_out ? io_r_746_b : _GEN_7585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7587 = 10'h2eb == r_count_9_io_out ? io_r_747_b : _GEN_7586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7588 = 10'h2ec == r_count_9_io_out ? io_r_748_b : _GEN_7587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7591 = 10'h1 == r_count_10_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7592 = 10'h2 == r_count_10_io_out ? io_r_2_b : _GEN_7591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7593 = 10'h3 == r_count_10_io_out ? io_r_3_b : _GEN_7592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7594 = 10'h4 == r_count_10_io_out ? io_r_4_b : _GEN_7593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7595 = 10'h5 == r_count_10_io_out ? io_r_5_b : _GEN_7594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7596 = 10'h6 == r_count_10_io_out ? io_r_6_b : _GEN_7595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7597 = 10'h7 == r_count_10_io_out ? io_r_7_b : _GEN_7596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7598 = 10'h8 == r_count_10_io_out ? io_r_8_b : _GEN_7597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7599 = 10'h9 == r_count_10_io_out ? io_r_9_b : _GEN_7598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7600 = 10'ha == r_count_10_io_out ? io_r_10_b : _GEN_7599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7601 = 10'hb == r_count_10_io_out ? io_r_11_b : _GEN_7600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7602 = 10'hc == r_count_10_io_out ? io_r_12_b : _GEN_7601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7603 = 10'hd == r_count_10_io_out ? io_r_13_b : _GEN_7602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7604 = 10'he == r_count_10_io_out ? io_r_14_b : _GEN_7603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7605 = 10'hf == r_count_10_io_out ? io_r_15_b : _GEN_7604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7606 = 10'h10 == r_count_10_io_out ? io_r_16_b : _GEN_7605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7607 = 10'h11 == r_count_10_io_out ? io_r_17_b : _GEN_7606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7608 = 10'h12 == r_count_10_io_out ? io_r_18_b : _GEN_7607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7609 = 10'h13 == r_count_10_io_out ? io_r_19_b : _GEN_7608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7610 = 10'h14 == r_count_10_io_out ? io_r_20_b : _GEN_7609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7611 = 10'h15 == r_count_10_io_out ? io_r_21_b : _GEN_7610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7612 = 10'h16 == r_count_10_io_out ? io_r_22_b : _GEN_7611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7613 = 10'h17 == r_count_10_io_out ? io_r_23_b : _GEN_7612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7614 = 10'h18 == r_count_10_io_out ? io_r_24_b : _GEN_7613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7615 = 10'h19 == r_count_10_io_out ? io_r_25_b : _GEN_7614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7616 = 10'h1a == r_count_10_io_out ? io_r_26_b : _GEN_7615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7617 = 10'h1b == r_count_10_io_out ? io_r_27_b : _GEN_7616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7618 = 10'h1c == r_count_10_io_out ? io_r_28_b : _GEN_7617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7619 = 10'h1d == r_count_10_io_out ? io_r_29_b : _GEN_7618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7620 = 10'h1e == r_count_10_io_out ? io_r_30_b : _GEN_7619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7621 = 10'h1f == r_count_10_io_out ? io_r_31_b : _GEN_7620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7622 = 10'h20 == r_count_10_io_out ? io_r_32_b : _GEN_7621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7623 = 10'h21 == r_count_10_io_out ? io_r_33_b : _GEN_7622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7624 = 10'h22 == r_count_10_io_out ? io_r_34_b : _GEN_7623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7625 = 10'h23 == r_count_10_io_out ? io_r_35_b : _GEN_7624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7626 = 10'h24 == r_count_10_io_out ? io_r_36_b : _GEN_7625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7627 = 10'h25 == r_count_10_io_out ? io_r_37_b : _GEN_7626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7628 = 10'h26 == r_count_10_io_out ? io_r_38_b : _GEN_7627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7629 = 10'h27 == r_count_10_io_out ? io_r_39_b : _GEN_7628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7630 = 10'h28 == r_count_10_io_out ? io_r_40_b : _GEN_7629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7631 = 10'h29 == r_count_10_io_out ? io_r_41_b : _GEN_7630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7632 = 10'h2a == r_count_10_io_out ? io_r_42_b : _GEN_7631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7633 = 10'h2b == r_count_10_io_out ? io_r_43_b : _GEN_7632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7634 = 10'h2c == r_count_10_io_out ? io_r_44_b : _GEN_7633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7635 = 10'h2d == r_count_10_io_out ? io_r_45_b : _GEN_7634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7636 = 10'h2e == r_count_10_io_out ? io_r_46_b : _GEN_7635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7637 = 10'h2f == r_count_10_io_out ? io_r_47_b : _GEN_7636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7638 = 10'h30 == r_count_10_io_out ? io_r_48_b : _GEN_7637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7639 = 10'h31 == r_count_10_io_out ? io_r_49_b : _GEN_7638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7640 = 10'h32 == r_count_10_io_out ? io_r_50_b : _GEN_7639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7641 = 10'h33 == r_count_10_io_out ? io_r_51_b : _GEN_7640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7642 = 10'h34 == r_count_10_io_out ? io_r_52_b : _GEN_7641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7643 = 10'h35 == r_count_10_io_out ? io_r_53_b : _GEN_7642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7644 = 10'h36 == r_count_10_io_out ? io_r_54_b : _GEN_7643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7645 = 10'h37 == r_count_10_io_out ? io_r_55_b : _GEN_7644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7646 = 10'h38 == r_count_10_io_out ? io_r_56_b : _GEN_7645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7647 = 10'h39 == r_count_10_io_out ? io_r_57_b : _GEN_7646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7648 = 10'h3a == r_count_10_io_out ? io_r_58_b : _GEN_7647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7649 = 10'h3b == r_count_10_io_out ? io_r_59_b : _GEN_7648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7650 = 10'h3c == r_count_10_io_out ? io_r_60_b : _GEN_7649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7651 = 10'h3d == r_count_10_io_out ? io_r_61_b : _GEN_7650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7652 = 10'h3e == r_count_10_io_out ? io_r_62_b : _GEN_7651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7653 = 10'h3f == r_count_10_io_out ? io_r_63_b : _GEN_7652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7654 = 10'h40 == r_count_10_io_out ? io_r_64_b : _GEN_7653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7655 = 10'h41 == r_count_10_io_out ? io_r_65_b : _GEN_7654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7656 = 10'h42 == r_count_10_io_out ? io_r_66_b : _GEN_7655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7657 = 10'h43 == r_count_10_io_out ? io_r_67_b : _GEN_7656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7658 = 10'h44 == r_count_10_io_out ? io_r_68_b : _GEN_7657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7659 = 10'h45 == r_count_10_io_out ? io_r_69_b : _GEN_7658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7660 = 10'h46 == r_count_10_io_out ? io_r_70_b : _GEN_7659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7661 = 10'h47 == r_count_10_io_out ? io_r_71_b : _GEN_7660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7662 = 10'h48 == r_count_10_io_out ? io_r_72_b : _GEN_7661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7663 = 10'h49 == r_count_10_io_out ? io_r_73_b : _GEN_7662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7664 = 10'h4a == r_count_10_io_out ? io_r_74_b : _GEN_7663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7665 = 10'h4b == r_count_10_io_out ? io_r_75_b : _GEN_7664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7666 = 10'h4c == r_count_10_io_out ? io_r_76_b : _GEN_7665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7667 = 10'h4d == r_count_10_io_out ? io_r_77_b : _GEN_7666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7668 = 10'h4e == r_count_10_io_out ? io_r_78_b : _GEN_7667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7669 = 10'h4f == r_count_10_io_out ? io_r_79_b : _GEN_7668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7670 = 10'h50 == r_count_10_io_out ? io_r_80_b : _GEN_7669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7671 = 10'h51 == r_count_10_io_out ? io_r_81_b : _GEN_7670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7672 = 10'h52 == r_count_10_io_out ? io_r_82_b : _GEN_7671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7673 = 10'h53 == r_count_10_io_out ? io_r_83_b : _GEN_7672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7674 = 10'h54 == r_count_10_io_out ? io_r_84_b : _GEN_7673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7675 = 10'h55 == r_count_10_io_out ? io_r_85_b : _GEN_7674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7676 = 10'h56 == r_count_10_io_out ? io_r_86_b : _GEN_7675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7677 = 10'h57 == r_count_10_io_out ? io_r_87_b : _GEN_7676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7678 = 10'h58 == r_count_10_io_out ? io_r_88_b : _GEN_7677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7679 = 10'h59 == r_count_10_io_out ? io_r_89_b : _GEN_7678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7680 = 10'h5a == r_count_10_io_out ? io_r_90_b : _GEN_7679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7681 = 10'h5b == r_count_10_io_out ? io_r_91_b : _GEN_7680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7682 = 10'h5c == r_count_10_io_out ? io_r_92_b : _GEN_7681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7683 = 10'h5d == r_count_10_io_out ? io_r_93_b : _GEN_7682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7684 = 10'h5e == r_count_10_io_out ? io_r_94_b : _GEN_7683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7685 = 10'h5f == r_count_10_io_out ? io_r_95_b : _GEN_7684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7686 = 10'h60 == r_count_10_io_out ? io_r_96_b : _GEN_7685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7687 = 10'h61 == r_count_10_io_out ? io_r_97_b : _GEN_7686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7688 = 10'h62 == r_count_10_io_out ? io_r_98_b : _GEN_7687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7689 = 10'h63 == r_count_10_io_out ? io_r_99_b : _GEN_7688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7690 = 10'h64 == r_count_10_io_out ? io_r_100_b : _GEN_7689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7691 = 10'h65 == r_count_10_io_out ? io_r_101_b : _GEN_7690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7692 = 10'h66 == r_count_10_io_out ? io_r_102_b : _GEN_7691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7693 = 10'h67 == r_count_10_io_out ? io_r_103_b : _GEN_7692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7694 = 10'h68 == r_count_10_io_out ? io_r_104_b : _GEN_7693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7695 = 10'h69 == r_count_10_io_out ? io_r_105_b : _GEN_7694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7696 = 10'h6a == r_count_10_io_out ? io_r_106_b : _GEN_7695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7697 = 10'h6b == r_count_10_io_out ? io_r_107_b : _GEN_7696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7698 = 10'h6c == r_count_10_io_out ? io_r_108_b : _GEN_7697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7699 = 10'h6d == r_count_10_io_out ? io_r_109_b : _GEN_7698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7700 = 10'h6e == r_count_10_io_out ? io_r_110_b : _GEN_7699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7701 = 10'h6f == r_count_10_io_out ? io_r_111_b : _GEN_7700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7702 = 10'h70 == r_count_10_io_out ? io_r_112_b : _GEN_7701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7703 = 10'h71 == r_count_10_io_out ? io_r_113_b : _GEN_7702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7704 = 10'h72 == r_count_10_io_out ? io_r_114_b : _GEN_7703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7705 = 10'h73 == r_count_10_io_out ? io_r_115_b : _GEN_7704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7706 = 10'h74 == r_count_10_io_out ? io_r_116_b : _GEN_7705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7707 = 10'h75 == r_count_10_io_out ? io_r_117_b : _GEN_7706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7708 = 10'h76 == r_count_10_io_out ? io_r_118_b : _GEN_7707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7709 = 10'h77 == r_count_10_io_out ? io_r_119_b : _GEN_7708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7710 = 10'h78 == r_count_10_io_out ? io_r_120_b : _GEN_7709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7711 = 10'h79 == r_count_10_io_out ? io_r_121_b : _GEN_7710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7712 = 10'h7a == r_count_10_io_out ? io_r_122_b : _GEN_7711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7713 = 10'h7b == r_count_10_io_out ? io_r_123_b : _GEN_7712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7714 = 10'h7c == r_count_10_io_out ? io_r_124_b : _GEN_7713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7715 = 10'h7d == r_count_10_io_out ? io_r_125_b : _GEN_7714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7716 = 10'h7e == r_count_10_io_out ? io_r_126_b : _GEN_7715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7717 = 10'h7f == r_count_10_io_out ? io_r_127_b : _GEN_7716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7718 = 10'h80 == r_count_10_io_out ? io_r_128_b : _GEN_7717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7719 = 10'h81 == r_count_10_io_out ? io_r_129_b : _GEN_7718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7720 = 10'h82 == r_count_10_io_out ? io_r_130_b : _GEN_7719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7721 = 10'h83 == r_count_10_io_out ? io_r_131_b : _GEN_7720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7722 = 10'h84 == r_count_10_io_out ? io_r_132_b : _GEN_7721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7723 = 10'h85 == r_count_10_io_out ? io_r_133_b : _GEN_7722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7724 = 10'h86 == r_count_10_io_out ? io_r_134_b : _GEN_7723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7725 = 10'h87 == r_count_10_io_out ? io_r_135_b : _GEN_7724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7726 = 10'h88 == r_count_10_io_out ? io_r_136_b : _GEN_7725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7727 = 10'h89 == r_count_10_io_out ? io_r_137_b : _GEN_7726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7728 = 10'h8a == r_count_10_io_out ? io_r_138_b : _GEN_7727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7729 = 10'h8b == r_count_10_io_out ? io_r_139_b : _GEN_7728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7730 = 10'h8c == r_count_10_io_out ? io_r_140_b : _GEN_7729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7731 = 10'h8d == r_count_10_io_out ? io_r_141_b : _GEN_7730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7732 = 10'h8e == r_count_10_io_out ? io_r_142_b : _GEN_7731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7733 = 10'h8f == r_count_10_io_out ? io_r_143_b : _GEN_7732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7734 = 10'h90 == r_count_10_io_out ? io_r_144_b : _GEN_7733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7735 = 10'h91 == r_count_10_io_out ? io_r_145_b : _GEN_7734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7736 = 10'h92 == r_count_10_io_out ? io_r_146_b : _GEN_7735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7737 = 10'h93 == r_count_10_io_out ? io_r_147_b : _GEN_7736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7738 = 10'h94 == r_count_10_io_out ? io_r_148_b : _GEN_7737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7739 = 10'h95 == r_count_10_io_out ? io_r_149_b : _GEN_7738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7740 = 10'h96 == r_count_10_io_out ? io_r_150_b : _GEN_7739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7741 = 10'h97 == r_count_10_io_out ? io_r_151_b : _GEN_7740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7742 = 10'h98 == r_count_10_io_out ? io_r_152_b : _GEN_7741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7743 = 10'h99 == r_count_10_io_out ? io_r_153_b : _GEN_7742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7744 = 10'h9a == r_count_10_io_out ? io_r_154_b : _GEN_7743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7745 = 10'h9b == r_count_10_io_out ? io_r_155_b : _GEN_7744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7746 = 10'h9c == r_count_10_io_out ? io_r_156_b : _GEN_7745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7747 = 10'h9d == r_count_10_io_out ? io_r_157_b : _GEN_7746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7748 = 10'h9e == r_count_10_io_out ? io_r_158_b : _GEN_7747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7749 = 10'h9f == r_count_10_io_out ? io_r_159_b : _GEN_7748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7750 = 10'ha0 == r_count_10_io_out ? io_r_160_b : _GEN_7749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7751 = 10'ha1 == r_count_10_io_out ? io_r_161_b : _GEN_7750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7752 = 10'ha2 == r_count_10_io_out ? io_r_162_b : _GEN_7751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7753 = 10'ha3 == r_count_10_io_out ? io_r_163_b : _GEN_7752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7754 = 10'ha4 == r_count_10_io_out ? io_r_164_b : _GEN_7753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7755 = 10'ha5 == r_count_10_io_out ? io_r_165_b : _GEN_7754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7756 = 10'ha6 == r_count_10_io_out ? io_r_166_b : _GEN_7755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7757 = 10'ha7 == r_count_10_io_out ? io_r_167_b : _GEN_7756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7758 = 10'ha8 == r_count_10_io_out ? io_r_168_b : _GEN_7757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7759 = 10'ha9 == r_count_10_io_out ? io_r_169_b : _GEN_7758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7760 = 10'haa == r_count_10_io_out ? io_r_170_b : _GEN_7759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7761 = 10'hab == r_count_10_io_out ? io_r_171_b : _GEN_7760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7762 = 10'hac == r_count_10_io_out ? io_r_172_b : _GEN_7761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7763 = 10'had == r_count_10_io_out ? io_r_173_b : _GEN_7762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7764 = 10'hae == r_count_10_io_out ? io_r_174_b : _GEN_7763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7765 = 10'haf == r_count_10_io_out ? io_r_175_b : _GEN_7764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7766 = 10'hb0 == r_count_10_io_out ? io_r_176_b : _GEN_7765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7767 = 10'hb1 == r_count_10_io_out ? io_r_177_b : _GEN_7766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7768 = 10'hb2 == r_count_10_io_out ? io_r_178_b : _GEN_7767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7769 = 10'hb3 == r_count_10_io_out ? io_r_179_b : _GEN_7768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7770 = 10'hb4 == r_count_10_io_out ? io_r_180_b : _GEN_7769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7771 = 10'hb5 == r_count_10_io_out ? io_r_181_b : _GEN_7770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7772 = 10'hb6 == r_count_10_io_out ? io_r_182_b : _GEN_7771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7773 = 10'hb7 == r_count_10_io_out ? io_r_183_b : _GEN_7772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7774 = 10'hb8 == r_count_10_io_out ? io_r_184_b : _GEN_7773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7775 = 10'hb9 == r_count_10_io_out ? io_r_185_b : _GEN_7774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7776 = 10'hba == r_count_10_io_out ? io_r_186_b : _GEN_7775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7777 = 10'hbb == r_count_10_io_out ? io_r_187_b : _GEN_7776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7778 = 10'hbc == r_count_10_io_out ? io_r_188_b : _GEN_7777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7779 = 10'hbd == r_count_10_io_out ? io_r_189_b : _GEN_7778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7780 = 10'hbe == r_count_10_io_out ? io_r_190_b : _GEN_7779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7781 = 10'hbf == r_count_10_io_out ? io_r_191_b : _GEN_7780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7782 = 10'hc0 == r_count_10_io_out ? io_r_192_b : _GEN_7781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7783 = 10'hc1 == r_count_10_io_out ? io_r_193_b : _GEN_7782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7784 = 10'hc2 == r_count_10_io_out ? io_r_194_b : _GEN_7783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7785 = 10'hc3 == r_count_10_io_out ? io_r_195_b : _GEN_7784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7786 = 10'hc4 == r_count_10_io_out ? io_r_196_b : _GEN_7785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7787 = 10'hc5 == r_count_10_io_out ? io_r_197_b : _GEN_7786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7788 = 10'hc6 == r_count_10_io_out ? io_r_198_b : _GEN_7787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7789 = 10'hc7 == r_count_10_io_out ? io_r_199_b : _GEN_7788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7790 = 10'hc8 == r_count_10_io_out ? io_r_200_b : _GEN_7789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7791 = 10'hc9 == r_count_10_io_out ? io_r_201_b : _GEN_7790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7792 = 10'hca == r_count_10_io_out ? io_r_202_b : _GEN_7791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7793 = 10'hcb == r_count_10_io_out ? io_r_203_b : _GEN_7792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7794 = 10'hcc == r_count_10_io_out ? io_r_204_b : _GEN_7793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7795 = 10'hcd == r_count_10_io_out ? io_r_205_b : _GEN_7794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7796 = 10'hce == r_count_10_io_out ? io_r_206_b : _GEN_7795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7797 = 10'hcf == r_count_10_io_out ? io_r_207_b : _GEN_7796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7798 = 10'hd0 == r_count_10_io_out ? io_r_208_b : _GEN_7797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7799 = 10'hd1 == r_count_10_io_out ? io_r_209_b : _GEN_7798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7800 = 10'hd2 == r_count_10_io_out ? io_r_210_b : _GEN_7799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7801 = 10'hd3 == r_count_10_io_out ? io_r_211_b : _GEN_7800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7802 = 10'hd4 == r_count_10_io_out ? io_r_212_b : _GEN_7801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7803 = 10'hd5 == r_count_10_io_out ? io_r_213_b : _GEN_7802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7804 = 10'hd6 == r_count_10_io_out ? io_r_214_b : _GEN_7803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7805 = 10'hd7 == r_count_10_io_out ? io_r_215_b : _GEN_7804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7806 = 10'hd8 == r_count_10_io_out ? io_r_216_b : _GEN_7805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7807 = 10'hd9 == r_count_10_io_out ? io_r_217_b : _GEN_7806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7808 = 10'hda == r_count_10_io_out ? io_r_218_b : _GEN_7807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7809 = 10'hdb == r_count_10_io_out ? io_r_219_b : _GEN_7808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7810 = 10'hdc == r_count_10_io_out ? io_r_220_b : _GEN_7809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7811 = 10'hdd == r_count_10_io_out ? io_r_221_b : _GEN_7810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7812 = 10'hde == r_count_10_io_out ? io_r_222_b : _GEN_7811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7813 = 10'hdf == r_count_10_io_out ? io_r_223_b : _GEN_7812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7814 = 10'he0 == r_count_10_io_out ? io_r_224_b : _GEN_7813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7815 = 10'he1 == r_count_10_io_out ? io_r_225_b : _GEN_7814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7816 = 10'he2 == r_count_10_io_out ? io_r_226_b : _GEN_7815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7817 = 10'he3 == r_count_10_io_out ? io_r_227_b : _GEN_7816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7818 = 10'he4 == r_count_10_io_out ? io_r_228_b : _GEN_7817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7819 = 10'he5 == r_count_10_io_out ? io_r_229_b : _GEN_7818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7820 = 10'he6 == r_count_10_io_out ? io_r_230_b : _GEN_7819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7821 = 10'he7 == r_count_10_io_out ? io_r_231_b : _GEN_7820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7822 = 10'he8 == r_count_10_io_out ? io_r_232_b : _GEN_7821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7823 = 10'he9 == r_count_10_io_out ? io_r_233_b : _GEN_7822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7824 = 10'hea == r_count_10_io_out ? io_r_234_b : _GEN_7823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7825 = 10'heb == r_count_10_io_out ? io_r_235_b : _GEN_7824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7826 = 10'hec == r_count_10_io_out ? io_r_236_b : _GEN_7825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7827 = 10'hed == r_count_10_io_out ? io_r_237_b : _GEN_7826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7828 = 10'hee == r_count_10_io_out ? io_r_238_b : _GEN_7827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7829 = 10'hef == r_count_10_io_out ? io_r_239_b : _GEN_7828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7830 = 10'hf0 == r_count_10_io_out ? io_r_240_b : _GEN_7829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7831 = 10'hf1 == r_count_10_io_out ? io_r_241_b : _GEN_7830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7832 = 10'hf2 == r_count_10_io_out ? io_r_242_b : _GEN_7831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7833 = 10'hf3 == r_count_10_io_out ? io_r_243_b : _GEN_7832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7834 = 10'hf4 == r_count_10_io_out ? io_r_244_b : _GEN_7833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7835 = 10'hf5 == r_count_10_io_out ? io_r_245_b : _GEN_7834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7836 = 10'hf6 == r_count_10_io_out ? io_r_246_b : _GEN_7835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7837 = 10'hf7 == r_count_10_io_out ? io_r_247_b : _GEN_7836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7838 = 10'hf8 == r_count_10_io_out ? io_r_248_b : _GEN_7837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7839 = 10'hf9 == r_count_10_io_out ? io_r_249_b : _GEN_7838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7840 = 10'hfa == r_count_10_io_out ? io_r_250_b : _GEN_7839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7841 = 10'hfb == r_count_10_io_out ? io_r_251_b : _GEN_7840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7842 = 10'hfc == r_count_10_io_out ? io_r_252_b : _GEN_7841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7843 = 10'hfd == r_count_10_io_out ? io_r_253_b : _GEN_7842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7844 = 10'hfe == r_count_10_io_out ? io_r_254_b : _GEN_7843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7845 = 10'hff == r_count_10_io_out ? io_r_255_b : _GEN_7844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7846 = 10'h100 == r_count_10_io_out ? io_r_256_b : _GEN_7845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7847 = 10'h101 == r_count_10_io_out ? io_r_257_b : _GEN_7846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7848 = 10'h102 == r_count_10_io_out ? io_r_258_b : _GEN_7847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7849 = 10'h103 == r_count_10_io_out ? io_r_259_b : _GEN_7848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7850 = 10'h104 == r_count_10_io_out ? io_r_260_b : _GEN_7849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7851 = 10'h105 == r_count_10_io_out ? io_r_261_b : _GEN_7850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7852 = 10'h106 == r_count_10_io_out ? io_r_262_b : _GEN_7851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7853 = 10'h107 == r_count_10_io_out ? io_r_263_b : _GEN_7852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7854 = 10'h108 == r_count_10_io_out ? io_r_264_b : _GEN_7853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7855 = 10'h109 == r_count_10_io_out ? io_r_265_b : _GEN_7854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7856 = 10'h10a == r_count_10_io_out ? io_r_266_b : _GEN_7855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7857 = 10'h10b == r_count_10_io_out ? io_r_267_b : _GEN_7856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7858 = 10'h10c == r_count_10_io_out ? io_r_268_b : _GEN_7857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7859 = 10'h10d == r_count_10_io_out ? io_r_269_b : _GEN_7858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7860 = 10'h10e == r_count_10_io_out ? io_r_270_b : _GEN_7859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7861 = 10'h10f == r_count_10_io_out ? io_r_271_b : _GEN_7860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7862 = 10'h110 == r_count_10_io_out ? io_r_272_b : _GEN_7861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7863 = 10'h111 == r_count_10_io_out ? io_r_273_b : _GEN_7862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7864 = 10'h112 == r_count_10_io_out ? io_r_274_b : _GEN_7863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7865 = 10'h113 == r_count_10_io_out ? io_r_275_b : _GEN_7864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7866 = 10'h114 == r_count_10_io_out ? io_r_276_b : _GEN_7865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7867 = 10'h115 == r_count_10_io_out ? io_r_277_b : _GEN_7866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7868 = 10'h116 == r_count_10_io_out ? io_r_278_b : _GEN_7867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7869 = 10'h117 == r_count_10_io_out ? io_r_279_b : _GEN_7868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7870 = 10'h118 == r_count_10_io_out ? io_r_280_b : _GEN_7869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7871 = 10'h119 == r_count_10_io_out ? io_r_281_b : _GEN_7870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7872 = 10'h11a == r_count_10_io_out ? io_r_282_b : _GEN_7871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7873 = 10'h11b == r_count_10_io_out ? io_r_283_b : _GEN_7872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7874 = 10'h11c == r_count_10_io_out ? io_r_284_b : _GEN_7873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7875 = 10'h11d == r_count_10_io_out ? io_r_285_b : _GEN_7874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7876 = 10'h11e == r_count_10_io_out ? io_r_286_b : _GEN_7875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7877 = 10'h11f == r_count_10_io_out ? io_r_287_b : _GEN_7876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7878 = 10'h120 == r_count_10_io_out ? io_r_288_b : _GEN_7877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7879 = 10'h121 == r_count_10_io_out ? io_r_289_b : _GEN_7878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7880 = 10'h122 == r_count_10_io_out ? io_r_290_b : _GEN_7879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7881 = 10'h123 == r_count_10_io_out ? io_r_291_b : _GEN_7880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7882 = 10'h124 == r_count_10_io_out ? io_r_292_b : _GEN_7881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7883 = 10'h125 == r_count_10_io_out ? io_r_293_b : _GEN_7882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7884 = 10'h126 == r_count_10_io_out ? io_r_294_b : _GEN_7883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7885 = 10'h127 == r_count_10_io_out ? io_r_295_b : _GEN_7884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7886 = 10'h128 == r_count_10_io_out ? io_r_296_b : _GEN_7885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7887 = 10'h129 == r_count_10_io_out ? io_r_297_b : _GEN_7886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7888 = 10'h12a == r_count_10_io_out ? io_r_298_b : _GEN_7887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7889 = 10'h12b == r_count_10_io_out ? io_r_299_b : _GEN_7888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7890 = 10'h12c == r_count_10_io_out ? io_r_300_b : _GEN_7889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7891 = 10'h12d == r_count_10_io_out ? io_r_301_b : _GEN_7890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7892 = 10'h12e == r_count_10_io_out ? io_r_302_b : _GEN_7891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7893 = 10'h12f == r_count_10_io_out ? io_r_303_b : _GEN_7892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7894 = 10'h130 == r_count_10_io_out ? io_r_304_b : _GEN_7893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7895 = 10'h131 == r_count_10_io_out ? io_r_305_b : _GEN_7894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7896 = 10'h132 == r_count_10_io_out ? io_r_306_b : _GEN_7895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7897 = 10'h133 == r_count_10_io_out ? io_r_307_b : _GEN_7896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7898 = 10'h134 == r_count_10_io_out ? io_r_308_b : _GEN_7897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7899 = 10'h135 == r_count_10_io_out ? io_r_309_b : _GEN_7898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7900 = 10'h136 == r_count_10_io_out ? io_r_310_b : _GEN_7899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7901 = 10'h137 == r_count_10_io_out ? io_r_311_b : _GEN_7900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7902 = 10'h138 == r_count_10_io_out ? io_r_312_b : _GEN_7901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7903 = 10'h139 == r_count_10_io_out ? io_r_313_b : _GEN_7902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7904 = 10'h13a == r_count_10_io_out ? io_r_314_b : _GEN_7903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7905 = 10'h13b == r_count_10_io_out ? io_r_315_b : _GEN_7904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7906 = 10'h13c == r_count_10_io_out ? io_r_316_b : _GEN_7905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7907 = 10'h13d == r_count_10_io_out ? io_r_317_b : _GEN_7906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7908 = 10'h13e == r_count_10_io_out ? io_r_318_b : _GEN_7907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7909 = 10'h13f == r_count_10_io_out ? io_r_319_b : _GEN_7908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7910 = 10'h140 == r_count_10_io_out ? io_r_320_b : _GEN_7909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7911 = 10'h141 == r_count_10_io_out ? io_r_321_b : _GEN_7910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7912 = 10'h142 == r_count_10_io_out ? io_r_322_b : _GEN_7911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7913 = 10'h143 == r_count_10_io_out ? io_r_323_b : _GEN_7912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7914 = 10'h144 == r_count_10_io_out ? io_r_324_b : _GEN_7913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7915 = 10'h145 == r_count_10_io_out ? io_r_325_b : _GEN_7914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7916 = 10'h146 == r_count_10_io_out ? io_r_326_b : _GEN_7915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7917 = 10'h147 == r_count_10_io_out ? io_r_327_b : _GEN_7916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7918 = 10'h148 == r_count_10_io_out ? io_r_328_b : _GEN_7917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7919 = 10'h149 == r_count_10_io_out ? io_r_329_b : _GEN_7918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7920 = 10'h14a == r_count_10_io_out ? io_r_330_b : _GEN_7919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7921 = 10'h14b == r_count_10_io_out ? io_r_331_b : _GEN_7920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7922 = 10'h14c == r_count_10_io_out ? io_r_332_b : _GEN_7921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7923 = 10'h14d == r_count_10_io_out ? io_r_333_b : _GEN_7922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7924 = 10'h14e == r_count_10_io_out ? io_r_334_b : _GEN_7923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7925 = 10'h14f == r_count_10_io_out ? io_r_335_b : _GEN_7924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7926 = 10'h150 == r_count_10_io_out ? io_r_336_b : _GEN_7925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7927 = 10'h151 == r_count_10_io_out ? io_r_337_b : _GEN_7926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7928 = 10'h152 == r_count_10_io_out ? io_r_338_b : _GEN_7927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7929 = 10'h153 == r_count_10_io_out ? io_r_339_b : _GEN_7928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7930 = 10'h154 == r_count_10_io_out ? io_r_340_b : _GEN_7929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7931 = 10'h155 == r_count_10_io_out ? io_r_341_b : _GEN_7930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7932 = 10'h156 == r_count_10_io_out ? io_r_342_b : _GEN_7931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7933 = 10'h157 == r_count_10_io_out ? io_r_343_b : _GEN_7932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7934 = 10'h158 == r_count_10_io_out ? io_r_344_b : _GEN_7933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7935 = 10'h159 == r_count_10_io_out ? io_r_345_b : _GEN_7934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7936 = 10'h15a == r_count_10_io_out ? io_r_346_b : _GEN_7935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7937 = 10'h15b == r_count_10_io_out ? io_r_347_b : _GEN_7936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7938 = 10'h15c == r_count_10_io_out ? io_r_348_b : _GEN_7937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7939 = 10'h15d == r_count_10_io_out ? io_r_349_b : _GEN_7938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7940 = 10'h15e == r_count_10_io_out ? io_r_350_b : _GEN_7939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7941 = 10'h15f == r_count_10_io_out ? io_r_351_b : _GEN_7940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7942 = 10'h160 == r_count_10_io_out ? io_r_352_b : _GEN_7941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7943 = 10'h161 == r_count_10_io_out ? io_r_353_b : _GEN_7942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7944 = 10'h162 == r_count_10_io_out ? io_r_354_b : _GEN_7943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7945 = 10'h163 == r_count_10_io_out ? io_r_355_b : _GEN_7944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7946 = 10'h164 == r_count_10_io_out ? io_r_356_b : _GEN_7945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7947 = 10'h165 == r_count_10_io_out ? io_r_357_b : _GEN_7946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7948 = 10'h166 == r_count_10_io_out ? io_r_358_b : _GEN_7947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7949 = 10'h167 == r_count_10_io_out ? io_r_359_b : _GEN_7948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7950 = 10'h168 == r_count_10_io_out ? io_r_360_b : _GEN_7949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7951 = 10'h169 == r_count_10_io_out ? io_r_361_b : _GEN_7950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7952 = 10'h16a == r_count_10_io_out ? io_r_362_b : _GEN_7951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7953 = 10'h16b == r_count_10_io_out ? io_r_363_b : _GEN_7952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7954 = 10'h16c == r_count_10_io_out ? io_r_364_b : _GEN_7953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7955 = 10'h16d == r_count_10_io_out ? io_r_365_b : _GEN_7954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7956 = 10'h16e == r_count_10_io_out ? io_r_366_b : _GEN_7955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7957 = 10'h16f == r_count_10_io_out ? io_r_367_b : _GEN_7956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7958 = 10'h170 == r_count_10_io_out ? io_r_368_b : _GEN_7957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7959 = 10'h171 == r_count_10_io_out ? io_r_369_b : _GEN_7958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7960 = 10'h172 == r_count_10_io_out ? io_r_370_b : _GEN_7959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7961 = 10'h173 == r_count_10_io_out ? io_r_371_b : _GEN_7960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7962 = 10'h174 == r_count_10_io_out ? io_r_372_b : _GEN_7961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7963 = 10'h175 == r_count_10_io_out ? io_r_373_b : _GEN_7962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7964 = 10'h176 == r_count_10_io_out ? io_r_374_b : _GEN_7963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7965 = 10'h177 == r_count_10_io_out ? io_r_375_b : _GEN_7964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7966 = 10'h178 == r_count_10_io_out ? io_r_376_b : _GEN_7965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7967 = 10'h179 == r_count_10_io_out ? io_r_377_b : _GEN_7966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7968 = 10'h17a == r_count_10_io_out ? io_r_378_b : _GEN_7967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7969 = 10'h17b == r_count_10_io_out ? io_r_379_b : _GEN_7968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7970 = 10'h17c == r_count_10_io_out ? io_r_380_b : _GEN_7969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7971 = 10'h17d == r_count_10_io_out ? io_r_381_b : _GEN_7970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7972 = 10'h17e == r_count_10_io_out ? io_r_382_b : _GEN_7971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7973 = 10'h17f == r_count_10_io_out ? io_r_383_b : _GEN_7972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7974 = 10'h180 == r_count_10_io_out ? io_r_384_b : _GEN_7973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7975 = 10'h181 == r_count_10_io_out ? io_r_385_b : _GEN_7974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7976 = 10'h182 == r_count_10_io_out ? io_r_386_b : _GEN_7975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7977 = 10'h183 == r_count_10_io_out ? io_r_387_b : _GEN_7976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7978 = 10'h184 == r_count_10_io_out ? io_r_388_b : _GEN_7977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7979 = 10'h185 == r_count_10_io_out ? io_r_389_b : _GEN_7978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7980 = 10'h186 == r_count_10_io_out ? io_r_390_b : _GEN_7979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7981 = 10'h187 == r_count_10_io_out ? io_r_391_b : _GEN_7980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7982 = 10'h188 == r_count_10_io_out ? io_r_392_b : _GEN_7981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7983 = 10'h189 == r_count_10_io_out ? io_r_393_b : _GEN_7982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7984 = 10'h18a == r_count_10_io_out ? io_r_394_b : _GEN_7983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7985 = 10'h18b == r_count_10_io_out ? io_r_395_b : _GEN_7984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7986 = 10'h18c == r_count_10_io_out ? io_r_396_b : _GEN_7985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7987 = 10'h18d == r_count_10_io_out ? io_r_397_b : _GEN_7986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7988 = 10'h18e == r_count_10_io_out ? io_r_398_b : _GEN_7987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7989 = 10'h18f == r_count_10_io_out ? io_r_399_b : _GEN_7988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7990 = 10'h190 == r_count_10_io_out ? io_r_400_b : _GEN_7989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7991 = 10'h191 == r_count_10_io_out ? io_r_401_b : _GEN_7990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7992 = 10'h192 == r_count_10_io_out ? io_r_402_b : _GEN_7991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7993 = 10'h193 == r_count_10_io_out ? io_r_403_b : _GEN_7992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7994 = 10'h194 == r_count_10_io_out ? io_r_404_b : _GEN_7993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7995 = 10'h195 == r_count_10_io_out ? io_r_405_b : _GEN_7994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7996 = 10'h196 == r_count_10_io_out ? io_r_406_b : _GEN_7995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7997 = 10'h197 == r_count_10_io_out ? io_r_407_b : _GEN_7996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7998 = 10'h198 == r_count_10_io_out ? io_r_408_b : _GEN_7997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7999 = 10'h199 == r_count_10_io_out ? io_r_409_b : _GEN_7998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8000 = 10'h19a == r_count_10_io_out ? io_r_410_b : _GEN_7999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8001 = 10'h19b == r_count_10_io_out ? io_r_411_b : _GEN_8000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8002 = 10'h19c == r_count_10_io_out ? io_r_412_b : _GEN_8001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8003 = 10'h19d == r_count_10_io_out ? io_r_413_b : _GEN_8002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8004 = 10'h19e == r_count_10_io_out ? io_r_414_b : _GEN_8003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8005 = 10'h19f == r_count_10_io_out ? io_r_415_b : _GEN_8004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8006 = 10'h1a0 == r_count_10_io_out ? io_r_416_b : _GEN_8005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8007 = 10'h1a1 == r_count_10_io_out ? io_r_417_b : _GEN_8006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8008 = 10'h1a2 == r_count_10_io_out ? io_r_418_b : _GEN_8007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8009 = 10'h1a3 == r_count_10_io_out ? io_r_419_b : _GEN_8008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8010 = 10'h1a4 == r_count_10_io_out ? io_r_420_b : _GEN_8009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8011 = 10'h1a5 == r_count_10_io_out ? io_r_421_b : _GEN_8010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8012 = 10'h1a6 == r_count_10_io_out ? io_r_422_b : _GEN_8011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8013 = 10'h1a7 == r_count_10_io_out ? io_r_423_b : _GEN_8012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8014 = 10'h1a8 == r_count_10_io_out ? io_r_424_b : _GEN_8013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8015 = 10'h1a9 == r_count_10_io_out ? io_r_425_b : _GEN_8014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8016 = 10'h1aa == r_count_10_io_out ? io_r_426_b : _GEN_8015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8017 = 10'h1ab == r_count_10_io_out ? io_r_427_b : _GEN_8016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8018 = 10'h1ac == r_count_10_io_out ? io_r_428_b : _GEN_8017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8019 = 10'h1ad == r_count_10_io_out ? io_r_429_b : _GEN_8018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8020 = 10'h1ae == r_count_10_io_out ? io_r_430_b : _GEN_8019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8021 = 10'h1af == r_count_10_io_out ? io_r_431_b : _GEN_8020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8022 = 10'h1b0 == r_count_10_io_out ? io_r_432_b : _GEN_8021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8023 = 10'h1b1 == r_count_10_io_out ? io_r_433_b : _GEN_8022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8024 = 10'h1b2 == r_count_10_io_out ? io_r_434_b : _GEN_8023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8025 = 10'h1b3 == r_count_10_io_out ? io_r_435_b : _GEN_8024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8026 = 10'h1b4 == r_count_10_io_out ? io_r_436_b : _GEN_8025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8027 = 10'h1b5 == r_count_10_io_out ? io_r_437_b : _GEN_8026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8028 = 10'h1b6 == r_count_10_io_out ? io_r_438_b : _GEN_8027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8029 = 10'h1b7 == r_count_10_io_out ? io_r_439_b : _GEN_8028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8030 = 10'h1b8 == r_count_10_io_out ? io_r_440_b : _GEN_8029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8031 = 10'h1b9 == r_count_10_io_out ? io_r_441_b : _GEN_8030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8032 = 10'h1ba == r_count_10_io_out ? io_r_442_b : _GEN_8031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8033 = 10'h1bb == r_count_10_io_out ? io_r_443_b : _GEN_8032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8034 = 10'h1bc == r_count_10_io_out ? io_r_444_b : _GEN_8033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8035 = 10'h1bd == r_count_10_io_out ? io_r_445_b : _GEN_8034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8036 = 10'h1be == r_count_10_io_out ? io_r_446_b : _GEN_8035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8037 = 10'h1bf == r_count_10_io_out ? io_r_447_b : _GEN_8036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8038 = 10'h1c0 == r_count_10_io_out ? io_r_448_b : _GEN_8037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8039 = 10'h1c1 == r_count_10_io_out ? io_r_449_b : _GEN_8038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8040 = 10'h1c2 == r_count_10_io_out ? io_r_450_b : _GEN_8039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8041 = 10'h1c3 == r_count_10_io_out ? io_r_451_b : _GEN_8040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8042 = 10'h1c4 == r_count_10_io_out ? io_r_452_b : _GEN_8041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8043 = 10'h1c5 == r_count_10_io_out ? io_r_453_b : _GEN_8042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8044 = 10'h1c6 == r_count_10_io_out ? io_r_454_b : _GEN_8043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8045 = 10'h1c7 == r_count_10_io_out ? io_r_455_b : _GEN_8044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8046 = 10'h1c8 == r_count_10_io_out ? io_r_456_b : _GEN_8045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8047 = 10'h1c9 == r_count_10_io_out ? io_r_457_b : _GEN_8046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8048 = 10'h1ca == r_count_10_io_out ? io_r_458_b : _GEN_8047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8049 = 10'h1cb == r_count_10_io_out ? io_r_459_b : _GEN_8048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8050 = 10'h1cc == r_count_10_io_out ? io_r_460_b : _GEN_8049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8051 = 10'h1cd == r_count_10_io_out ? io_r_461_b : _GEN_8050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8052 = 10'h1ce == r_count_10_io_out ? io_r_462_b : _GEN_8051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8053 = 10'h1cf == r_count_10_io_out ? io_r_463_b : _GEN_8052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8054 = 10'h1d0 == r_count_10_io_out ? io_r_464_b : _GEN_8053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8055 = 10'h1d1 == r_count_10_io_out ? io_r_465_b : _GEN_8054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8056 = 10'h1d2 == r_count_10_io_out ? io_r_466_b : _GEN_8055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8057 = 10'h1d3 == r_count_10_io_out ? io_r_467_b : _GEN_8056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8058 = 10'h1d4 == r_count_10_io_out ? io_r_468_b : _GEN_8057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8059 = 10'h1d5 == r_count_10_io_out ? io_r_469_b : _GEN_8058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8060 = 10'h1d6 == r_count_10_io_out ? io_r_470_b : _GEN_8059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8061 = 10'h1d7 == r_count_10_io_out ? io_r_471_b : _GEN_8060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8062 = 10'h1d8 == r_count_10_io_out ? io_r_472_b : _GEN_8061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8063 = 10'h1d9 == r_count_10_io_out ? io_r_473_b : _GEN_8062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8064 = 10'h1da == r_count_10_io_out ? io_r_474_b : _GEN_8063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8065 = 10'h1db == r_count_10_io_out ? io_r_475_b : _GEN_8064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8066 = 10'h1dc == r_count_10_io_out ? io_r_476_b : _GEN_8065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8067 = 10'h1dd == r_count_10_io_out ? io_r_477_b : _GEN_8066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8068 = 10'h1de == r_count_10_io_out ? io_r_478_b : _GEN_8067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8069 = 10'h1df == r_count_10_io_out ? io_r_479_b : _GEN_8068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8070 = 10'h1e0 == r_count_10_io_out ? io_r_480_b : _GEN_8069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8071 = 10'h1e1 == r_count_10_io_out ? io_r_481_b : _GEN_8070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8072 = 10'h1e2 == r_count_10_io_out ? io_r_482_b : _GEN_8071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8073 = 10'h1e3 == r_count_10_io_out ? io_r_483_b : _GEN_8072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8074 = 10'h1e4 == r_count_10_io_out ? io_r_484_b : _GEN_8073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8075 = 10'h1e5 == r_count_10_io_out ? io_r_485_b : _GEN_8074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8076 = 10'h1e6 == r_count_10_io_out ? io_r_486_b : _GEN_8075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8077 = 10'h1e7 == r_count_10_io_out ? io_r_487_b : _GEN_8076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8078 = 10'h1e8 == r_count_10_io_out ? io_r_488_b : _GEN_8077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8079 = 10'h1e9 == r_count_10_io_out ? io_r_489_b : _GEN_8078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8080 = 10'h1ea == r_count_10_io_out ? io_r_490_b : _GEN_8079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8081 = 10'h1eb == r_count_10_io_out ? io_r_491_b : _GEN_8080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8082 = 10'h1ec == r_count_10_io_out ? io_r_492_b : _GEN_8081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8083 = 10'h1ed == r_count_10_io_out ? io_r_493_b : _GEN_8082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8084 = 10'h1ee == r_count_10_io_out ? io_r_494_b : _GEN_8083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8085 = 10'h1ef == r_count_10_io_out ? io_r_495_b : _GEN_8084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8086 = 10'h1f0 == r_count_10_io_out ? io_r_496_b : _GEN_8085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8087 = 10'h1f1 == r_count_10_io_out ? io_r_497_b : _GEN_8086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8088 = 10'h1f2 == r_count_10_io_out ? io_r_498_b : _GEN_8087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8089 = 10'h1f3 == r_count_10_io_out ? io_r_499_b : _GEN_8088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8090 = 10'h1f4 == r_count_10_io_out ? io_r_500_b : _GEN_8089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8091 = 10'h1f5 == r_count_10_io_out ? io_r_501_b : _GEN_8090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8092 = 10'h1f6 == r_count_10_io_out ? io_r_502_b : _GEN_8091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8093 = 10'h1f7 == r_count_10_io_out ? io_r_503_b : _GEN_8092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8094 = 10'h1f8 == r_count_10_io_out ? io_r_504_b : _GEN_8093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8095 = 10'h1f9 == r_count_10_io_out ? io_r_505_b : _GEN_8094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8096 = 10'h1fa == r_count_10_io_out ? io_r_506_b : _GEN_8095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8097 = 10'h1fb == r_count_10_io_out ? io_r_507_b : _GEN_8096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8098 = 10'h1fc == r_count_10_io_out ? io_r_508_b : _GEN_8097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8099 = 10'h1fd == r_count_10_io_out ? io_r_509_b : _GEN_8098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8100 = 10'h1fe == r_count_10_io_out ? io_r_510_b : _GEN_8099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8101 = 10'h1ff == r_count_10_io_out ? io_r_511_b : _GEN_8100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8102 = 10'h200 == r_count_10_io_out ? io_r_512_b : _GEN_8101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8103 = 10'h201 == r_count_10_io_out ? io_r_513_b : _GEN_8102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8104 = 10'h202 == r_count_10_io_out ? io_r_514_b : _GEN_8103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8105 = 10'h203 == r_count_10_io_out ? io_r_515_b : _GEN_8104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8106 = 10'h204 == r_count_10_io_out ? io_r_516_b : _GEN_8105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8107 = 10'h205 == r_count_10_io_out ? io_r_517_b : _GEN_8106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8108 = 10'h206 == r_count_10_io_out ? io_r_518_b : _GEN_8107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8109 = 10'h207 == r_count_10_io_out ? io_r_519_b : _GEN_8108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8110 = 10'h208 == r_count_10_io_out ? io_r_520_b : _GEN_8109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8111 = 10'h209 == r_count_10_io_out ? io_r_521_b : _GEN_8110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8112 = 10'h20a == r_count_10_io_out ? io_r_522_b : _GEN_8111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8113 = 10'h20b == r_count_10_io_out ? io_r_523_b : _GEN_8112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8114 = 10'h20c == r_count_10_io_out ? io_r_524_b : _GEN_8113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8115 = 10'h20d == r_count_10_io_out ? io_r_525_b : _GEN_8114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8116 = 10'h20e == r_count_10_io_out ? io_r_526_b : _GEN_8115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8117 = 10'h20f == r_count_10_io_out ? io_r_527_b : _GEN_8116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8118 = 10'h210 == r_count_10_io_out ? io_r_528_b : _GEN_8117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8119 = 10'h211 == r_count_10_io_out ? io_r_529_b : _GEN_8118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8120 = 10'h212 == r_count_10_io_out ? io_r_530_b : _GEN_8119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8121 = 10'h213 == r_count_10_io_out ? io_r_531_b : _GEN_8120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8122 = 10'h214 == r_count_10_io_out ? io_r_532_b : _GEN_8121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8123 = 10'h215 == r_count_10_io_out ? io_r_533_b : _GEN_8122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8124 = 10'h216 == r_count_10_io_out ? io_r_534_b : _GEN_8123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8125 = 10'h217 == r_count_10_io_out ? io_r_535_b : _GEN_8124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8126 = 10'h218 == r_count_10_io_out ? io_r_536_b : _GEN_8125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8127 = 10'h219 == r_count_10_io_out ? io_r_537_b : _GEN_8126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8128 = 10'h21a == r_count_10_io_out ? io_r_538_b : _GEN_8127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8129 = 10'h21b == r_count_10_io_out ? io_r_539_b : _GEN_8128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8130 = 10'h21c == r_count_10_io_out ? io_r_540_b : _GEN_8129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8131 = 10'h21d == r_count_10_io_out ? io_r_541_b : _GEN_8130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8132 = 10'h21e == r_count_10_io_out ? io_r_542_b : _GEN_8131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8133 = 10'h21f == r_count_10_io_out ? io_r_543_b : _GEN_8132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8134 = 10'h220 == r_count_10_io_out ? io_r_544_b : _GEN_8133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8135 = 10'h221 == r_count_10_io_out ? io_r_545_b : _GEN_8134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8136 = 10'h222 == r_count_10_io_out ? io_r_546_b : _GEN_8135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8137 = 10'h223 == r_count_10_io_out ? io_r_547_b : _GEN_8136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8138 = 10'h224 == r_count_10_io_out ? io_r_548_b : _GEN_8137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8139 = 10'h225 == r_count_10_io_out ? io_r_549_b : _GEN_8138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8140 = 10'h226 == r_count_10_io_out ? io_r_550_b : _GEN_8139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8141 = 10'h227 == r_count_10_io_out ? io_r_551_b : _GEN_8140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8142 = 10'h228 == r_count_10_io_out ? io_r_552_b : _GEN_8141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8143 = 10'h229 == r_count_10_io_out ? io_r_553_b : _GEN_8142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8144 = 10'h22a == r_count_10_io_out ? io_r_554_b : _GEN_8143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8145 = 10'h22b == r_count_10_io_out ? io_r_555_b : _GEN_8144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8146 = 10'h22c == r_count_10_io_out ? io_r_556_b : _GEN_8145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8147 = 10'h22d == r_count_10_io_out ? io_r_557_b : _GEN_8146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8148 = 10'h22e == r_count_10_io_out ? io_r_558_b : _GEN_8147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8149 = 10'h22f == r_count_10_io_out ? io_r_559_b : _GEN_8148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8150 = 10'h230 == r_count_10_io_out ? io_r_560_b : _GEN_8149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8151 = 10'h231 == r_count_10_io_out ? io_r_561_b : _GEN_8150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8152 = 10'h232 == r_count_10_io_out ? io_r_562_b : _GEN_8151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8153 = 10'h233 == r_count_10_io_out ? io_r_563_b : _GEN_8152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8154 = 10'h234 == r_count_10_io_out ? io_r_564_b : _GEN_8153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8155 = 10'h235 == r_count_10_io_out ? io_r_565_b : _GEN_8154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8156 = 10'h236 == r_count_10_io_out ? io_r_566_b : _GEN_8155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8157 = 10'h237 == r_count_10_io_out ? io_r_567_b : _GEN_8156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8158 = 10'h238 == r_count_10_io_out ? io_r_568_b : _GEN_8157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8159 = 10'h239 == r_count_10_io_out ? io_r_569_b : _GEN_8158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8160 = 10'h23a == r_count_10_io_out ? io_r_570_b : _GEN_8159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8161 = 10'h23b == r_count_10_io_out ? io_r_571_b : _GEN_8160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8162 = 10'h23c == r_count_10_io_out ? io_r_572_b : _GEN_8161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8163 = 10'h23d == r_count_10_io_out ? io_r_573_b : _GEN_8162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8164 = 10'h23e == r_count_10_io_out ? io_r_574_b : _GEN_8163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8165 = 10'h23f == r_count_10_io_out ? io_r_575_b : _GEN_8164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8166 = 10'h240 == r_count_10_io_out ? io_r_576_b : _GEN_8165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8167 = 10'h241 == r_count_10_io_out ? io_r_577_b : _GEN_8166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8168 = 10'h242 == r_count_10_io_out ? io_r_578_b : _GEN_8167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8169 = 10'h243 == r_count_10_io_out ? io_r_579_b : _GEN_8168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8170 = 10'h244 == r_count_10_io_out ? io_r_580_b : _GEN_8169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8171 = 10'h245 == r_count_10_io_out ? io_r_581_b : _GEN_8170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8172 = 10'h246 == r_count_10_io_out ? io_r_582_b : _GEN_8171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8173 = 10'h247 == r_count_10_io_out ? io_r_583_b : _GEN_8172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8174 = 10'h248 == r_count_10_io_out ? io_r_584_b : _GEN_8173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8175 = 10'h249 == r_count_10_io_out ? io_r_585_b : _GEN_8174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8176 = 10'h24a == r_count_10_io_out ? io_r_586_b : _GEN_8175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8177 = 10'h24b == r_count_10_io_out ? io_r_587_b : _GEN_8176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8178 = 10'h24c == r_count_10_io_out ? io_r_588_b : _GEN_8177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8179 = 10'h24d == r_count_10_io_out ? io_r_589_b : _GEN_8178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8180 = 10'h24e == r_count_10_io_out ? io_r_590_b : _GEN_8179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8181 = 10'h24f == r_count_10_io_out ? io_r_591_b : _GEN_8180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8182 = 10'h250 == r_count_10_io_out ? io_r_592_b : _GEN_8181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8183 = 10'h251 == r_count_10_io_out ? io_r_593_b : _GEN_8182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8184 = 10'h252 == r_count_10_io_out ? io_r_594_b : _GEN_8183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8185 = 10'h253 == r_count_10_io_out ? io_r_595_b : _GEN_8184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8186 = 10'h254 == r_count_10_io_out ? io_r_596_b : _GEN_8185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8187 = 10'h255 == r_count_10_io_out ? io_r_597_b : _GEN_8186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8188 = 10'h256 == r_count_10_io_out ? io_r_598_b : _GEN_8187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8189 = 10'h257 == r_count_10_io_out ? io_r_599_b : _GEN_8188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8190 = 10'h258 == r_count_10_io_out ? io_r_600_b : _GEN_8189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8191 = 10'h259 == r_count_10_io_out ? io_r_601_b : _GEN_8190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8192 = 10'h25a == r_count_10_io_out ? io_r_602_b : _GEN_8191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8193 = 10'h25b == r_count_10_io_out ? io_r_603_b : _GEN_8192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8194 = 10'h25c == r_count_10_io_out ? io_r_604_b : _GEN_8193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8195 = 10'h25d == r_count_10_io_out ? io_r_605_b : _GEN_8194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8196 = 10'h25e == r_count_10_io_out ? io_r_606_b : _GEN_8195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8197 = 10'h25f == r_count_10_io_out ? io_r_607_b : _GEN_8196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8198 = 10'h260 == r_count_10_io_out ? io_r_608_b : _GEN_8197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8199 = 10'h261 == r_count_10_io_out ? io_r_609_b : _GEN_8198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8200 = 10'h262 == r_count_10_io_out ? io_r_610_b : _GEN_8199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8201 = 10'h263 == r_count_10_io_out ? io_r_611_b : _GEN_8200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8202 = 10'h264 == r_count_10_io_out ? io_r_612_b : _GEN_8201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8203 = 10'h265 == r_count_10_io_out ? io_r_613_b : _GEN_8202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8204 = 10'h266 == r_count_10_io_out ? io_r_614_b : _GEN_8203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8205 = 10'h267 == r_count_10_io_out ? io_r_615_b : _GEN_8204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8206 = 10'h268 == r_count_10_io_out ? io_r_616_b : _GEN_8205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8207 = 10'h269 == r_count_10_io_out ? io_r_617_b : _GEN_8206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8208 = 10'h26a == r_count_10_io_out ? io_r_618_b : _GEN_8207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8209 = 10'h26b == r_count_10_io_out ? io_r_619_b : _GEN_8208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8210 = 10'h26c == r_count_10_io_out ? io_r_620_b : _GEN_8209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8211 = 10'h26d == r_count_10_io_out ? io_r_621_b : _GEN_8210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8212 = 10'h26e == r_count_10_io_out ? io_r_622_b : _GEN_8211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8213 = 10'h26f == r_count_10_io_out ? io_r_623_b : _GEN_8212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8214 = 10'h270 == r_count_10_io_out ? io_r_624_b : _GEN_8213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8215 = 10'h271 == r_count_10_io_out ? io_r_625_b : _GEN_8214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8216 = 10'h272 == r_count_10_io_out ? io_r_626_b : _GEN_8215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8217 = 10'h273 == r_count_10_io_out ? io_r_627_b : _GEN_8216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8218 = 10'h274 == r_count_10_io_out ? io_r_628_b : _GEN_8217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8219 = 10'h275 == r_count_10_io_out ? io_r_629_b : _GEN_8218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8220 = 10'h276 == r_count_10_io_out ? io_r_630_b : _GEN_8219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8221 = 10'h277 == r_count_10_io_out ? io_r_631_b : _GEN_8220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8222 = 10'h278 == r_count_10_io_out ? io_r_632_b : _GEN_8221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8223 = 10'h279 == r_count_10_io_out ? io_r_633_b : _GEN_8222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8224 = 10'h27a == r_count_10_io_out ? io_r_634_b : _GEN_8223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8225 = 10'h27b == r_count_10_io_out ? io_r_635_b : _GEN_8224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8226 = 10'h27c == r_count_10_io_out ? io_r_636_b : _GEN_8225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8227 = 10'h27d == r_count_10_io_out ? io_r_637_b : _GEN_8226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8228 = 10'h27e == r_count_10_io_out ? io_r_638_b : _GEN_8227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8229 = 10'h27f == r_count_10_io_out ? io_r_639_b : _GEN_8228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8230 = 10'h280 == r_count_10_io_out ? io_r_640_b : _GEN_8229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8231 = 10'h281 == r_count_10_io_out ? io_r_641_b : _GEN_8230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8232 = 10'h282 == r_count_10_io_out ? io_r_642_b : _GEN_8231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8233 = 10'h283 == r_count_10_io_out ? io_r_643_b : _GEN_8232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8234 = 10'h284 == r_count_10_io_out ? io_r_644_b : _GEN_8233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8235 = 10'h285 == r_count_10_io_out ? io_r_645_b : _GEN_8234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8236 = 10'h286 == r_count_10_io_out ? io_r_646_b : _GEN_8235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8237 = 10'h287 == r_count_10_io_out ? io_r_647_b : _GEN_8236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8238 = 10'h288 == r_count_10_io_out ? io_r_648_b : _GEN_8237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8239 = 10'h289 == r_count_10_io_out ? io_r_649_b : _GEN_8238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8240 = 10'h28a == r_count_10_io_out ? io_r_650_b : _GEN_8239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8241 = 10'h28b == r_count_10_io_out ? io_r_651_b : _GEN_8240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8242 = 10'h28c == r_count_10_io_out ? io_r_652_b : _GEN_8241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8243 = 10'h28d == r_count_10_io_out ? io_r_653_b : _GEN_8242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8244 = 10'h28e == r_count_10_io_out ? io_r_654_b : _GEN_8243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8245 = 10'h28f == r_count_10_io_out ? io_r_655_b : _GEN_8244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8246 = 10'h290 == r_count_10_io_out ? io_r_656_b : _GEN_8245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8247 = 10'h291 == r_count_10_io_out ? io_r_657_b : _GEN_8246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8248 = 10'h292 == r_count_10_io_out ? io_r_658_b : _GEN_8247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8249 = 10'h293 == r_count_10_io_out ? io_r_659_b : _GEN_8248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8250 = 10'h294 == r_count_10_io_out ? io_r_660_b : _GEN_8249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8251 = 10'h295 == r_count_10_io_out ? io_r_661_b : _GEN_8250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8252 = 10'h296 == r_count_10_io_out ? io_r_662_b : _GEN_8251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8253 = 10'h297 == r_count_10_io_out ? io_r_663_b : _GEN_8252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8254 = 10'h298 == r_count_10_io_out ? io_r_664_b : _GEN_8253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8255 = 10'h299 == r_count_10_io_out ? io_r_665_b : _GEN_8254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8256 = 10'h29a == r_count_10_io_out ? io_r_666_b : _GEN_8255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8257 = 10'h29b == r_count_10_io_out ? io_r_667_b : _GEN_8256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8258 = 10'h29c == r_count_10_io_out ? io_r_668_b : _GEN_8257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8259 = 10'h29d == r_count_10_io_out ? io_r_669_b : _GEN_8258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8260 = 10'h29e == r_count_10_io_out ? io_r_670_b : _GEN_8259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8261 = 10'h29f == r_count_10_io_out ? io_r_671_b : _GEN_8260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8262 = 10'h2a0 == r_count_10_io_out ? io_r_672_b : _GEN_8261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8263 = 10'h2a1 == r_count_10_io_out ? io_r_673_b : _GEN_8262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8264 = 10'h2a2 == r_count_10_io_out ? io_r_674_b : _GEN_8263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8265 = 10'h2a3 == r_count_10_io_out ? io_r_675_b : _GEN_8264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8266 = 10'h2a4 == r_count_10_io_out ? io_r_676_b : _GEN_8265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8267 = 10'h2a5 == r_count_10_io_out ? io_r_677_b : _GEN_8266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8268 = 10'h2a6 == r_count_10_io_out ? io_r_678_b : _GEN_8267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8269 = 10'h2a7 == r_count_10_io_out ? io_r_679_b : _GEN_8268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8270 = 10'h2a8 == r_count_10_io_out ? io_r_680_b : _GEN_8269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8271 = 10'h2a9 == r_count_10_io_out ? io_r_681_b : _GEN_8270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8272 = 10'h2aa == r_count_10_io_out ? io_r_682_b : _GEN_8271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8273 = 10'h2ab == r_count_10_io_out ? io_r_683_b : _GEN_8272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8274 = 10'h2ac == r_count_10_io_out ? io_r_684_b : _GEN_8273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8275 = 10'h2ad == r_count_10_io_out ? io_r_685_b : _GEN_8274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8276 = 10'h2ae == r_count_10_io_out ? io_r_686_b : _GEN_8275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8277 = 10'h2af == r_count_10_io_out ? io_r_687_b : _GEN_8276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8278 = 10'h2b0 == r_count_10_io_out ? io_r_688_b : _GEN_8277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8279 = 10'h2b1 == r_count_10_io_out ? io_r_689_b : _GEN_8278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8280 = 10'h2b2 == r_count_10_io_out ? io_r_690_b : _GEN_8279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8281 = 10'h2b3 == r_count_10_io_out ? io_r_691_b : _GEN_8280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8282 = 10'h2b4 == r_count_10_io_out ? io_r_692_b : _GEN_8281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8283 = 10'h2b5 == r_count_10_io_out ? io_r_693_b : _GEN_8282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8284 = 10'h2b6 == r_count_10_io_out ? io_r_694_b : _GEN_8283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8285 = 10'h2b7 == r_count_10_io_out ? io_r_695_b : _GEN_8284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8286 = 10'h2b8 == r_count_10_io_out ? io_r_696_b : _GEN_8285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8287 = 10'h2b9 == r_count_10_io_out ? io_r_697_b : _GEN_8286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8288 = 10'h2ba == r_count_10_io_out ? io_r_698_b : _GEN_8287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8289 = 10'h2bb == r_count_10_io_out ? io_r_699_b : _GEN_8288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8290 = 10'h2bc == r_count_10_io_out ? io_r_700_b : _GEN_8289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8291 = 10'h2bd == r_count_10_io_out ? io_r_701_b : _GEN_8290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8292 = 10'h2be == r_count_10_io_out ? io_r_702_b : _GEN_8291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8293 = 10'h2bf == r_count_10_io_out ? io_r_703_b : _GEN_8292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8294 = 10'h2c0 == r_count_10_io_out ? io_r_704_b : _GEN_8293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8295 = 10'h2c1 == r_count_10_io_out ? io_r_705_b : _GEN_8294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8296 = 10'h2c2 == r_count_10_io_out ? io_r_706_b : _GEN_8295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8297 = 10'h2c3 == r_count_10_io_out ? io_r_707_b : _GEN_8296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8298 = 10'h2c4 == r_count_10_io_out ? io_r_708_b : _GEN_8297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8299 = 10'h2c5 == r_count_10_io_out ? io_r_709_b : _GEN_8298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8300 = 10'h2c6 == r_count_10_io_out ? io_r_710_b : _GEN_8299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8301 = 10'h2c7 == r_count_10_io_out ? io_r_711_b : _GEN_8300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8302 = 10'h2c8 == r_count_10_io_out ? io_r_712_b : _GEN_8301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8303 = 10'h2c9 == r_count_10_io_out ? io_r_713_b : _GEN_8302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8304 = 10'h2ca == r_count_10_io_out ? io_r_714_b : _GEN_8303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8305 = 10'h2cb == r_count_10_io_out ? io_r_715_b : _GEN_8304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8306 = 10'h2cc == r_count_10_io_out ? io_r_716_b : _GEN_8305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8307 = 10'h2cd == r_count_10_io_out ? io_r_717_b : _GEN_8306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8308 = 10'h2ce == r_count_10_io_out ? io_r_718_b : _GEN_8307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8309 = 10'h2cf == r_count_10_io_out ? io_r_719_b : _GEN_8308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8310 = 10'h2d0 == r_count_10_io_out ? io_r_720_b : _GEN_8309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8311 = 10'h2d1 == r_count_10_io_out ? io_r_721_b : _GEN_8310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8312 = 10'h2d2 == r_count_10_io_out ? io_r_722_b : _GEN_8311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8313 = 10'h2d3 == r_count_10_io_out ? io_r_723_b : _GEN_8312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8314 = 10'h2d4 == r_count_10_io_out ? io_r_724_b : _GEN_8313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8315 = 10'h2d5 == r_count_10_io_out ? io_r_725_b : _GEN_8314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8316 = 10'h2d6 == r_count_10_io_out ? io_r_726_b : _GEN_8315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8317 = 10'h2d7 == r_count_10_io_out ? io_r_727_b : _GEN_8316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8318 = 10'h2d8 == r_count_10_io_out ? io_r_728_b : _GEN_8317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8319 = 10'h2d9 == r_count_10_io_out ? io_r_729_b : _GEN_8318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8320 = 10'h2da == r_count_10_io_out ? io_r_730_b : _GEN_8319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8321 = 10'h2db == r_count_10_io_out ? io_r_731_b : _GEN_8320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8322 = 10'h2dc == r_count_10_io_out ? io_r_732_b : _GEN_8321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8323 = 10'h2dd == r_count_10_io_out ? io_r_733_b : _GEN_8322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8324 = 10'h2de == r_count_10_io_out ? io_r_734_b : _GEN_8323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8325 = 10'h2df == r_count_10_io_out ? io_r_735_b : _GEN_8324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8326 = 10'h2e0 == r_count_10_io_out ? io_r_736_b : _GEN_8325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8327 = 10'h2e1 == r_count_10_io_out ? io_r_737_b : _GEN_8326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8328 = 10'h2e2 == r_count_10_io_out ? io_r_738_b : _GEN_8327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8329 = 10'h2e3 == r_count_10_io_out ? io_r_739_b : _GEN_8328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8330 = 10'h2e4 == r_count_10_io_out ? io_r_740_b : _GEN_8329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8331 = 10'h2e5 == r_count_10_io_out ? io_r_741_b : _GEN_8330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8332 = 10'h2e6 == r_count_10_io_out ? io_r_742_b : _GEN_8331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8333 = 10'h2e7 == r_count_10_io_out ? io_r_743_b : _GEN_8332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8334 = 10'h2e8 == r_count_10_io_out ? io_r_744_b : _GEN_8333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8335 = 10'h2e9 == r_count_10_io_out ? io_r_745_b : _GEN_8334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8336 = 10'h2ea == r_count_10_io_out ? io_r_746_b : _GEN_8335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8337 = 10'h2eb == r_count_10_io_out ? io_r_747_b : _GEN_8336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8338 = 10'h2ec == r_count_10_io_out ? io_r_748_b : _GEN_8337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8341 = 10'h1 == r_count_11_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8342 = 10'h2 == r_count_11_io_out ? io_r_2_b : _GEN_8341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8343 = 10'h3 == r_count_11_io_out ? io_r_3_b : _GEN_8342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8344 = 10'h4 == r_count_11_io_out ? io_r_4_b : _GEN_8343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8345 = 10'h5 == r_count_11_io_out ? io_r_5_b : _GEN_8344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8346 = 10'h6 == r_count_11_io_out ? io_r_6_b : _GEN_8345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8347 = 10'h7 == r_count_11_io_out ? io_r_7_b : _GEN_8346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8348 = 10'h8 == r_count_11_io_out ? io_r_8_b : _GEN_8347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8349 = 10'h9 == r_count_11_io_out ? io_r_9_b : _GEN_8348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8350 = 10'ha == r_count_11_io_out ? io_r_10_b : _GEN_8349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8351 = 10'hb == r_count_11_io_out ? io_r_11_b : _GEN_8350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8352 = 10'hc == r_count_11_io_out ? io_r_12_b : _GEN_8351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8353 = 10'hd == r_count_11_io_out ? io_r_13_b : _GEN_8352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8354 = 10'he == r_count_11_io_out ? io_r_14_b : _GEN_8353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8355 = 10'hf == r_count_11_io_out ? io_r_15_b : _GEN_8354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8356 = 10'h10 == r_count_11_io_out ? io_r_16_b : _GEN_8355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8357 = 10'h11 == r_count_11_io_out ? io_r_17_b : _GEN_8356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8358 = 10'h12 == r_count_11_io_out ? io_r_18_b : _GEN_8357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8359 = 10'h13 == r_count_11_io_out ? io_r_19_b : _GEN_8358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8360 = 10'h14 == r_count_11_io_out ? io_r_20_b : _GEN_8359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8361 = 10'h15 == r_count_11_io_out ? io_r_21_b : _GEN_8360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8362 = 10'h16 == r_count_11_io_out ? io_r_22_b : _GEN_8361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8363 = 10'h17 == r_count_11_io_out ? io_r_23_b : _GEN_8362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8364 = 10'h18 == r_count_11_io_out ? io_r_24_b : _GEN_8363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8365 = 10'h19 == r_count_11_io_out ? io_r_25_b : _GEN_8364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8366 = 10'h1a == r_count_11_io_out ? io_r_26_b : _GEN_8365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8367 = 10'h1b == r_count_11_io_out ? io_r_27_b : _GEN_8366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8368 = 10'h1c == r_count_11_io_out ? io_r_28_b : _GEN_8367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8369 = 10'h1d == r_count_11_io_out ? io_r_29_b : _GEN_8368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8370 = 10'h1e == r_count_11_io_out ? io_r_30_b : _GEN_8369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8371 = 10'h1f == r_count_11_io_out ? io_r_31_b : _GEN_8370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8372 = 10'h20 == r_count_11_io_out ? io_r_32_b : _GEN_8371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8373 = 10'h21 == r_count_11_io_out ? io_r_33_b : _GEN_8372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8374 = 10'h22 == r_count_11_io_out ? io_r_34_b : _GEN_8373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8375 = 10'h23 == r_count_11_io_out ? io_r_35_b : _GEN_8374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8376 = 10'h24 == r_count_11_io_out ? io_r_36_b : _GEN_8375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8377 = 10'h25 == r_count_11_io_out ? io_r_37_b : _GEN_8376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8378 = 10'h26 == r_count_11_io_out ? io_r_38_b : _GEN_8377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8379 = 10'h27 == r_count_11_io_out ? io_r_39_b : _GEN_8378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8380 = 10'h28 == r_count_11_io_out ? io_r_40_b : _GEN_8379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8381 = 10'h29 == r_count_11_io_out ? io_r_41_b : _GEN_8380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8382 = 10'h2a == r_count_11_io_out ? io_r_42_b : _GEN_8381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8383 = 10'h2b == r_count_11_io_out ? io_r_43_b : _GEN_8382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8384 = 10'h2c == r_count_11_io_out ? io_r_44_b : _GEN_8383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8385 = 10'h2d == r_count_11_io_out ? io_r_45_b : _GEN_8384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8386 = 10'h2e == r_count_11_io_out ? io_r_46_b : _GEN_8385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8387 = 10'h2f == r_count_11_io_out ? io_r_47_b : _GEN_8386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8388 = 10'h30 == r_count_11_io_out ? io_r_48_b : _GEN_8387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8389 = 10'h31 == r_count_11_io_out ? io_r_49_b : _GEN_8388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8390 = 10'h32 == r_count_11_io_out ? io_r_50_b : _GEN_8389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8391 = 10'h33 == r_count_11_io_out ? io_r_51_b : _GEN_8390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8392 = 10'h34 == r_count_11_io_out ? io_r_52_b : _GEN_8391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8393 = 10'h35 == r_count_11_io_out ? io_r_53_b : _GEN_8392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8394 = 10'h36 == r_count_11_io_out ? io_r_54_b : _GEN_8393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8395 = 10'h37 == r_count_11_io_out ? io_r_55_b : _GEN_8394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8396 = 10'h38 == r_count_11_io_out ? io_r_56_b : _GEN_8395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8397 = 10'h39 == r_count_11_io_out ? io_r_57_b : _GEN_8396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8398 = 10'h3a == r_count_11_io_out ? io_r_58_b : _GEN_8397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8399 = 10'h3b == r_count_11_io_out ? io_r_59_b : _GEN_8398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8400 = 10'h3c == r_count_11_io_out ? io_r_60_b : _GEN_8399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8401 = 10'h3d == r_count_11_io_out ? io_r_61_b : _GEN_8400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8402 = 10'h3e == r_count_11_io_out ? io_r_62_b : _GEN_8401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8403 = 10'h3f == r_count_11_io_out ? io_r_63_b : _GEN_8402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8404 = 10'h40 == r_count_11_io_out ? io_r_64_b : _GEN_8403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8405 = 10'h41 == r_count_11_io_out ? io_r_65_b : _GEN_8404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8406 = 10'h42 == r_count_11_io_out ? io_r_66_b : _GEN_8405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8407 = 10'h43 == r_count_11_io_out ? io_r_67_b : _GEN_8406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8408 = 10'h44 == r_count_11_io_out ? io_r_68_b : _GEN_8407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8409 = 10'h45 == r_count_11_io_out ? io_r_69_b : _GEN_8408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8410 = 10'h46 == r_count_11_io_out ? io_r_70_b : _GEN_8409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8411 = 10'h47 == r_count_11_io_out ? io_r_71_b : _GEN_8410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8412 = 10'h48 == r_count_11_io_out ? io_r_72_b : _GEN_8411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8413 = 10'h49 == r_count_11_io_out ? io_r_73_b : _GEN_8412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8414 = 10'h4a == r_count_11_io_out ? io_r_74_b : _GEN_8413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8415 = 10'h4b == r_count_11_io_out ? io_r_75_b : _GEN_8414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8416 = 10'h4c == r_count_11_io_out ? io_r_76_b : _GEN_8415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8417 = 10'h4d == r_count_11_io_out ? io_r_77_b : _GEN_8416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8418 = 10'h4e == r_count_11_io_out ? io_r_78_b : _GEN_8417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8419 = 10'h4f == r_count_11_io_out ? io_r_79_b : _GEN_8418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8420 = 10'h50 == r_count_11_io_out ? io_r_80_b : _GEN_8419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8421 = 10'h51 == r_count_11_io_out ? io_r_81_b : _GEN_8420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8422 = 10'h52 == r_count_11_io_out ? io_r_82_b : _GEN_8421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8423 = 10'h53 == r_count_11_io_out ? io_r_83_b : _GEN_8422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8424 = 10'h54 == r_count_11_io_out ? io_r_84_b : _GEN_8423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8425 = 10'h55 == r_count_11_io_out ? io_r_85_b : _GEN_8424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8426 = 10'h56 == r_count_11_io_out ? io_r_86_b : _GEN_8425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8427 = 10'h57 == r_count_11_io_out ? io_r_87_b : _GEN_8426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8428 = 10'h58 == r_count_11_io_out ? io_r_88_b : _GEN_8427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8429 = 10'h59 == r_count_11_io_out ? io_r_89_b : _GEN_8428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8430 = 10'h5a == r_count_11_io_out ? io_r_90_b : _GEN_8429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8431 = 10'h5b == r_count_11_io_out ? io_r_91_b : _GEN_8430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8432 = 10'h5c == r_count_11_io_out ? io_r_92_b : _GEN_8431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8433 = 10'h5d == r_count_11_io_out ? io_r_93_b : _GEN_8432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8434 = 10'h5e == r_count_11_io_out ? io_r_94_b : _GEN_8433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8435 = 10'h5f == r_count_11_io_out ? io_r_95_b : _GEN_8434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8436 = 10'h60 == r_count_11_io_out ? io_r_96_b : _GEN_8435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8437 = 10'h61 == r_count_11_io_out ? io_r_97_b : _GEN_8436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8438 = 10'h62 == r_count_11_io_out ? io_r_98_b : _GEN_8437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8439 = 10'h63 == r_count_11_io_out ? io_r_99_b : _GEN_8438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8440 = 10'h64 == r_count_11_io_out ? io_r_100_b : _GEN_8439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8441 = 10'h65 == r_count_11_io_out ? io_r_101_b : _GEN_8440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8442 = 10'h66 == r_count_11_io_out ? io_r_102_b : _GEN_8441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8443 = 10'h67 == r_count_11_io_out ? io_r_103_b : _GEN_8442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8444 = 10'h68 == r_count_11_io_out ? io_r_104_b : _GEN_8443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8445 = 10'h69 == r_count_11_io_out ? io_r_105_b : _GEN_8444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8446 = 10'h6a == r_count_11_io_out ? io_r_106_b : _GEN_8445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8447 = 10'h6b == r_count_11_io_out ? io_r_107_b : _GEN_8446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8448 = 10'h6c == r_count_11_io_out ? io_r_108_b : _GEN_8447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8449 = 10'h6d == r_count_11_io_out ? io_r_109_b : _GEN_8448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8450 = 10'h6e == r_count_11_io_out ? io_r_110_b : _GEN_8449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8451 = 10'h6f == r_count_11_io_out ? io_r_111_b : _GEN_8450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8452 = 10'h70 == r_count_11_io_out ? io_r_112_b : _GEN_8451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8453 = 10'h71 == r_count_11_io_out ? io_r_113_b : _GEN_8452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8454 = 10'h72 == r_count_11_io_out ? io_r_114_b : _GEN_8453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8455 = 10'h73 == r_count_11_io_out ? io_r_115_b : _GEN_8454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8456 = 10'h74 == r_count_11_io_out ? io_r_116_b : _GEN_8455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8457 = 10'h75 == r_count_11_io_out ? io_r_117_b : _GEN_8456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8458 = 10'h76 == r_count_11_io_out ? io_r_118_b : _GEN_8457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8459 = 10'h77 == r_count_11_io_out ? io_r_119_b : _GEN_8458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8460 = 10'h78 == r_count_11_io_out ? io_r_120_b : _GEN_8459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8461 = 10'h79 == r_count_11_io_out ? io_r_121_b : _GEN_8460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8462 = 10'h7a == r_count_11_io_out ? io_r_122_b : _GEN_8461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8463 = 10'h7b == r_count_11_io_out ? io_r_123_b : _GEN_8462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8464 = 10'h7c == r_count_11_io_out ? io_r_124_b : _GEN_8463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8465 = 10'h7d == r_count_11_io_out ? io_r_125_b : _GEN_8464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8466 = 10'h7e == r_count_11_io_out ? io_r_126_b : _GEN_8465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8467 = 10'h7f == r_count_11_io_out ? io_r_127_b : _GEN_8466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8468 = 10'h80 == r_count_11_io_out ? io_r_128_b : _GEN_8467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8469 = 10'h81 == r_count_11_io_out ? io_r_129_b : _GEN_8468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8470 = 10'h82 == r_count_11_io_out ? io_r_130_b : _GEN_8469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8471 = 10'h83 == r_count_11_io_out ? io_r_131_b : _GEN_8470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8472 = 10'h84 == r_count_11_io_out ? io_r_132_b : _GEN_8471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8473 = 10'h85 == r_count_11_io_out ? io_r_133_b : _GEN_8472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8474 = 10'h86 == r_count_11_io_out ? io_r_134_b : _GEN_8473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8475 = 10'h87 == r_count_11_io_out ? io_r_135_b : _GEN_8474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8476 = 10'h88 == r_count_11_io_out ? io_r_136_b : _GEN_8475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8477 = 10'h89 == r_count_11_io_out ? io_r_137_b : _GEN_8476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8478 = 10'h8a == r_count_11_io_out ? io_r_138_b : _GEN_8477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8479 = 10'h8b == r_count_11_io_out ? io_r_139_b : _GEN_8478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8480 = 10'h8c == r_count_11_io_out ? io_r_140_b : _GEN_8479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8481 = 10'h8d == r_count_11_io_out ? io_r_141_b : _GEN_8480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8482 = 10'h8e == r_count_11_io_out ? io_r_142_b : _GEN_8481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8483 = 10'h8f == r_count_11_io_out ? io_r_143_b : _GEN_8482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8484 = 10'h90 == r_count_11_io_out ? io_r_144_b : _GEN_8483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8485 = 10'h91 == r_count_11_io_out ? io_r_145_b : _GEN_8484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8486 = 10'h92 == r_count_11_io_out ? io_r_146_b : _GEN_8485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8487 = 10'h93 == r_count_11_io_out ? io_r_147_b : _GEN_8486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8488 = 10'h94 == r_count_11_io_out ? io_r_148_b : _GEN_8487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8489 = 10'h95 == r_count_11_io_out ? io_r_149_b : _GEN_8488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8490 = 10'h96 == r_count_11_io_out ? io_r_150_b : _GEN_8489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8491 = 10'h97 == r_count_11_io_out ? io_r_151_b : _GEN_8490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8492 = 10'h98 == r_count_11_io_out ? io_r_152_b : _GEN_8491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8493 = 10'h99 == r_count_11_io_out ? io_r_153_b : _GEN_8492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8494 = 10'h9a == r_count_11_io_out ? io_r_154_b : _GEN_8493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8495 = 10'h9b == r_count_11_io_out ? io_r_155_b : _GEN_8494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8496 = 10'h9c == r_count_11_io_out ? io_r_156_b : _GEN_8495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8497 = 10'h9d == r_count_11_io_out ? io_r_157_b : _GEN_8496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8498 = 10'h9e == r_count_11_io_out ? io_r_158_b : _GEN_8497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8499 = 10'h9f == r_count_11_io_out ? io_r_159_b : _GEN_8498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8500 = 10'ha0 == r_count_11_io_out ? io_r_160_b : _GEN_8499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8501 = 10'ha1 == r_count_11_io_out ? io_r_161_b : _GEN_8500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8502 = 10'ha2 == r_count_11_io_out ? io_r_162_b : _GEN_8501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8503 = 10'ha3 == r_count_11_io_out ? io_r_163_b : _GEN_8502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8504 = 10'ha4 == r_count_11_io_out ? io_r_164_b : _GEN_8503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8505 = 10'ha5 == r_count_11_io_out ? io_r_165_b : _GEN_8504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8506 = 10'ha6 == r_count_11_io_out ? io_r_166_b : _GEN_8505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8507 = 10'ha7 == r_count_11_io_out ? io_r_167_b : _GEN_8506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8508 = 10'ha8 == r_count_11_io_out ? io_r_168_b : _GEN_8507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8509 = 10'ha9 == r_count_11_io_out ? io_r_169_b : _GEN_8508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8510 = 10'haa == r_count_11_io_out ? io_r_170_b : _GEN_8509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8511 = 10'hab == r_count_11_io_out ? io_r_171_b : _GEN_8510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8512 = 10'hac == r_count_11_io_out ? io_r_172_b : _GEN_8511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8513 = 10'had == r_count_11_io_out ? io_r_173_b : _GEN_8512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8514 = 10'hae == r_count_11_io_out ? io_r_174_b : _GEN_8513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8515 = 10'haf == r_count_11_io_out ? io_r_175_b : _GEN_8514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8516 = 10'hb0 == r_count_11_io_out ? io_r_176_b : _GEN_8515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8517 = 10'hb1 == r_count_11_io_out ? io_r_177_b : _GEN_8516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8518 = 10'hb2 == r_count_11_io_out ? io_r_178_b : _GEN_8517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8519 = 10'hb3 == r_count_11_io_out ? io_r_179_b : _GEN_8518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8520 = 10'hb4 == r_count_11_io_out ? io_r_180_b : _GEN_8519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8521 = 10'hb5 == r_count_11_io_out ? io_r_181_b : _GEN_8520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8522 = 10'hb6 == r_count_11_io_out ? io_r_182_b : _GEN_8521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8523 = 10'hb7 == r_count_11_io_out ? io_r_183_b : _GEN_8522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8524 = 10'hb8 == r_count_11_io_out ? io_r_184_b : _GEN_8523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8525 = 10'hb9 == r_count_11_io_out ? io_r_185_b : _GEN_8524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8526 = 10'hba == r_count_11_io_out ? io_r_186_b : _GEN_8525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8527 = 10'hbb == r_count_11_io_out ? io_r_187_b : _GEN_8526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8528 = 10'hbc == r_count_11_io_out ? io_r_188_b : _GEN_8527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8529 = 10'hbd == r_count_11_io_out ? io_r_189_b : _GEN_8528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8530 = 10'hbe == r_count_11_io_out ? io_r_190_b : _GEN_8529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8531 = 10'hbf == r_count_11_io_out ? io_r_191_b : _GEN_8530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8532 = 10'hc0 == r_count_11_io_out ? io_r_192_b : _GEN_8531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8533 = 10'hc1 == r_count_11_io_out ? io_r_193_b : _GEN_8532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8534 = 10'hc2 == r_count_11_io_out ? io_r_194_b : _GEN_8533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8535 = 10'hc3 == r_count_11_io_out ? io_r_195_b : _GEN_8534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8536 = 10'hc4 == r_count_11_io_out ? io_r_196_b : _GEN_8535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8537 = 10'hc5 == r_count_11_io_out ? io_r_197_b : _GEN_8536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8538 = 10'hc6 == r_count_11_io_out ? io_r_198_b : _GEN_8537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8539 = 10'hc7 == r_count_11_io_out ? io_r_199_b : _GEN_8538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8540 = 10'hc8 == r_count_11_io_out ? io_r_200_b : _GEN_8539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8541 = 10'hc9 == r_count_11_io_out ? io_r_201_b : _GEN_8540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8542 = 10'hca == r_count_11_io_out ? io_r_202_b : _GEN_8541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8543 = 10'hcb == r_count_11_io_out ? io_r_203_b : _GEN_8542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8544 = 10'hcc == r_count_11_io_out ? io_r_204_b : _GEN_8543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8545 = 10'hcd == r_count_11_io_out ? io_r_205_b : _GEN_8544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8546 = 10'hce == r_count_11_io_out ? io_r_206_b : _GEN_8545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8547 = 10'hcf == r_count_11_io_out ? io_r_207_b : _GEN_8546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8548 = 10'hd0 == r_count_11_io_out ? io_r_208_b : _GEN_8547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8549 = 10'hd1 == r_count_11_io_out ? io_r_209_b : _GEN_8548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8550 = 10'hd2 == r_count_11_io_out ? io_r_210_b : _GEN_8549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8551 = 10'hd3 == r_count_11_io_out ? io_r_211_b : _GEN_8550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8552 = 10'hd4 == r_count_11_io_out ? io_r_212_b : _GEN_8551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8553 = 10'hd5 == r_count_11_io_out ? io_r_213_b : _GEN_8552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8554 = 10'hd6 == r_count_11_io_out ? io_r_214_b : _GEN_8553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8555 = 10'hd7 == r_count_11_io_out ? io_r_215_b : _GEN_8554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8556 = 10'hd8 == r_count_11_io_out ? io_r_216_b : _GEN_8555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8557 = 10'hd9 == r_count_11_io_out ? io_r_217_b : _GEN_8556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8558 = 10'hda == r_count_11_io_out ? io_r_218_b : _GEN_8557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8559 = 10'hdb == r_count_11_io_out ? io_r_219_b : _GEN_8558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8560 = 10'hdc == r_count_11_io_out ? io_r_220_b : _GEN_8559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8561 = 10'hdd == r_count_11_io_out ? io_r_221_b : _GEN_8560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8562 = 10'hde == r_count_11_io_out ? io_r_222_b : _GEN_8561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8563 = 10'hdf == r_count_11_io_out ? io_r_223_b : _GEN_8562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8564 = 10'he0 == r_count_11_io_out ? io_r_224_b : _GEN_8563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8565 = 10'he1 == r_count_11_io_out ? io_r_225_b : _GEN_8564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8566 = 10'he2 == r_count_11_io_out ? io_r_226_b : _GEN_8565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8567 = 10'he3 == r_count_11_io_out ? io_r_227_b : _GEN_8566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8568 = 10'he4 == r_count_11_io_out ? io_r_228_b : _GEN_8567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8569 = 10'he5 == r_count_11_io_out ? io_r_229_b : _GEN_8568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8570 = 10'he6 == r_count_11_io_out ? io_r_230_b : _GEN_8569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8571 = 10'he7 == r_count_11_io_out ? io_r_231_b : _GEN_8570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8572 = 10'he8 == r_count_11_io_out ? io_r_232_b : _GEN_8571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8573 = 10'he9 == r_count_11_io_out ? io_r_233_b : _GEN_8572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8574 = 10'hea == r_count_11_io_out ? io_r_234_b : _GEN_8573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8575 = 10'heb == r_count_11_io_out ? io_r_235_b : _GEN_8574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8576 = 10'hec == r_count_11_io_out ? io_r_236_b : _GEN_8575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8577 = 10'hed == r_count_11_io_out ? io_r_237_b : _GEN_8576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8578 = 10'hee == r_count_11_io_out ? io_r_238_b : _GEN_8577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8579 = 10'hef == r_count_11_io_out ? io_r_239_b : _GEN_8578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8580 = 10'hf0 == r_count_11_io_out ? io_r_240_b : _GEN_8579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8581 = 10'hf1 == r_count_11_io_out ? io_r_241_b : _GEN_8580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8582 = 10'hf2 == r_count_11_io_out ? io_r_242_b : _GEN_8581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8583 = 10'hf3 == r_count_11_io_out ? io_r_243_b : _GEN_8582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8584 = 10'hf4 == r_count_11_io_out ? io_r_244_b : _GEN_8583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8585 = 10'hf5 == r_count_11_io_out ? io_r_245_b : _GEN_8584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8586 = 10'hf6 == r_count_11_io_out ? io_r_246_b : _GEN_8585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8587 = 10'hf7 == r_count_11_io_out ? io_r_247_b : _GEN_8586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8588 = 10'hf8 == r_count_11_io_out ? io_r_248_b : _GEN_8587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8589 = 10'hf9 == r_count_11_io_out ? io_r_249_b : _GEN_8588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8590 = 10'hfa == r_count_11_io_out ? io_r_250_b : _GEN_8589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8591 = 10'hfb == r_count_11_io_out ? io_r_251_b : _GEN_8590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8592 = 10'hfc == r_count_11_io_out ? io_r_252_b : _GEN_8591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8593 = 10'hfd == r_count_11_io_out ? io_r_253_b : _GEN_8592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8594 = 10'hfe == r_count_11_io_out ? io_r_254_b : _GEN_8593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8595 = 10'hff == r_count_11_io_out ? io_r_255_b : _GEN_8594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8596 = 10'h100 == r_count_11_io_out ? io_r_256_b : _GEN_8595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8597 = 10'h101 == r_count_11_io_out ? io_r_257_b : _GEN_8596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8598 = 10'h102 == r_count_11_io_out ? io_r_258_b : _GEN_8597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8599 = 10'h103 == r_count_11_io_out ? io_r_259_b : _GEN_8598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8600 = 10'h104 == r_count_11_io_out ? io_r_260_b : _GEN_8599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8601 = 10'h105 == r_count_11_io_out ? io_r_261_b : _GEN_8600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8602 = 10'h106 == r_count_11_io_out ? io_r_262_b : _GEN_8601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8603 = 10'h107 == r_count_11_io_out ? io_r_263_b : _GEN_8602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8604 = 10'h108 == r_count_11_io_out ? io_r_264_b : _GEN_8603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8605 = 10'h109 == r_count_11_io_out ? io_r_265_b : _GEN_8604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8606 = 10'h10a == r_count_11_io_out ? io_r_266_b : _GEN_8605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8607 = 10'h10b == r_count_11_io_out ? io_r_267_b : _GEN_8606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8608 = 10'h10c == r_count_11_io_out ? io_r_268_b : _GEN_8607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8609 = 10'h10d == r_count_11_io_out ? io_r_269_b : _GEN_8608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8610 = 10'h10e == r_count_11_io_out ? io_r_270_b : _GEN_8609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8611 = 10'h10f == r_count_11_io_out ? io_r_271_b : _GEN_8610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8612 = 10'h110 == r_count_11_io_out ? io_r_272_b : _GEN_8611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8613 = 10'h111 == r_count_11_io_out ? io_r_273_b : _GEN_8612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8614 = 10'h112 == r_count_11_io_out ? io_r_274_b : _GEN_8613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8615 = 10'h113 == r_count_11_io_out ? io_r_275_b : _GEN_8614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8616 = 10'h114 == r_count_11_io_out ? io_r_276_b : _GEN_8615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8617 = 10'h115 == r_count_11_io_out ? io_r_277_b : _GEN_8616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8618 = 10'h116 == r_count_11_io_out ? io_r_278_b : _GEN_8617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8619 = 10'h117 == r_count_11_io_out ? io_r_279_b : _GEN_8618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8620 = 10'h118 == r_count_11_io_out ? io_r_280_b : _GEN_8619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8621 = 10'h119 == r_count_11_io_out ? io_r_281_b : _GEN_8620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8622 = 10'h11a == r_count_11_io_out ? io_r_282_b : _GEN_8621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8623 = 10'h11b == r_count_11_io_out ? io_r_283_b : _GEN_8622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8624 = 10'h11c == r_count_11_io_out ? io_r_284_b : _GEN_8623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8625 = 10'h11d == r_count_11_io_out ? io_r_285_b : _GEN_8624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8626 = 10'h11e == r_count_11_io_out ? io_r_286_b : _GEN_8625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8627 = 10'h11f == r_count_11_io_out ? io_r_287_b : _GEN_8626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8628 = 10'h120 == r_count_11_io_out ? io_r_288_b : _GEN_8627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8629 = 10'h121 == r_count_11_io_out ? io_r_289_b : _GEN_8628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8630 = 10'h122 == r_count_11_io_out ? io_r_290_b : _GEN_8629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8631 = 10'h123 == r_count_11_io_out ? io_r_291_b : _GEN_8630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8632 = 10'h124 == r_count_11_io_out ? io_r_292_b : _GEN_8631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8633 = 10'h125 == r_count_11_io_out ? io_r_293_b : _GEN_8632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8634 = 10'h126 == r_count_11_io_out ? io_r_294_b : _GEN_8633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8635 = 10'h127 == r_count_11_io_out ? io_r_295_b : _GEN_8634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8636 = 10'h128 == r_count_11_io_out ? io_r_296_b : _GEN_8635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8637 = 10'h129 == r_count_11_io_out ? io_r_297_b : _GEN_8636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8638 = 10'h12a == r_count_11_io_out ? io_r_298_b : _GEN_8637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8639 = 10'h12b == r_count_11_io_out ? io_r_299_b : _GEN_8638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8640 = 10'h12c == r_count_11_io_out ? io_r_300_b : _GEN_8639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8641 = 10'h12d == r_count_11_io_out ? io_r_301_b : _GEN_8640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8642 = 10'h12e == r_count_11_io_out ? io_r_302_b : _GEN_8641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8643 = 10'h12f == r_count_11_io_out ? io_r_303_b : _GEN_8642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8644 = 10'h130 == r_count_11_io_out ? io_r_304_b : _GEN_8643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8645 = 10'h131 == r_count_11_io_out ? io_r_305_b : _GEN_8644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8646 = 10'h132 == r_count_11_io_out ? io_r_306_b : _GEN_8645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8647 = 10'h133 == r_count_11_io_out ? io_r_307_b : _GEN_8646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8648 = 10'h134 == r_count_11_io_out ? io_r_308_b : _GEN_8647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8649 = 10'h135 == r_count_11_io_out ? io_r_309_b : _GEN_8648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8650 = 10'h136 == r_count_11_io_out ? io_r_310_b : _GEN_8649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8651 = 10'h137 == r_count_11_io_out ? io_r_311_b : _GEN_8650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8652 = 10'h138 == r_count_11_io_out ? io_r_312_b : _GEN_8651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8653 = 10'h139 == r_count_11_io_out ? io_r_313_b : _GEN_8652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8654 = 10'h13a == r_count_11_io_out ? io_r_314_b : _GEN_8653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8655 = 10'h13b == r_count_11_io_out ? io_r_315_b : _GEN_8654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8656 = 10'h13c == r_count_11_io_out ? io_r_316_b : _GEN_8655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8657 = 10'h13d == r_count_11_io_out ? io_r_317_b : _GEN_8656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8658 = 10'h13e == r_count_11_io_out ? io_r_318_b : _GEN_8657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8659 = 10'h13f == r_count_11_io_out ? io_r_319_b : _GEN_8658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8660 = 10'h140 == r_count_11_io_out ? io_r_320_b : _GEN_8659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8661 = 10'h141 == r_count_11_io_out ? io_r_321_b : _GEN_8660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8662 = 10'h142 == r_count_11_io_out ? io_r_322_b : _GEN_8661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8663 = 10'h143 == r_count_11_io_out ? io_r_323_b : _GEN_8662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8664 = 10'h144 == r_count_11_io_out ? io_r_324_b : _GEN_8663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8665 = 10'h145 == r_count_11_io_out ? io_r_325_b : _GEN_8664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8666 = 10'h146 == r_count_11_io_out ? io_r_326_b : _GEN_8665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8667 = 10'h147 == r_count_11_io_out ? io_r_327_b : _GEN_8666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8668 = 10'h148 == r_count_11_io_out ? io_r_328_b : _GEN_8667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8669 = 10'h149 == r_count_11_io_out ? io_r_329_b : _GEN_8668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8670 = 10'h14a == r_count_11_io_out ? io_r_330_b : _GEN_8669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8671 = 10'h14b == r_count_11_io_out ? io_r_331_b : _GEN_8670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8672 = 10'h14c == r_count_11_io_out ? io_r_332_b : _GEN_8671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8673 = 10'h14d == r_count_11_io_out ? io_r_333_b : _GEN_8672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8674 = 10'h14e == r_count_11_io_out ? io_r_334_b : _GEN_8673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8675 = 10'h14f == r_count_11_io_out ? io_r_335_b : _GEN_8674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8676 = 10'h150 == r_count_11_io_out ? io_r_336_b : _GEN_8675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8677 = 10'h151 == r_count_11_io_out ? io_r_337_b : _GEN_8676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8678 = 10'h152 == r_count_11_io_out ? io_r_338_b : _GEN_8677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8679 = 10'h153 == r_count_11_io_out ? io_r_339_b : _GEN_8678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8680 = 10'h154 == r_count_11_io_out ? io_r_340_b : _GEN_8679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8681 = 10'h155 == r_count_11_io_out ? io_r_341_b : _GEN_8680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8682 = 10'h156 == r_count_11_io_out ? io_r_342_b : _GEN_8681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8683 = 10'h157 == r_count_11_io_out ? io_r_343_b : _GEN_8682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8684 = 10'h158 == r_count_11_io_out ? io_r_344_b : _GEN_8683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8685 = 10'h159 == r_count_11_io_out ? io_r_345_b : _GEN_8684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8686 = 10'h15a == r_count_11_io_out ? io_r_346_b : _GEN_8685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8687 = 10'h15b == r_count_11_io_out ? io_r_347_b : _GEN_8686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8688 = 10'h15c == r_count_11_io_out ? io_r_348_b : _GEN_8687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8689 = 10'h15d == r_count_11_io_out ? io_r_349_b : _GEN_8688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8690 = 10'h15e == r_count_11_io_out ? io_r_350_b : _GEN_8689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8691 = 10'h15f == r_count_11_io_out ? io_r_351_b : _GEN_8690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8692 = 10'h160 == r_count_11_io_out ? io_r_352_b : _GEN_8691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8693 = 10'h161 == r_count_11_io_out ? io_r_353_b : _GEN_8692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8694 = 10'h162 == r_count_11_io_out ? io_r_354_b : _GEN_8693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8695 = 10'h163 == r_count_11_io_out ? io_r_355_b : _GEN_8694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8696 = 10'h164 == r_count_11_io_out ? io_r_356_b : _GEN_8695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8697 = 10'h165 == r_count_11_io_out ? io_r_357_b : _GEN_8696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8698 = 10'h166 == r_count_11_io_out ? io_r_358_b : _GEN_8697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8699 = 10'h167 == r_count_11_io_out ? io_r_359_b : _GEN_8698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8700 = 10'h168 == r_count_11_io_out ? io_r_360_b : _GEN_8699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8701 = 10'h169 == r_count_11_io_out ? io_r_361_b : _GEN_8700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8702 = 10'h16a == r_count_11_io_out ? io_r_362_b : _GEN_8701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8703 = 10'h16b == r_count_11_io_out ? io_r_363_b : _GEN_8702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8704 = 10'h16c == r_count_11_io_out ? io_r_364_b : _GEN_8703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8705 = 10'h16d == r_count_11_io_out ? io_r_365_b : _GEN_8704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8706 = 10'h16e == r_count_11_io_out ? io_r_366_b : _GEN_8705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8707 = 10'h16f == r_count_11_io_out ? io_r_367_b : _GEN_8706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8708 = 10'h170 == r_count_11_io_out ? io_r_368_b : _GEN_8707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8709 = 10'h171 == r_count_11_io_out ? io_r_369_b : _GEN_8708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8710 = 10'h172 == r_count_11_io_out ? io_r_370_b : _GEN_8709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8711 = 10'h173 == r_count_11_io_out ? io_r_371_b : _GEN_8710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8712 = 10'h174 == r_count_11_io_out ? io_r_372_b : _GEN_8711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8713 = 10'h175 == r_count_11_io_out ? io_r_373_b : _GEN_8712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8714 = 10'h176 == r_count_11_io_out ? io_r_374_b : _GEN_8713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8715 = 10'h177 == r_count_11_io_out ? io_r_375_b : _GEN_8714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8716 = 10'h178 == r_count_11_io_out ? io_r_376_b : _GEN_8715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8717 = 10'h179 == r_count_11_io_out ? io_r_377_b : _GEN_8716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8718 = 10'h17a == r_count_11_io_out ? io_r_378_b : _GEN_8717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8719 = 10'h17b == r_count_11_io_out ? io_r_379_b : _GEN_8718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8720 = 10'h17c == r_count_11_io_out ? io_r_380_b : _GEN_8719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8721 = 10'h17d == r_count_11_io_out ? io_r_381_b : _GEN_8720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8722 = 10'h17e == r_count_11_io_out ? io_r_382_b : _GEN_8721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8723 = 10'h17f == r_count_11_io_out ? io_r_383_b : _GEN_8722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8724 = 10'h180 == r_count_11_io_out ? io_r_384_b : _GEN_8723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8725 = 10'h181 == r_count_11_io_out ? io_r_385_b : _GEN_8724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8726 = 10'h182 == r_count_11_io_out ? io_r_386_b : _GEN_8725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8727 = 10'h183 == r_count_11_io_out ? io_r_387_b : _GEN_8726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8728 = 10'h184 == r_count_11_io_out ? io_r_388_b : _GEN_8727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8729 = 10'h185 == r_count_11_io_out ? io_r_389_b : _GEN_8728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8730 = 10'h186 == r_count_11_io_out ? io_r_390_b : _GEN_8729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8731 = 10'h187 == r_count_11_io_out ? io_r_391_b : _GEN_8730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8732 = 10'h188 == r_count_11_io_out ? io_r_392_b : _GEN_8731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8733 = 10'h189 == r_count_11_io_out ? io_r_393_b : _GEN_8732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8734 = 10'h18a == r_count_11_io_out ? io_r_394_b : _GEN_8733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8735 = 10'h18b == r_count_11_io_out ? io_r_395_b : _GEN_8734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8736 = 10'h18c == r_count_11_io_out ? io_r_396_b : _GEN_8735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8737 = 10'h18d == r_count_11_io_out ? io_r_397_b : _GEN_8736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8738 = 10'h18e == r_count_11_io_out ? io_r_398_b : _GEN_8737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8739 = 10'h18f == r_count_11_io_out ? io_r_399_b : _GEN_8738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8740 = 10'h190 == r_count_11_io_out ? io_r_400_b : _GEN_8739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8741 = 10'h191 == r_count_11_io_out ? io_r_401_b : _GEN_8740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8742 = 10'h192 == r_count_11_io_out ? io_r_402_b : _GEN_8741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8743 = 10'h193 == r_count_11_io_out ? io_r_403_b : _GEN_8742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8744 = 10'h194 == r_count_11_io_out ? io_r_404_b : _GEN_8743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8745 = 10'h195 == r_count_11_io_out ? io_r_405_b : _GEN_8744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8746 = 10'h196 == r_count_11_io_out ? io_r_406_b : _GEN_8745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8747 = 10'h197 == r_count_11_io_out ? io_r_407_b : _GEN_8746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8748 = 10'h198 == r_count_11_io_out ? io_r_408_b : _GEN_8747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8749 = 10'h199 == r_count_11_io_out ? io_r_409_b : _GEN_8748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8750 = 10'h19a == r_count_11_io_out ? io_r_410_b : _GEN_8749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8751 = 10'h19b == r_count_11_io_out ? io_r_411_b : _GEN_8750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8752 = 10'h19c == r_count_11_io_out ? io_r_412_b : _GEN_8751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8753 = 10'h19d == r_count_11_io_out ? io_r_413_b : _GEN_8752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8754 = 10'h19e == r_count_11_io_out ? io_r_414_b : _GEN_8753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8755 = 10'h19f == r_count_11_io_out ? io_r_415_b : _GEN_8754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8756 = 10'h1a0 == r_count_11_io_out ? io_r_416_b : _GEN_8755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8757 = 10'h1a1 == r_count_11_io_out ? io_r_417_b : _GEN_8756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8758 = 10'h1a2 == r_count_11_io_out ? io_r_418_b : _GEN_8757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8759 = 10'h1a3 == r_count_11_io_out ? io_r_419_b : _GEN_8758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8760 = 10'h1a4 == r_count_11_io_out ? io_r_420_b : _GEN_8759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8761 = 10'h1a5 == r_count_11_io_out ? io_r_421_b : _GEN_8760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8762 = 10'h1a6 == r_count_11_io_out ? io_r_422_b : _GEN_8761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8763 = 10'h1a7 == r_count_11_io_out ? io_r_423_b : _GEN_8762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8764 = 10'h1a8 == r_count_11_io_out ? io_r_424_b : _GEN_8763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8765 = 10'h1a9 == r_count_11_io_out ? io_r_425_b : _GEN_8764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8766 = 10'h1aa == r_count_11_io_out ? io_r_426_b : _GEN_8765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8767 = 10'h1ab == r_count_11_io_out ? io_r_427_b : _GEN_8766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8768 = 10'h1ac == r_count_11_io_out ? io_r_428_b : _GEN_8767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8769 = 10'h1ad == r_count_11_io_out ? io_r_429_b : _GEN_8768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8770 = 10'h1ae == r_count_11_io_out ? io_r_430_b : _GEN_8769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8771 = 10'h1af == r_count_11_io_out ? io_r_431_b : _GEN_8770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8772 = 10'h1b0 == r_count_11_io_out ? io_r_432_b : _GEN_8771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8773 = 10'h1b1 == r_count_11_io_out ? io_r_433_b : _GEN_8772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8774 = 10'h1b2 == r_count_11_io_out ? io_r_434_b : _GEN_8773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8775 = 10'h1b3 == r_count_11_io_out ? io_r_435_b : _GEN_8774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8776 = 10'h1b4 == r_count_11_io_out ? io_r_436_b : _GEN_8775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8777 = 10'h1b5 == r_count_11_io_out ? io_r_437_b : _GEN_8776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8778 = 10'h1b6 == r_count_11_io_out ? io_r_438_b : _GEN_8777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8779 = 10'h1b7 == r_count_11_io_out ? io_r_439_b : _GEN_8778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8780 = 10'h1b8 == r_count_11_io_out ? io_r_440_b : _GEN_8779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8781 = 10'h1b9 == r_count_11_io_out ? io_r_441_b : _GEN_8780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8782 = 10'h1ba == r_count_11_io_out ? io_r_442_b : _GEN_8781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8783 = 10'h1bb == r_count_11_io_out ? io_r_443_b : _GEN_8782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8784 = 10'h1bc == r_count_11_io_out ? io_r_444_b : _GEN_8783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8785 = 10'h1bd == r_count_11_io_out ? io_r_445_b : _GEN_8784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8786 = 10'h1be == r_count_11_io_out ? io_r_446_b : _GEN_8785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8787 = 10'h1bf == r_count_11_io_out ? io_r_447_b : _GEN_8786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8788 = 10'h1c0 == r_count_11_io_out ? io_r_448_b : _GEN_8787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8789 = 10'h1c1 == r_count_11_io_out ? io_r_449_b : _GEN_8788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8790 = 10'h1c2 == r_count_11_io_out ? io_r_450_b : _GEN_8789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8791 = 10'h1c3 == r_count_11_io_out ? io_r_451_b : _GEN_8790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8792 = 10'h1c4 == r_count_11_io_out ? io_r_452_b : _GEN_8791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8793 = 10'h1c5 == r_count_11_io_out ? io_r_453_b : _GEN_8792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8794 = 10'h1c6 == r_count_11_io_out ? io_r_454_b : _GEN_8793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8795 = 10'h1c7 == r_count_11_io_out ? io_r_455_b : _GEN_8794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8796 = 10'h1c8 == r_count_11_io_out ? io_r_456_b : _GEN_8795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8797 = 10'h1c9 == r_count_11_io_out ? io_r_457_b : _GEN_8796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8798 = 10'h1ca == r_count_11_io_out ? io_r_458_b : _GEN_8797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8799 = 10'h1cb == r_count_11_io_out ? io_r_459_b : _GEN_8798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8800 = 10'h1cc == r_count_11_io_out ? io_r_460_b : _GEN_8799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8801 = 10'h1cd == r_count_11_io_out ? io_r_461_b : _GEN_8800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8802 = 10'h1ce == r_count_11_io_out ? io_r_462_b : _GEN_8801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8803 = 10'h1cf == r_count_11_io_out ? io_r_463_b : _GEN_8802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8804 = 10'h1d0 == r_count_11_io_out ? io_r_464_b : _GEN_8803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8805 = 10'h1d1 == r_count_11_io_out ? io_r_465_b : _GEN_8804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8806 = 10'h1d2 == r_count_11_io_out ? io_r_466_b : _GEN_8805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8807 = 10'h1d3 == r_count_11_io_out ? io_r_467_b : _GEN_8806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8808 = 10'h1d4 == r_count_11_io_out ? io_r_468_b : _GEN_8807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8809 = 10'h1d5 == r_count_11_io_out ? io_r_469_b : _GEN_8808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8810 = 10'h1d6 == r_count_11_io_out ? io_r_470_b : _GEN_8809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8811 = 10'h1d7 == r_count_11_io_out ? io_r_471_b : _GEN_8810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8812 = 10'h1d8 == r_count_11_io_out ? io_r_472_b : _GEN_8811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8813 = 10'h1d9 == r_count_11_io_out ? io_r_473_b : _GEN_8812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8814 = 10'h1da == r_count_11_io_out ? io_r_474_b : _GEN_8813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8815 = 10'h1db == r_count_11_io_out ? io_r_475_b : _GEN_8814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8816 = 10'h1dc == r_count_11_io_out ? io_r_476_b : _GEN_8815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8817 = 10'h1dd == r_count_11_io_out ? io_r_477_b : _GEN_8816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8818 = 10'h1de == r_count_11_io_out ? io_r_478_b : _GEN_8817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8819 = 10'h1df == r_count_11_io_out ? io_r_479_b : _GEN_8818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8820 = 10'h1e0 == r_count_11_io_out ? io_r_480_b : _GEN_8819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8821 = 10'h1e1 == r_count_11_io_out ? io_r_481_b : _GEN_8820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8822 = 10'h1e2 == r_count_11_io_out ? io_r_482_b : _GEN_8821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8823 = 10'h1e3 == r_count_11_io_out ? io_r_483_b : _GEN_8822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8824 = 10'h1e4 == r_count_11_io_out ? io_r_484_b : _GEN_8823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8825 = 10'h1e5 == r_count_11_io_out ? io_r_485_b : _GEN_8824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8826 = 10'h1e6 == r_count_11_io_out ? io_r_486_b : _GEN_8825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8827 = 10'h1e7 == r_count_11_io_out ? io_r_487_b : _GEN_8826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8828 = 10'h1e8 == r_count_11_io_out ? io_r_488_b : _GEN_8827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8829 = 10'h1e9 == r_count_11_io_out ? io_r_489_b : _GEN_8828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8830 = 10'h1ea == r_count_11_io_out ? io_r_490_b : _GEN_8829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8831 = 10'h1eb == r_count_11_io_out ? io_r_491_b : _GEN_8830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8832 = 10'h1ec == r_count_11_io_out ? io_r_492_b : _GEN_8831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8833 = 10'h1ed == r_count_11_io_out ? io_r_493_b : _GEN_8832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8834 = 10'h1ee == r_count_11_io_out ? io_r_494_b : _GEN_8833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8835 = 10'h1ef == r_count_11_io_out ? io_r_495_b : _GEN_8834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8836 = 10'h1f0 == r_count_11_io_out ? io_r_496_b : _GEN_8835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8837 = 10'h1f1 == r_count_11_io_out ? io_r_497_b : _GEN_8836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8838 = 10'h1f2 == r_count_11_io_out ? io_r_498_b : _GEN_8837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8839 = 10'h1f3 == r_count_11_io_out ? io_r_499_b : _GEN_8838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8840 = 10'h1f4 == r_count_11_io_out ? io_r_500_b : _GEN_8839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8841 = 10'h1f5 == r_count_11_io_out ? io_r_501_b : _GEN_8840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8842 = 10'h1f6 == r_count_11_io_out ? io_r_502_b : _GEN_8841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8843 = 10'h1f7 == r_count_11_io_out ? io_r_503_b : _GEN_8842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8844 = 10'h1f8 == r_count_11_io_out ? io_r_504_b : _GEN_8843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8845 = 10'h1f9 == r_count_11_io_out ? io_r_505_b : _GEN_8844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8846 = 10'h1fa == r_count_11_io_out ? io_r_506_b : _GEN_8845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8847 = 10'h1fb == r_count_11_io_out ? io_r_507_b : _GEN_8846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8848 = 10'h1fc == r_count_11_io_out ? io_r_508_b : _GEN_8847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8849 = 10'h1fd == r_count_11_io_out ? io_r_509_b : _GEN_8848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8850 = 10'h1fe == r_count_11_io_out ? io_r_510_b : _GEN_8849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8851 = 10'h1ff == r_count_11_io_out ? io_r_511_b : _GEN_8850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8852 = 10'h200 == r_count_11_io_out ? io_r_512_b : _GEN_8851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8853 = 10'h201 == r_count_11_io_out ? io_r_513_b : _GEN_8852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8854 = 10'h202 == r_count_11_io_out ? io_r_514_b : _GEN_8853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8855 = 10'h203 == r_count_11_io_out ? io_r_515_b : _GEN_8854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8856 = 10'h204 == r_count_11_io_out ? io_r_516_b : _GEN_8855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8857 = 10'h205 == r_count_11_io_out ? io_r_517_b : _GEN_8856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8858 = 10'h206 == r_count_11_io_out ? io_r_518_b : _GEN_8857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8859 = 10'h207 == r_count_11_io_out ? io_r_519_b : _GEN_8858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8860 = 10'h208 == r_count_11_io_out ? io_r_520_b : _GEN_8859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8861 = 10'h209 == r_count_11_io_out ? io_r_521_b : _GEN_8860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8862 = 10'h20a == r_count_11_io_out ? io_r_522_b : _GEN_8861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8863 = 10'h20b == r_count_11_io_out ? io_r_523_b : _GEN_8862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8864 = 10'h20c == r_count_11_io_out ? io_r_524_b : _GEN_8863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8865 = 10'h20d == r_count_11_io_out ? io_r_525_b : _GEN_8864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8866 = 10'h20e == r_count_11_io_out ? io_r_526_b : _GEN_8865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8867 = 10'h20f == r_count_11_io_out ? io_r_527_b : _GEN_8866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8868 = 10'h210 == r_count_11_io_out ? io_r_528_b : _GEN_8867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8869 = 10'h211 == r_count_11_io_out ? io_r_529_b : _GEN_8868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8870 = 10'h212 == r_count_11_io_out ? io_r_530_b : _GEN_8869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8871 = 10'h213 == r_count_11_io_out ? io_r_531_b : _GEN_8870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8872 = 10'h214 == r_count_11_io_out ? io_r_532_b : _GEN_8871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8873 = 10'h215 == r_count_11_io_out ? io_r_533_b : _GEN_8872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8874 = 10'h216 == r_count_11_io_out ? io_r_534_b : _GEN_8873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8875 = 10'h217 == r_count_11_io_out ? io_r_535_b : _GEN_8874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8876 = 10'h218 == r_count_11_io_out ? io_r_536_b : _GEN_8875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8877 = 10'h219 == r_count_11_io_out ? io_r_537_b : _GEN_8876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8878 = 10'h21a == r_count_11_io_out ? io_r_538_b : _GEN_8877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8879 = 10'h21b == r_count_11_io_out ? io_r_539_b : _GEN_8878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8880 = 10'h21c == r_count_11_io_out ? io_r_540_b : _GEN_8879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8881 = 10'h21d == r_count_11_io_out ? io_r_541_b : _GEN_8880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8882 = 10'h21e == r_count_11_io_out ? io_r_542_b : _GEN_8881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8883 = 10'h21f == r_count_11_io_out ? io_r_543_b : _GEN_8882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8884 = 10'h220 == r_count_11_io_out ? io_r_544_b : _GEN_8883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8885 = 10'h221 == r_count_11_io_out ? io_r_545_b : _GEN_8884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8886 = 10'h222 == r_count_11_io_out ? io_r_546_b : _GEN_8885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8887 = 10'h223 == r_count_11_io_out ? io_r_547_b : _GEN_8886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8888 = 10'h224 == r_count_11_io_out ? io_r_548_b : _GEN_8887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8889 = 10'h225 == r_count_11_io_out ? io_r_549_b : _GEN_8888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8890 = 10'h226 == r_count_11_io_out ? io_r_550_b : _GEN_8889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8891 = 10'h227 == r_count_11_io_out ? io_r_551_b : _GEN_8890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8892 = 10'h228 == r_count_11_io_out ? io_r_552_b : _GEN_8891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8893 = 10'h229 == r_count_11_io_out ? io_r_553_b : _GEN_8892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8894 = 10'h22a == r_count_11_io_out ? io_r_554_b : _GEN_8893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8895 = 10'h22b == r_count_11_io_out ? io_r_555_b : _GEN_8894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8896 = 10'h22c == r_count_11_io_out ? io_r_556_b : _GEN_8895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8897 = 10'h22d == r_count_11_io_out ? io_r_557_b : _GEN_8896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8898 = 10'h22e == r_count_11_io_out ? io_r_558_b : _GEN_8897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8899 = 10'h22f == r_count_11_io_out ? io_r_559_b : _GEN_8898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8900 = 10'h230 == r_count_11_io_out ? io_r_560_b : _GEN_8899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8901 = 10'h231 == r_count_11_io_out ? io_r_561_b : _GEN_8900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8902 = 10'h232 == r_count_11_io_out ? io_r_562_b : _GEN_8901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8903 = 10'h233 == r_count_11_io_out ? io_r_563_b : _GEN_8902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8904 = 10'h234 == r_count_11_io_out ? io_r_564_b : _GEN_8903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8905 = 10'h235 == r_count_11_io_out ? io_r_565_b : _GEN_8904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8906 = 10'h236 == r_count_11_io_out ? io_r_566_b : _GEN_8905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8907 = 10'h237 == r_count_11_io_out ? io_r_567_b : _GEN_8906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8908 = 10'h238 == r_count_11_io_out ? io_r_568_b : _GEN_8907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8909 = 10'h239 == r_count_11_io_out ? io_r_569_b : _GEN_8908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8910 = 10'h23a == r_count_11_io_out ? io_r_570_b : _GEN_8909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8911 = 10'h23b == r_count_11_io_out ? io_r_571_b : _GEN_8910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8912 = 10'h23c == r_count_11_io_out ? io_r_572_b : _GEN_8911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8913 = 10'h23d == r_count_11_io_out ? io_r_573_b : _GEN_8912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8914 = 10'h23e == r_count_11_io_out ? io_r_574_b : _GEN_8913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8915 = 10'h23f == r_count_11_io_out ? io_r_575_b : _GEN_8914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8916 = 10'h240 == r_count_11_io_out ? io_r_576_b : _GEN_8915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8917 = 10'h241 == r_count_11_io_out ? io_r_577_b : _GEN_8916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8918 = 10'h242 == r_count_11_io_out ? io_r_578_b : _GEN_8917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8919 = 10'h243 == r_count_11_io_out ? io_r_579_b : _GEN_8918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8920 = 10'h244 == r_count_11_io_out ? io_r_580_b : _GEN_8919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8921 = 10'h245 == r_count_11_io_out ? io_r_581_b : _GEN_8920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8922 = 10'h246 == r_count_11_io_out ? io_r_582_b : _GEN_8921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8923 = 10'h247 == r_count_11_io_out ? io_r_583_b : _GEN_8922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8924 = 10'h248 == r_count_11_io_out ? io_r_584_b : _GEN_8923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8925 = 10'h249 == r_count_11_io_out ? io_r_585_b : _GEN_8924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8926 = 10'h24a == r_count_11_io_out ? io_r_586_b : _GEN_8925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8927 = 10'h24b == r_count_11_io_out ? io_r_587_b : _GEN_8926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8928 = 10'h24c == r_count_11_io_out ? io_r_588_b : _GEN_8927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8929 = 10'h24d == r_count_11_io_out ? io_r_589_b : _GEN_8928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8930 = 10'h24e == r_count_11_io_out ? io_r_590_b : _GEN_8929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8931 = 10'h24f == r_count_11_io_out ? io_r_591_b : _GEN_8930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8932 = 10'h250 == r_count_11_io_out ? io_r_592_b : _GEN_8931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8933 = 10'h251 == r_count_11_io_out ? io_r_593_b : _GEN_8932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8934 = 10'h252 == r_count_11_io_out ? io_r_594_b : _GEN_8933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8935 = 10'h253 == r_count_11_io_out ? io_r_595_b : _GEN_8934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8936 = 10'h254 == r_count_11_io_out ? io_r_596_b : _GEN_8935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8937 = 10'h255 == r_count_11_io_out ? io_r_597_b : _GEN_8936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8938 = 10'h256 == r_count_11_io_out ? io_r_598_b : _GEN_8937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8939 = 10'h257 == r_count_11_io_out ? io_r_599_b : _GEN_8938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8940 = 10'h258 == r_count_11_io_out ? io_r_600_b : _GEN_8939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8941 = 10'h259 == r_count_11_io_out ? io_r_601_b : _GEN_8940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8942 = 10'h25a == r_count_11_io_out ? io_r_602_b : _GEN_8941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8943 = 10'h25b == r_count_11_io_out ? io_r_603_b : _GEN_8942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8944 = 10'h25c == r_count_11_io_out ? io_r_604_b : _GEN_8943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8945 = 10'h25d == r_count_11_io_out ? io_r_605_b : _GEN_8944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8946 = 10'h25e == r_count_11_io_out ? io_r_606_b : _GEN_8945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8947 = 10'h25f == r_count_11_io_out ? io_r_607_b : _GEN_8946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8948 = 10'h260 == r_count_11_io_out ? io_r_608_b : _GEN_8947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8949 = 10'h261 == r_count_11_io_out ? io_r_609_b : _GEN_8948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8950 = 10'h262 == r_count_11_io_out ? io_r_610_b : _GEN_8949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8951 = 10'h263 == r_count_11_io_out ? io_r_611_b : _GEN_8950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8952 = 10'h264 == r_count_11_io_out ? io_r_612_b : _GEN_8951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8953 = 10'h265 == r_count_11_io_out ? io_r_613_b : _GEN_8952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8954 = 10'h266 == r_count_11_io_out ? io_r_614_b : _GEN_8953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8955 = 10'h267 == r_count_11_io_out ? io_r_615_b : _GEN_8954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8956 = 10'h268 == r_count_11_io_out ? io_r_616_b : _GEN_8955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8957 = 10'h269 == r_count_11_io_out ? io_r_617_b : _GEN_8956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8958 = 10'h26a == r_count_11_io_out ? io_r_618_b : _GEN_8957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8959 = 10'h26b == r_count_11_io_out ? io_r_619_b : _GEN_8958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8960 = 10'h26c == r_count_11_io_out ? io_r_620_b : _GEN_8959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8961 = 10'h26d == r_count_11_io_out ? io_r_621_b : _GEN_8960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8962 = 10'h26e == r_count_11_io_out ? io_r_622_b : _GEN_8961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8963 = 10'h26f == r_count_11_io_out ? io_r_623_b : _GEN_8962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8964 = 10'h270 == r_count_11_io_out ? io_r_624_b : _GEN_8963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8965 = 10'h271 == r_count_11_io_out ? io_r_625_b : _GEN_8964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8966 = 10'h272 == r_count_11_io_out ? io_r_626_b : _GEN_8965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8967 = 10'h273 == r_count_11_io_out ? io_r_627_b : _GEN_8966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8968 = 10'h274 == r_count_11_io_out ? io_r_628_b : _GEN_8967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8969 = 10'h275 == r_count_11_io_out ? io_r_629_b : _GEN_8968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8970 = 10'h276 == r_count_11_io_out ? io_r_630_b : _GEN_8969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8971 = 10'h277 == r_count_11_io_out ? io_r_631_b : _GEN_8970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8972 = 10'h278 == r_count_11_io_out ? io_r_632_b : _GEN_8971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8973 = 10'h279 == r_count_11_io_out ? io_r_633_b : _GEN_8972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8974 = 10'h27a == r_count_11_io_out ? io_r_634_b : _GEN_8973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8975 = 10'h27b == r_count_11_io_out ? io_r_635_b : _GEN_8974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8976 = 10'h27c == r_count_11_io_out ? io_r_636_b : _GEN_8975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8977 = 10'h27d == r_count_11_io_out ? io_r_637_b : _GEN_8976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8978 = 10'h27e == r_count_11_io_out ? io_r_638_b : _GEN_8977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8979 = 10'h27f == r_count_11_io_out ? io_r_639_b : _GEN_8978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8980 = 10'h280 == r_count_11_io_out ? io_r_640_b : _GEN_8979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8981 = 10'h281 == r_count_11_io_out ? io_r_641_b : _GEN_8980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8982 = 10'h282 == r_count_11_io_out ? io_r_642_b : _GEN_8981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8983 = 10'h283 == r_count_11_io_out ? io_r_643_b : _GEN_8982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8984 = 10'h284 == r_count_11_io_out ? io_r_644_b : _GEN_8983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8985 = 10'h285 == r_count_11_io_out ? io_r_645_b : _GEN_8984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8986 = 10'h286 == r_count_11_io_out ? io_r_646_b : _GEN_8985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8987 = 10'h287 == r_count_11_io_out ? io_r_647_b : _GEN_8986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8988 = 10'h288 == r_count_11_io_out ? io_r_648_b : _GEN_8987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8989 = 10'h289 == r_count_11_io_out ? io_r_649_b : _GEN_8988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8990 = 10'h28a == r_count_11_io_out ? io_r_650_b : _GEN_8989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8991 = 10'h28b == r_count_11_io_out ? io_r_651_b : _GEN_8990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8992 = 10'h28c == r_count_11_io_out ? io_r_652_b : _GEN_8991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8993 = 10'h28d == r_count_11_io_out ? io_r_653_b : _GEN_8992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8994 = 10'h28e == r_count_11_io_out ? io_r_654_b : _GEN_8993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8995 = 10'h28f == r_count_11_io_out ? io_r_655_b : _GEN_8994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8996 = 10'h290 == r_count_11_io_out ? io_r_656_b : _GEN_8995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8997 = 10'h291 == r_count_11_io_out ? io_r_657_b : _GEN_8996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8998 = 10'h292 == r_count_11_io_out ? io_r_658_b : _GEN_8997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8999 = 10'h293 == r_count_11_io_out ? io_r_659_b : _GEN_8998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9000 = 10'h294 == r_count_11_io_out ? io_r_660_b : _GEN_8999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9001 = 10'h295 == r_count_11_io_out ? io_r_661_b : _GEN_9000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9002 = 10'h296 == r_count_11_io_out ? io_r_662_b : _GEN_9001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9003 = 10'h297 == r_count_11_io_out ? io_r_663_b : _GEN_9002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9004 = 10'h298 == r_count_11_io_out ? io_r_664_b : _GEN_9003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9005 = 10'h299 == r_count_11_io_out ? io_r_665_b : _GEN_9004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9006 = 10'h29a == r_count_11_io_out ? io_r_666_b : _GEN_9005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9007 = 10'h29b == r_count_11_io_out ? io_r_667_b : _GEN_9006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9008 = 10'h29c == r_count_11_io_out ? io_r_668_b : _GEN_9007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9009 = 10'h29d == r_count_11_io_out ? io_r_669_b : _GEN_9008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9010 = 10'h29e == r_count_11_io_out ? io_r_670_b : _GEN_9009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9011 = 10'h29f == r_count_11_io_out ? io_r_671_b : _GEN_9010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9012 = 10'h2a0 == r_count_11_io_out ? io_r_672_b : _GEN_9011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9013 = 10'h2a1 == r_count_11_io_out ? io_r_673_b : _GEN_9012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9014 = 10'h2a2 == r_count_11_io_out ? io_r_674_b : _GEN_9013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9015 = 10'h2a3 == r_count_11_io_out ? io_r_675_b : _GEN_9014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9016 = 10'h2a4 == r_count_11_io_out ? io_r_676_b : _GEN_9015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9017 = 10'h2a5 == r_count_11_io_out ? io_r_677_b : _GEN_9016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9018 = 10'h2a6 == r_count_11_io_out ? io_r_678_b : _GEN_9017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9019 = 10'h2a7 == r_count_11_io_out ? io_r_679_b : _GEN_9018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9020 = 10'h2a8 == r_count_11_io_out ? io_r_680_b : _GEN_9019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9021 = 10'h2a9 == r_count_11_io_out ? io_r_681_b : _GEN_9020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9022 = 10'h2aa == r_count_11_io_out ? io_r_682_b : _GEN_9021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9023 = 10'h2ab == r_count_11_io_out ? io_r_683_b : _GEN_9022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9024 = 10'h2ac == r_count_11_io_out ? io_r_684_b : _GEN_9023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9025 = 10'h2ad == r_count_11_io_out ? io_r_685_b : _GEN_9024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9026 = 10'h2ae == r_count_11_io_out ? io_r_686_b : _GEN_9025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9027 = 10'h2af == r_count_11_io_out ? io_r_687_b : _GEN_9026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9028 = 10'h2b0 == r_count_11_io_out ? io_r_688_b : _GEN_9027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9029 = 10'h2b1 == r_count_11_io_out ? io_r_689_b : _GEN_9028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9030 = 10'h2b2 == r_count_11_io_out ? io_r_690_b : _GEN_9029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9031 = 10'h2b3 == r_count_11_io_out ? io_r_691_b : _GEN_9030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9032 = 10'h2b4 == r_count_11_io_out ? io_r_692_b : _GEN_9031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9033 = 10'h2b5 == r_count_11_io_out ? io_r_693_b : _GEN_9032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9034 = 10'h2b6 == r_count_11_io_out ? io_r_694_b : _GEN_9033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9035 = 10'h2b7 == r_count_11_io_out ? io_r_695_b : _GEN_9034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9036 = 10'h2b8 == r_count_11_io_out ? io_r_696_b : _GEN_9035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9037 = 10'h2b9 == r_count_11_io_out ? io_r_697_b : _GEN_9036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9038 = 10'h2ba == r_count_11_io_out ? io_r_698_b : _GEN_9037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9039 = 10'h2bb == r_count_11_io_out ? io_r_699_b : _GEN_9038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9040 = 10'h2bc == r_count_11_io_out ? io_r_700_b : _GEN_9039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9041 = 10'h2bd == r_count_11_io_out ? io_r_701_b : _GEN_9040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9042 = 10'h2be == r_count_11_io_out ? io_r_702_b : _GEN_9041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9043 = 10'h2bf == r_count_11_io_out ? io_r_703_b : _GEN_9042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9044 = 10'h2c0 == r_count_11_io_out ? io_r_704_b : _GEN_9043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9045 = 10'h2c1 == r_count_11_io_out ? io_r_705_b : _GEN_9044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9046 = 10'h2c2 == r_count_11_io_out ? io_r_706_b : _GEN_9045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9047 = 10'h2c3 == r_count_11_io_out ? io_r_707_b : _GEN_9046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9048 = 10'h2c4 == r_count_11_io_out ? io_r_708_b : _GEN_9047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9049 = 10'h2c5 == r_count_11_io_out ? io_r_709_b : _GEN_9048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9050 = 10'h2c6 == r_count_11_io_out ? io_r_710_b : _GEN_9049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9051 = 10'h2c7 == r_count_11_io_out ? io_r_711_b : _GEN_9050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9052 = 10'h2c8 == r_count_11_io_out ? io_r_712_b : _GEN_9051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9053 = 10'h2c9 == r_count_11_io_out ? io_r_713_b : _GEN_9052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9054 = 10'h2ca == r_count_11_io_out ? io_r_714_b : _GEN_9053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9055 = 10'h2cb == r_count_11_io_out ? io_r_715_b : _GEN_9054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9056 = 10'h2cc == r_count_11_io_out ? io_r_716_b : _GEN_9055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9057 = 10'h2cd == r_count_11_io_out ? io_r_717_b : _GEN_9056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9058 = 10'h2ce == r_count_11_io_out ? io_r_718_b : _GEN_9057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9059 = 10'h2cf == r_count_11_io_out ? io_r_719_b : _GEN_9058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9060 = 10'h2d0 == r_count_11_io_out ? io_r_720_b : _GEN_9059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9061 = 10'h2d1 == r_count_11_io_out ? io_r_721_b : _GEN_9060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9062 = 10'h2d2 == r_count_11_io_out ? io_r_722_b : _GEN_9061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9063 = 10'h2d3 == r_count_11_io_out ? io_r_723_b : _GEN_9062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9064 = 10'h2d4 == r_count_11_io_out ? io_r_724_b : _GEN_9063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9065 = 10'h2d5 == r_count_11_io_out ? io_r_725_b : _GEN_9064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9066 = 10'h2d6 == r_count_11_io_out ? io_r_726_b : _GEN_9065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9067 = 10'h2d7 == r_count_11_io_out ? io_r_727_b : _GEN_9066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9068 = 10'h2d8 == r_count_11_io_out ? io_r_728_b : _GEN_9067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9069 = 10'h2d9 == r_count_11_io_out ? io_r_729_b : _GEN_9068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9070 = 10'h2da == r_count_11_io_out ? io_r_730_b : _GEN_9069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9071 = 10'h2db == r_count_11_io_out ? io_r_731_b : _GEN_9070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9072 = 10'h2dc == r_count_11_io_out ? io_r_732_b : _GEN_9071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9073 = 10'h2dd == r_count_11_io_out ? io_r_733_b : _GEN_9072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9074 = 10'h2de == r_count_11_io_out ? io_r_734_b : _GEN_9073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9075 = 10'h2df == r_count_11_io_out ? io_r_735_b : _GEN_9074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9076 = 10'h2e0 == r_count_11_io_out ? io_r_736_b : _GEN_9075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9077 = 10'h2e1 == r_count_11_io_out ? io_r_737_b : _GEN_9076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9078 = 10'h2e2 == r_count_11_io_out ? io_r_738_b : _GEN_9077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9079 = 10'h2e3 == r_count_11_io_out ? io_r_739_b : _GEN_9078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9080 = 10'h2e4 == r_count_11_io_out ? io_r_740_b : _GEN_9079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9081 = 10'h2e5 == r_count_11_io_out ? io_r_741_b : _GEN_9080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9082 = 10'h2e6 == r_count_11_io_out ? io_r_742_b : _GEN_9081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9083 = 10'h2e7 == r_count_11_io_out ? io_r_743_b : _GEN_9082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9084 = 10'h2e8 == r_count_11_io_out ? io_r_744_b : _GEN_9083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9085 = 10'h2e9 == r_count_11_io_out ? io_r_745_b : _GEN_9084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9086 = 10'h2ea == r_count_11_io_out ? io_r_746_b : _GEN_9085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9087 = 10'h2eb == r_count_11_io_out ? io_r_747_b : _GEN_9086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9088 = 10'h2ec == r_count_11_io_out ? io_r_748_b : _GEN_9087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9091 = 10'h1 == r_count_12_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9092 = 10'h2 == r_count_12_io_out ? io_r_2_b : _GEN_9091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9093 = 10'h3 == r_count_12_io_out ? io_r_3_b : _GEN_9092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9094 = 10'h4 == r_count_12_io_out ? io_r_4_b : _GEN_9093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9095 = 10'h5 == r_count_12_io_out ? io_r_5_b : _GEN_9094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9096 = 10'h6 == r_count_12_io_out ? io_r_6_b : _GEN_9095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9097 = 10'h7 == r_count_12_io_out ? io_r_7_b : _GEN_9096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9098 = 10'h8 == r_count_12_io_out ? io_r_8_b : _GEN_9097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9099 = 10'h9 == r_count_12_io_out ? io_r_9_b : _GEN_9098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9100 = 10'ha == r_count_12_io_out ? io_r_10_b : _GEN_9099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9101 = 10'hb == r_count_12_io_out ? io_r_11_b : _GEN_9100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9102 = 10'hc == r_count_12_io_out ? io_r_12_b : _GEN_9101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9103 = 10'hd == r_count_12_io_out ? io_r_13_b : _GEN_9102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9104 = 10'he == r_count_12_io_out ? io_r_14_b : _GEN_9103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9105 = 10'hf == r_count_12_io_out ? io_r_15_b : _GEN_9104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9106 = 10'h10 == r_count_12_io_out ? io_r_16_b : _GEN_9105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9107 = 10'h11 == r_count_12_io_out ? io_r_17_b : _GEN_9106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9108 = 10'h12 == r_count_12_io_out ? io_r_18_b : _GEN_9107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9109 = 10'h13 == r_count_12_io_out ? io_r_19_b : _GEN_9108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9110 = 10'h14 == r_count_12_io_out ? io_r_20_b : _GEN_9109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9111 = 10'h15 == r_count_12_io_out ? io_r_21_b : _GEN_9110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9112 = 10'h16 == r_count_12_io_out ? io_r_22_b : _GEN_9111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9113 = 10'h17 == r_count_12_io_out ? io_r_23_b : _GEN_9112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9114 = 10'h18 == r_count_12_io_out ? io_r_24_b : _GEN_9113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9115 = 10'h19 == r_count_12_io_out ? io_r_25_b : _GEN_9114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9116 = 10'h1a == r_count_12_io_out ? io_r_26_b : _GEN_9115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9117 = 10'h1b == r_count_12_io_out ? io_r_27_b : _GEN_9116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9118 = 10'h1c == r_count_12_io_out ? io_r_28_b : _GEN_9117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9119 = 10'h1d == r_count_12_io_out ? io_r_29_b : _GEN_9118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9120 = 10'h1e == r_count_12_io_out ? io_r_30_b : _GEN_9119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9121 = 10'h1f == r_count_12_io_out ? io_r_31_b : _GEN_9120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9122 = 10'h20 == r_count_12_io_out ? io_r_32_b : _GEN_9121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9123 = 10'h21 == r_count_12_io_out ? io_r_33_b : _GEN_9122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9124 = 10'h22 == r_count_12_io_out ? io_r_34_b : _GEN_9123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9125 = 10'h23 == r_count_12_io_out ? io_r_35_b : _GEN_9124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9126 = 10'h24 == r_count_12_io_out ? io_r_36_b : _GEN_9125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9127 = 10'h25 == r_count_12_io_out ? io_r_37_b : _GEN_9126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9128 = 10'h26 == r_count_12_io_out ? io_r_38_b : _GEN_9127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9129 = 10'h27 == r_count_12_io_out ? io_r_39_b : _GEN_9128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9130 = 10'h28 == r_count_12_io_out ? io_r_40_b : _GEN_9129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9131 = 10'h29 == r_count_12_io_out ? io_r_41_b : _GEN_9130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9132 = 10'h2a == r_count_12_io_out ? io_r_42_b : _GEN_9131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9133 = 10'h2b == r_count_12_io_out ? io_r_43_b : _GEN_9132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9134 = 10'h2c == r_count_12_io_out ? io_r_44_b : _GEN_9133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9135 = 10'h2d == r_count_12_io_out ? io_r_45_b : _GEN_9134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9136 = 10'h2e == r_count_12_io_out ? io_r_46_b : _GEN_9135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9137 = 10'h2f == r_count_12_io_out ? io_r_47_b : _GEN_9136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9138 = 10'h30 == r_count_12_io_out ? io_r_48_b : _GEN_9137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9139 = 10'h31 == r_count_12_io_out ? io_r_49_b : _GEN_9138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9140 = 10'h32 == r_count_12_io_out ? io_r_50_b : _GEN_9139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9141 = 10'h33 == r_count_12_io_out ? io_r_51_b : _GEN_9140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9142 = 10'h34 == r_count_12_io_out ? io_r_52_b : _GEN_9141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9143 = 10'h35 == r_count_12_io_out ? io_r_53_b : _GEN_9142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9144 = 10'h36 == r_count_12_io_out ? io_r_54_b : _GEN_9143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9145 = 10'h37 == r_count_12_io_out ? io_r_55_b : _GEN_9144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9146 = 10'h38 == r_count_12_io_out ? io_r_56_b : _GEN_9145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9147 = 10'h39 == r_count_12_io_out ? io_r_57_b : _GEN_9146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9148 = 10'h3a == r_count_12_io_out ? io_r_58_b : _GEN_9147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9149 = 10'h3b == r_count_12_io_out ? io_r_59_b : _GEN_9148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9150 = 10'h3c == r_count_12_io_out ? io_r_60_b : _GEN_9149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9151 = 10'h3d == r_count_12_io_out ? io_r_61_b : _GEN_9150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9152 = 10'h3e == r_count_12_io_out ? io_r_62_b : _GEN_9151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9153 = 10'h3f == r_count_12_io_out ? io_r_63_b : _GEN_9152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9154 = 10'h40 == r_count_12_io_out ? io_r_64_b : _GEN_9153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9155 = 10'h41 == r_count_12_io_out ? io_r_65_b : _GEN_9154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9156 = 10'h42 == r_count_12_io_out ? io_r_66_b : _GEN_9155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9157 = 10'h43 == r_count_12_io_out ? io_r_67_b : _GEN_9156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9158 = 10'h44 == r_count_12_io_out ? io_r_68_b : _GEN_9157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9159 = 10'h45 == r_count_12_io_out ? io_r_69_b : _GEN_9158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9160 = 10'h46 == r_count_12_io_out ? io_r_70_b : _GEN_9159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9161 = 10'h47 == r_count_12_io_out ? io_r_71_b : _GEN_9160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9162 = 10'h48 == r_count_12_io_out ? io_r_72_b : _GEN_9161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9163 = 10'h49 == r_count_12_io_out ? io_r_73_b : _GEN_9162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9164 = 10'h4a == r_count_12_io_out ? io_r_74_b : _GEN_9163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9165 = 10'h4b == r_count_12_io_out ? io_r_75_b : _GEN_9164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9166 = 10'h4c == r_count_12_io_out ? io_r_76_b : _GEN_9165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9167 = 10'h4d == r_count_12_io_out ? io_r_77_b : _GEN_9166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9168 = 10'h4e == r_count_12_io_out ? io_r_78_b : _GEN_9167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9169 = 10'h4f == r_count_12_io_out ? io_r_79_b : _GEN_9168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9170 = 10'h50 == r_count_12_io_out ? io_r_80_b : _GEN_9169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9171 = 10'h51 == r_count_12_io_out ? io_r_81_b : _GEN_9170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9172 = 10'h52 == r_count_12_io_out ? io_r_82_b : _GEN_9171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9173 = 10'h53 == r_count_12_io_out ? io_r_83_b : _GEN_9172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9174 = 10'h54 == r_count_12_io_out ? io_r_84_b : _GEN_9173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9175 = 10'h55 == r_count_12_io_out ? io_r_85_b : _GEN_9174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9176 = 10'h56 == r_count_12_io_out ? io_r_86_b : _GEN_9175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9177 = 10'h57 == r_count_12_io_out ? io_r_87_b : _GEN_9176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9178 = 10'h58 == r_count_12_io_out ? io_r_88_b : _GEN_9177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9179 = 10'h59 == r_count_12_io_out ? io_r_89_b : _GEN_9178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9180 = 10'h5a == r_count_12_io_out ? io_r_90_b : _GEN_9179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9181 = 10'h5b == r_count_12_io_out ? io_r_91_b : _GEN_9180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9182 = 10'h5c == r_count_12_io_out ? io_r_92_b : _GEN_9181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9183 = 10'h5d == r_count_12_io_out ? io_r_93_b : _GEN_9182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9184 = 10'h5e == r_count_12_io_out ? io_r_94_b : _GEN_9183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9185 = 10'h5f == r_count_12_io_out ? io_r_95_b : _GEN_9184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9186 = 10'h60 == r_count_12_io_out ? io_r_96_b : _GEN_9185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9187 = 10'h61 == r_count_12_io_out ? io_r_97_b : _GEN_9186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9188 = 10'h62 == r_count_12_io_out ? io_r_98_b : _GEN_9187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9189 = 10'h63 == r_count_12_io_out ? io_r_99_b : _GEN_9188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9190 = 10'h64 == r_count_12_io_out ? io_r_100_b : _GEN_9189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9191 = 10'h65 == r_count_12_io_out ? io_r_101_b : _GEN_9190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9192 = 10'h66 == r_count_12_io_out ? io_r_102_b : _GEN_9191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9193 = 10'h67 == r_count_12_io_out ? io_r_103_b : _GEN_9192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9194 = 10'h68 == r_count_12_io_out ? io_r_104_b : _GEN_9193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9195 = 10'h69 == r_count_12_io_out ? io_r_105_b : _GEN_9194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9196 = 10'h6a == r_count_12_io_out ? io_r_106_b : _GEN_9195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9197 = 10'h6b == r_count_12_io_out ? io_r_107_b : _GEN_9196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9198 = 10'h6c == r_count_12_io_out ? io_r_108_b : _GEN_9197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9199 = 10'h6d == r_count_12_io_out ? io_r_109_b : _GEN_9198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9200 = 10'h6e == r_count_12_io_out ? io_r_110_b : _GEN_9199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9201 = 10'h6f == r_count_12_io_out ? io_r_111_b : _GEN_9200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9202 = 10'h70 == r_count_12_io_out ? io_r_112_b : _GEN_9201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9203 = 10'h71 == r_count_12_io_out ? io_r_113_b : _GEN_9202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9204 = 10'h72 == r_count_12_io_out ? io_r_114_b : _GEN_9203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9205 = 10'h73 == r_count_12_io_out ? io_r_115_b : _GEN_9204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9206 = 10'h74 == r_count_12_io_out ? io_r_116_b : _GEN_9205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9207 = 10'h75 == r_count_12_io_out ? io_r_117_b : _GEN_9206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9208 = 10'h76 == r_count_12_io_out ? io_r_118_b : _GEN_9207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9209 = 10'h77 == r_count_12_io_out ? io_r_119_b : _GEN_9208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9210 = 10'h78 == r_count_12_io_out ? io_r_120_b : _GEN_9209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9211 = 10'h79 == r_count_12_io_out ? io_r_121_b : _GEN_9210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9212 = 10'h7a == r_count_12_io_out ? io_r_122_b : _GEN_9211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9213 = 10'h7b == r_count_12_io_out ? io_r_123_b : _GEN_9212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9214 = 10'h7c == r_count_12_io_out ? io_r_124_b : _GEN_9213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9215 = 10'h7d == r_count_12_io_out ? io_r_125_b : _GEN_9214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9216 = 10'h7e == r_count_12_io_out ? io_r_126_b : _GEN_9215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9217 = 10'h7f == r_count_12_io_out ? io_r_127_b : _GEN_9216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9218 = 10'h80 == r_count_12_io_out ? io_r_128_b : _GEN_9217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9219 = 10'h81 == r_count_12_io_out ? io_r_129_b : _GEN_9218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9220 = 10'h82 == r_count_12_io_out ? io_r_130_b : _GEN_9219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9221 = 10'h83 == r_count_12_io_out ? io_r_131_b : _GEN_9220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9222 = 10'h84 == r_count_12_io_out ? io_r_132_b : _GEN_9221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9223 = 10'h85 == r_count_12_io_out ? io_r_133_b : _GEN_9222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9224 = 10'h86 == r_count_12_io_out ? io_r_134_b : _GEN_9223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9225 = 10'h87 == r_count_12_io_out ? io_r_135_b : _GEN_9224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9226 = 10'h88 == r_count_12_io_out ? io_r_136_b : _GEN_9225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9227 = 10'h89 == r_count_12_io_out ? io_r_137_b : _GEN_9226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9228 = 10'h8a == r_count_12_io_out ? io_r_138_b : _GEN_9227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9229 = 10'h8b == r_count_12_io_out ? io_r_139_b : _GEN_9228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9230 = 10'h8c == r_count_12_io_out ? io_r_140_b : _GEN_9229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9231 = 10'h8d == r_count_12_io_out ? io_r_141_b : _GEN_9230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9232 = 10'h8e == r_count_12_io_out ? io_r_142_b : _GEN_9231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9233 = 10'h8f == r_count_12_io_out ? io_r_143_b : _GEN_9232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9234 = 10'h90 == r_count_12_io_out ? io_r_144_b : _GEN_9233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9235 = 10'h91 == r_count_12_io_out ? io_r_145_b : _GEN_9234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9236 = 10'h92 == r_count_12_io_out ? io_r_146_b : _GEN_9235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9237 = 10'h93 == r_count_12_io_out ? io_r_147_b : _GEN_9236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9238 = 10'h94 == r_count_12_io_out ? io_r_148_b : _GEN_9237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9239 = 10'h95 == r_count_12_io_out ? io_r_149_b : _GEN_9238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9240 = 10'h96 == r_count_12_io_out ? io_r_150_b : _GEN_9239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9241 = 10'h97 == r_count_12_io_out ? io_r_151_b : _GEN_9240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9242 = 10'h98 == r_count_12_io_out ? io_r_152_b : _GEN_9241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9243 = 10'h99 == r_count_12_io_out ? io_r_153_b : _GEN_9242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9244 = 10'h9a == r_count_12_io_out ? io_r_154_b : _GEN_9243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9245 = 10'h9b == r_count_12_io_out ? io_r_155_b : _GEN_9244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9246 = 10'h9c == r_count_12_io_out ? io_r_156_b : _GEN_9245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9247 = 10'h9d == r_count_12_io_out ? io_r_157_b : _GEN_9246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9248 = 10'h9e == r_count_12_io_out ? io_r_158_b : _GEN_9247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9249 = 10'h9f == r_count_12_io_out ? io_r_159_b : _GEN_9248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9250 = 10'ha0 == r_count_12_io_out ? io_r_160_b : _GEN_9249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9251 = 10'ha1 == r_count_12_io_out ? io_r_161_b : _GEN_9250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9252 = 10'ha2 == r_count_12_io_out ? io_r_162_b : _GEN_9251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9253 = 10'ha3 == r_count_12_io_out ? io_r_163_b : _GEN_9252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9254 = 10'ha4 == r_count_12_io_out ? io_r_164_b : _GEN_9253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9255 = 10'ha5 == r_count_12_io_out ? io_r_165_b : _GEN_9254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9256 = 10'ha6 == r_count_12_io_out ? io_r_166_b : _GEN_9255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9257 = 10'ha7 == r_count_12_io_out ? io_r_167_b : _GEN_9256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9258 = 10'ha8 == r_count_12_io_out ? io_r_168_b : _GEN_9257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9259 = 10'ha9 == r_count_12_io_out ? io_r_169_b : _GEN_9258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9260 = 10'haa == r_count_12_io_out ? io_r_170_b : _GEN_9259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9261 = 10'hab == r_count_12_io_out ? io_r_171_b : _GEN_9260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9262 = 10'hac == r_count_12_io_out ? io_r_172_b : _GEN_9261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9263 = 10'had == r_count_12_io_out ? io_r_173_b : _GEN_9262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9264 = 10'hae == r_count_12_io_out ? io_r_174_b : _GEN_9263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9265 = 10'haf == r_count_12_io_out ? io_r_175_b : _GEN_9264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9266 = 10'hb0 == r_count_12_io_out ? io_r_176_b : _GEN_9265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9267 = 10'hb1 == r_count_12_io_out ? io_r_177_b : _GEN_9266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9268 = 10'hb2 == r_count_12_io_out ? io_r_178_b : _GEN_9267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9269 = 10'hb3 == r_count_12_io_out ? io_r_179_b : _GEN_9268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9270 = 10'hb4 == r_count_12_io_out ? io_r_180_b : _GEN_9269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9271 = 10'hb5 == r_count_12_io_out ? io_r_181_b : _GEN_9270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9272 = 10'hb6 == r_count_12_io_out ? io_r_182_b : _GEN_9271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9273 = 10'hb7 == r_count_12_io_out ? io_r_183_b : _GEN_9272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9274 = 10'hb8 == r_count_12_io_out ? io_r_184_b : _GEN_9273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9275 = 10'hb9 == r_count_12_io_out ? io_r_185_b : _GEN_9274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9276 = 10'hba == r_count_12_io_out ? io_r_186_b : _GEN_9275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9277 = 10'hbb == r_count_12_io_out ? io_r_187_b : _GEN_9276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9278 = 10'hbc == r_count_12_io_out ? io_r_188_b : _GEN_9277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9279 = 10'hbd == r_count_12_io_out ? io_r_189_b : _GEN_9278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9280 = 10'hbe == r_count_12_io_out ? io_r_190_b : _GEN_9279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9281 = 10'hbf == r_count_12_io_out ? io_r_191_b : _GEN_9280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9282 = 10'hc0 == r_count_12_io_out ? io_r_192_b : _GEN_9281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9283 = 10'hc1 == r_count_12_io_out ? io_r_193_b : _GEN_9282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9284 = 10'hc2 == r_count_12_io_out ? io_r_194_b : _GEN_9283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9285 = 10'hc3 == r_count_12_io_out ? io_r_195_b : _GEN_9284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9286 = 10'hc4 == r_count_12_io_out ? io_r_196_b : _GEN_9285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9287 = 10'hc5 == r_count_12_io_out ? io_r_197_b : _GEN_9286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9288 = 10'hc6 == r_count_12_io_out ? io_r_198_b : _GEN_9287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9289 = 10'hc7 == r_count_12_io_out ? io_r_199_b : _GEN_9288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9290 = 10'hc8 == r_count_12_io_out ? io_r_200_b : _GEN_9289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9291 = 10'hc9 == r_count_12_io_out ? io_r_201_b : _GEN_9290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9292 = 10'hca == r_count_12_io_out ? io_r_202_b : _GEN_9291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9293 = 10'hcb == r_count_12_io_out ? io_r_203_b : _GEN_9292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9294 = 10'hcc == r_count_12_io_out ? io_r_204_b : _GEN_9293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9295 = 10'hcd == r_count_12_io_out ? io_r_205_b : _GEN_9294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9296 = 10'hce == r_count_12_io_out ? io_r_206_b : _GEN_9295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9297 = 10'hcf == r_count_12_io_out ? io_r_207_b : _GEN_9296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9298 = 10'hd0 == r_count_12_io_out ? io_r_208_b : _GEN_9297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9299 = 10'hd1 == r_count_12_io_out ? io_r_209_b : _GEN_9298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9300 = 10'hd2 == r_count_12_io_out ? io_r_210_b : _GEN_9299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9301 = 10'hd3 == r_count_12_io_out ? io_r_211_b : _GEN_9300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9302 = 10'hd4 == r_count_12_io_out ? io_r_212_b : _GEN_9301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9303 = 10'hd5 == r_count_12_io_out ? io_r_213_b : _GEN_9302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9304 = 10'hd6 == r_count_12_io_out ? io_r_214_b : _GEN_9303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9305 = 10'hd7 == r_count_12_io_out ? io_r_215_b : _GEN_9304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9306 = 10'hd8 == r_count_12_io_out ? io_r_216_b : _GEN_9305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9307 = 10'hd9 == r_count_12_io_out ? io_r_217_b : _GEN_9306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9308 = 10'hda == r_count_12_io_out ? io_r_218_b : _GEN_9307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9309 = 10'hdb == r_count_12_io_out ? io_r_219_b : _GEN_9308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9310 = 10'hdc == r_count_12_io_out ? io_r_220_b : _GEN_9309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9311 = 10'hdd == r_count_12_io_out ? io_r_221_b : _GEN_9310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9312 = 10'hde == r_count_12_io_out ? io_r_222_b : _GEN_9311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9313 = 10'hdf == r_count_12_io_out ? io_r_223_b : _GEN_9312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9314 = 10'he0 == r_count_12_io_out ? io_r_224_b : _GEN_9313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9315 = 10'he1 == r_count_12_io_out ? io_r_225_b : _GEN_9314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9316 = 10'he2 == r_count_12_io_out ? io_r_226_b : _GEN_9315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9317 = 10'he3 == r_count_12_io_out ? io_r_227_b : _GEN_9316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9318 = 10'he4 == r_count_12_io_out ? io_r_228_b : _GEN_9317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9319 = 10'he5 == r_count_12_io_out ? io_r_229_b : _GEN_9318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9320 = 10'he6 == r_count_12_io_out ? io_r_230_b : _GEN_9319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9321 = 10'he7 == r_count_12_io_out ? io_r_231_b : _GEN_9320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9322 = 10'he8 == r_count_12_io_out ? io_r_232_b : _GEN_9321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9323 = 10'he9 == r_count_12_io_out ? io_r_233_b : _GEN_9322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9324 = 10'hea == r_count_12_io_out ? io_r_234_b : _GEN_9323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9325 = 10'heb == r_count_12_io_out ? io_r_235_b : _GEN_9324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9326 = 10'hec == r_count_12_io_out ? io_r_236_b : _GEN_9325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9327 = 10'hed == r_count_12_io_out ? io_r_237_b : _GEN_9326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9328 = 10'hee == r_count_12_io_out ? io_r_238_b : _GEN_9327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9329 = 10'hef == r_count_12_io_out ? io_r_239_b : _GEN_9328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9330 = 10'hf0 == r_count_12_io_out ? io_r_240_b : _GEN_9329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9331 = 10'hf1 == r_count_12_io_out ? io_r_241_b : _GEN_9330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9332 = 10'hf2 == r_count_12_io_out ? io_r_242_b : _GEN_9331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9333 = 10'hf3 == r_count_12_io_out ? io_r_243_b : _GEN_9332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9334 = 10'hf4 == r_count_12_io_out ? io_r_244_b : _GEN_9333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9335 = 10'hf5 == r_count_12_io_out ? io_r_245_b : _GEN_9334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9336 = 10'hf6 == r_count_12_io_out ? io_r_246_b : _GEN_9335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9337 = 10'hf7 == r_count_12_io_out ? io_r_247_b : _GEN_9336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9338 = 10'hf8 == r_count_12_io_out ? io_r_248_b : _GEN_9337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9339 = 10'hf9 == r_count_12_io_out ? io_r_249_b : _GEN_9338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9340 = 10'hfa == r_count_12_io_out ? io_r_250_b : _GEN_9339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9341 = 10'hfb == r_count_12_io_out ? io_r_251_b : _GEN_9340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9342 = 10'hfc == r_count_12_io_out ? io_r_252_b : _GEN_9341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9343 = 10'hfd == r_count_12_io_out ? io_r_253_b : _GEN_9342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9344 = 10'hfe == r_count_12_io_out ? io_r_254_b : _GEN_9343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9345 = 10'hff == r_count_12_io_out ? io_r_255_b : _GEN_9344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9346 = 10'h100 == r_count_12_io_out ? io_r_256_b : _GEN_9345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9347 = 10'h101 == r_count_12_io_out ? io_r_257_b : _GEN_9346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9348 = 10'h102 == r_count_12_io_out ? io_r_258_b : _GEN_9347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9349 = 10'h103 == r_count_12_io_out ? io_r_259_b : _GEN_9348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9350 = 10'h104 == r_count_12_io_out ? io_r_260_b : _GEN_9349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9351 = 10'h105 == r_count_12_io_out ? io_r_261_b : _GEN_9350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9352 = 10'h106 == r_count_12_io_out ? io_r_262_b : _GEN_9351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9353 = 10'h107 == r_count_12_io_out ? io_r_263_b : _GEN_9352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9354 = 10'h108 == r_count_12_io_out ? io_r_264_b : _GEN_9353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9355 = 10'h109 == r_count_12_io_out ? io_r_265_b : _GEN_9354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9356 = 10'h10a == r_count_12_io_out ? io_r_266_b : _GEN_9355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9357 = 10'h10b == r_count_12_io_out ? io_r_267_b : _GEN_9356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9358 = 10'h10c == r_count_12_io_out ? io_r_268_b : _GEN_9357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9359 = 10'h10d == r_count_12_io_out ? io_r_269_b : _GEN_9358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9360 = 10'h10e == r_count_12_io_out ? io_r_270_b : _GEN_9359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9361 = 10'h10f == r_count_12_io_out ? io_r_271_b : _GEN_9360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9362 = 10'h110 == r_count_12_io_out ? io_r_272_b : _GEN_9361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9363 = 10'h111 == r_count_12_io_out ? io_r_273_b : _GEN_9362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9364 = 10'h112 == r_count_12_io_out ? io_r_274_b : _GEN_9363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9365 = 10'h113 == r_count_12_io_out ? io_r_275_b : _GEN_9364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9366 = 10'h114 == r_count_12_io_out ? io_r_276_b : _GEN_9365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9367 = 10'h115 == r_count_12_io_out ? io_r_277_b : _GEN_9366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9368 = 10'h116 == r_count_12_io_out ? io_r_278_b : _GEN_9367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9369 = 10'h117 == r_count_12_io_out ? io_r_279_b : _GEN_9368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9370 = 10'h118 == r_count_12_io_out ? io_r_280_b : _GEN_9369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9371 = 10'h119 == r_count_12_io_out ? io_r_281_b : _GEN_9370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9372 = 10'h11a == r_count_12_io_out ? io_r_282_b : _GEN_9371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9373 = 10'h11b == r_count_12_io_out ? io_r_283_b : _GEN_9372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9374 = 10'h11c == r_count_12_io_out ? io_r_284_b : _GEN_9373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9375 = 10'h11d == r_count_12_io_out ? io_r_285_b : _GEN_9374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9376 = 10'h11e == r_count_12_io_out ? io_r_286_b : _GEN_9375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9377 = 10'h11f == r_count_12_io_out ? io_r_287_b : _GEN_9376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9378 = 10'h120 == r_count_12_io_out ? io_r_288_b : _GEN_9377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9379 = 10'h121 == r_count_12_io_out ? io_r_289_b : _GEN_9378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9380 = 10'h122 == r_count_12_io_out ? io_r_290_b : _GEN_9379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9381 = 10'h123 == r_count_12_io_out ? io_r_291_b : _GEN_9380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9382 = 10'h124 == r_count_12_io_out ? io_r_292_b : _GEN_9381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9383 = 10'h125 == r_count_12_io_out ? io_r_293_b : _GEN_9382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9384 = 10'h126 == r_count_12_io_out ? io_r_294_b : _GEN_9383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9385 = 10'h127 == r_count_12_io_out ? io_r_295_b : _GEN_9384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9386 = 10'h128 == r_count_12_io_out ? io_r_296_b : _GEN_9385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9387 = 10'h129 == r_count_12_io_out ? io_r_297_b : _GEN_9386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9388 = 10'h12a == r_count_12_io_out ? io_r_298_b : _GEN_9387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9389 = 10'h12b == r_count_12_io_out ? io_r_299_b : _GEN_9388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9390 = 10'h12c == r_count_12_io_out ? io_r_300_b : _GEN_9389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9391 = 10'h12d == r_count_12_io_out ? io_r_301_b : _GEN_9390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9392 = 10'h12e == r_count_12_io_out ? io_r_302_b : _GEN_9391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9393 = 10'h12f == r_count_12_io_out ? io_r_303_b : _GEN_9392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9394 = 10'h130 == r_count_12_io_out ? io_r_304_b : _GEN_9393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9395 = 10'h131 == r_count_12_io_out ? io_r_305_b : _GEN_9394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9396 = 10'h132 == r_count_12_io_out ? io_r_306_b : _GEN_9395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9397 = 10'h133 == r_count_12_io_out ? io_r_307_b : _GEN_9396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9398 = 10'h134 == r_count_12_io_out ? io_r_308_b : _GEN_9397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9399 = 10'h135 == r_count_12_io_out ? io_r_309_b : _GEN_9398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9400 = 10'h136 == r_count_12_io_out ? io_r_310_b : _GEN_9399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9401 = 10'h137 == r_count_12_io_out ? io_r_311_b : _GEN_9400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9402 = 10'h138 == r_count_12_io_out ? io_r_312_b : _GEN_9401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9403 = 10'h139 == r_count_12_io_out ? io_r_313_b : _GEN_9402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9404 = 10'h13a == r_count_12_io_out ? io_r_314_b : _GEN_9403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9405 = 10'h13b == r_count_12_io_out ? io_r_315_b : _GEN_9404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9406 = 10'h13c == r_count_12_io_out ? io_r_316_b : _GEN_9405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9407 = 10'h13d == r_count_12_io_out ? io_r_317_b : _GEN_9406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9408 = 10'h13e == r_count_12_io_out ? io_r_318_b : _GEN_9407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9409 = 10'h13f == r_count_12_io_out ? io_r_319_b : _GEN_9408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9410 = 10'h140 == r_count_12_io_out ? io_r_320_b : _GEN_9409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9411 = 10'h141 == r_count_12_io_out ? io_r_321_b : _GEN_9410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9412 = 10'h142 == r_count_12_io_out ? io_r_322_b : _GEN_9411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9413 = 10'h143 == r_count_12_io_out ? io_r_323_b : _GEN_9412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9414 = 10'h144 == r_count_12_io_out ? io_r_324_b : _GEN_9413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9415 = 10'h145 == r_count_12_io_out ? io_r_325_b : _GEN_9414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9416 = 10'h146 == r_count_12_io_out ? io_r_326_b : _GEN_9415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9417 = 10'h147 == r_count_12_io_out ? io_r_327_b : _GEN_9416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9418 = 10'h148 == r_count_12_io_out ? io_r_328_b : _GEN_9417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9419 = 10'h149 == r_count_12_io_out ? io_r_329_b : _GEN_9418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9420 = 10'h14a == r_count_12_io_out ? io_r_330_b : _GEN_9419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9421 = 10'h14b == r_count_12_io_out ? io_r_331_b : _GEN_9420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9422 = 10'h14c == r_count_12_io_out ? io_r_332_b : _GEN_9421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9423 = 10'h14d == r_count_12_io_out ? io_r_333_b : _GEN_9422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9424 = 10'h14e == r_count_12_io_out ? io_r_334_b : _GEN_9423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9425 = 10'h14f == r_count_12_io_out ? io_r_335_b : _GEN_9424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9426 = 10'h150 == r_count_12_io_out ? io_r_336_b : _GEN_9425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9427 = 10'h151 == r_count_12_io_out ? io_r_337_b : _GEN_9426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9428 = 10'h152 == r_count_12_io_out ? io_r_338_b : _GEN_9427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9429 = 10'h153 == r_count_12_io_out ? io_r_339_b : _GEN_9428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9430 = 10'h154 == r_count_12_io_out ? io_r_340_b : _GEN_9429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9431 = 10'h155 == r_count_12_io_out ? io_r_341_b : _GEN_9430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9432 = 10'h156 == r_count_12_io_out ? io_r_342_b : _GEN_9431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9433 = 10'h157 == r_count_12_io_out ? io_r_343_b : _GEN_9432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9434 = 10'h158 == r_count_12_io_out ? io_r_344_b : _GEN_9433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9435 = 10'h159 == r_count_12_io_out ? io_r_345_b : _GEN_9434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9436 = 10'h15a == r_count_12_io_out ? io_r_346_b : _GEN_9435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9437 = 10'h15b == r_count_12_io_out ? io_r_347_b : _GEN_9436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9438 = 10'h15c == r_count_12_io_out ? io_r_348_b : _GEN_9437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9439 = 10'h15d == r_count_12_io_out ? io_r_349_b : _GEN_9438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9440 = 10'h15e == r_count_12_io_out ? io_r_350_b : _GEN_9439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9441 = 10'h15f == r_count_12_io_out ? io_r_351_b : _GEN_9440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9442 = 10'h160 == r_count_12_io_out ? io_r_352_b : _GEN_9441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9443 = 10'h161 == r_count_12_io_out ? io_r_353_b : _GEN_9442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9444 = 10'h162 == r_count_12_io_out ? io_r_354_b : _GEN_9443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9445 = 10'h163 == r_count_12_io_out ? io_r_355_b : _GEN_9444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9446 = 10'h164 == r_count_12_io_out ? io_r_356_b : _GEN_9445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9447 = 10'h165 == r_count_12_io_out ? io_r_357_b : _GEN_9446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9448 = 10'h166 == r_count_12_io_out ? io_r_358_b : _GEN_9447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9449 = 10'h167 == r_count_12_io_out ? io_r_359_b : _GEN_9448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9450 = 10'h168 == r_count_12_io_out ? io_r_360_b : _GEN_9449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9451 = 10'h169 == r_count_12_io_out ? io_r_361_b : _GEN_9450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9452 = 10'h16a == r_count_12_io_out ? io_r_362_b : _GEN_9451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9453 = 10'h16b == r_count_12_io_out ? io_r_363_b : _GEN_9452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9454 = 10'h16c == r_count_12_io_out ? io_r_364_b : _GEN_9453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9455 = 10'h16d == r_count_12_io_out ? io_r_365_b : _GEN_9454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9456 = 10'h16e == r_count_12_io_out ? io_r_366_b : _GEN_9455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9457 = 10'h16f == r_count_12_io_out ? io_r_367_b : _GEN_9456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9458 = 10'h170 == r_count_12_io_out ? io_r_368_b : _GEN_9457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9459 = 10'h171 == r_count_12_io_out ? io_r_369_b : _GEN_9458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9460 = 10'h172 == r_count_12_io_out ? io_r_370_b : _GEN_9459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9461 = 10'h173 == r_count_12_io_out ? io_r_371_b : _GEN_9460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9462 = 10'h174 == r_count_12_io_out ? io_r_372_b : _GEN_9461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9463 = 10'h175 == r_count_12_io_out ? io_r_373_b : _GEN_9462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9464 = 10'h176 == r_count_12_io_out ? io_r_374_b : _GEN_9463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9465 = 10'h177 == r_count_12_io_out ? io_r_375_b : _GEN_9464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9466 = 10'h178 == r_count_12_io_out ? io_r_376_b : _GEN_9465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9467 = 10'h179 == r_count_12_io_out ? io_r_377_b : _GEN_9466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9468 = 10'h17a == r_count_12_io_out ? io_r_378_b : _GEN_9467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9469 = 10'h17b == r_count_12_io_out ? io_r_379_b : _GEN_9468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9470 = 10'h17c == r_count_12_io_out ? io_r_380_b : _GEN_9469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9471 = 10'h17d == r_count_12_io_out ? io_r_381_b : _GEN_9470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9472 = 10'h17e == r_count_12_io_out ? io_r_382_b : _GEN_9471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9473 = 10'h17f == r_count_12_io_out ? io_r_383_b : _GEN_9472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9474 = 10'h180 == r_count_12_io_out ? io_r_384_b : _GEN_9473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9475 = 10'h181 == r_count_12_io_out ? io_r_385_b : _GEN_9474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9476 = 10'h182 == r_count_12_io_out ? io_r_386_b : _GEN_9475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9477 = 10'h183 == r_count_12_io_out ? io_r_387_b : _GEN_9476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9478 = 10'h184 == r_count_12_io_out ? io_r_388_b : _GEN_9477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9479 = 10'h185 == r_count_12_io_out ? io_r_389_b : _GEN_9478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9480 = 10'h186 == r_count_12_io_out ? io_r_390_b : _GEN_9479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9481 = 10'h187 == r_count_12_io_out ? io_r_391_b : _GEN_9480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9482 = 10'h188 == r_count_12_io_out ? io_r_392_b : _GEN_9481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9483 = 10'h189 == r_count_12_io_out ? io_r_393_b : _GEN_9482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9484 = 10'h18a == r_count_12_io_out ? io_r_394_b : _GEN_9483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9485 = 10'h18b == r_count_12_io_out ? io_r_395_b : _GEN_9484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9486 = 10'h18c == r_count_12_io_out ? io_r_396_b : _GEN_9485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9487 = 10'h18d == r_count_12_io_out ? io_r_397_b : _GEN_9486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9488 = 10'h18e == r_count_12_io_out ? io_r_398_b : _GEN_9487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9489 = 10'h18f == r_count_12_io_out ? io_r_399_b : _GEN_9488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9490 = 10'h190 == r_count_12_io_out ? io_r_400_b : _GEN_9489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9491 = 10'h191 == r_count_12_io_out ? io_r_401_b : _GEN_9490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9492 = 10'h192 == r_count_12_io_out ? io_r_402_b : _GEN_9491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9493 = 10'h193 == r_count_12_io_out ? io_r_403_b : _GEN_9492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9494 = 10'h194 == r_count_12_io_out ? io_r_404_b : _GEN_9493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9495 = 10'h195 == r_count_12_io_out ? io_r_405_b : _GEN_9494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9496 = 10'h196 == r_count_12_io_out ? io_r_406_b : _GEN_9495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9497 = 10'h197 == r_count_12_io_out ? io_r_407_b : _GEN_9496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9498 = 10'h198 == r_count_12_io_out ? io_r_408_b : _GEN_9497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9499 = 10'h199 == r_count_12_io_out ? io_r_409_b : _GEN_9498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9500 = 10'h19a == r_count_12_io_out ? io_r_410_b : _GEN_9499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9501 = 10'h19b == r_count_12_io_out ? io_r_411_b : _GEN_9500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9502 = 10'h19c == r_count_12_io_out ? io_r_412_b : _GEN_9501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9503 = 10'h19d == r_count_12_io_out ? io_r_413_b : _GEN_9502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9504 = 10'h19e == r_count_12_io_out ? io_r_414_b : _GEN_9503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9505 = 10'h19f == r_count_12_io_out ? io_r_415_b : _GEN_9504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9506 = 10'h1a0 == r_count_12_io_out ? io_r_416_b : _GEN_9505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9507 = 10'h1a1 == r_count_12_io_out ? io_r_417_b : _GEN_9506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9508 = 10'h1a2 == r_count_12_io_out ? io_r_418_b : _GEN_9507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9509 = 10'h1a3 == r_count_12_io_out ? io_r_419_b : _GEN_9508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9510 = 10'h1a4 == r_count_12_io_out ? io_r_420_b : _GEN_9509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9511 = 10'h1a5 == r_count_12_io_out ? io_r_421_b : _GEN_9510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9512 = 10'h1a6 == r_count_12_io_out ? io_r_422_b : _GEN_9511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9513 = 10'h1a7 == r_count_12_io_out ? io_r_423_b : _GEN_9512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9514 = 10'h1a8 == r_count_12_io_out ? io_r_424_b : _GEN_9513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9515 = 10'h1a9 == r_count_12_io_out ? io_r_425_b : _GEN_9514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9516 = 10'h1aa == r_count_12_io_out ? io_r_426_b : _GEN_9515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9517 = 10'h1ab == r_count_12_io_out ? io_r_427_b : _GEN_9516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9518 = 10'h1ac == r_count_12_io_out ? io_r_428_b : _GEN_9517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9519 = 10'h1ad == r_count_12_io_out ? io_r_429_b : _GEN_9518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9520 = 10'h1ae == r_count_12_io_out ? io_r_430_b : _GEN_9519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9521 = 10'h1af == r_count_12_io_out ? io_r_431_b : _GEN_9520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9522 = 10'h1b0 == r_count_12_io_out ? io_r_432_b : _GEN_9521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9523 = 10'h1b1 == r_count_12_io_out ? io_r_433_b : _GEN_9522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9524 = 10'h1b2 == r_count_12_io_out ? io_r_434_b : _GEN_9523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9525 = 10'h1b3 == r_count_12_io_out ? io_r_435_b : _GEN_9524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9526 = 10'h1b4 == r_count_12_io_out ? io_r_436_b : _GEN_9525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9527 = 10'h1b5 == r_count_12_io_out ? io_r_437_b : _GEN_9526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9528 = 10'h1b6 == r_count_12_io_out ? io_r_438_b : _GEN_9527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9529 = 10'h1b7 == r_count_12_io_out ? io_r_439_b : _GEN_9528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9530 = 10'h1b8 == r_count_12_io_out ? io_r_440_b : _GEN_9529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9531 = 10'h1b9 == r_count_12_io_out ? io_r_441_b : _GEN_9530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9532 = 10'h1ba == r_count_12_io_out ? io_r_442_b : _GEN_9531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9533 = 10'h1bb == r_count_12_io_out ? io_r_443_b : _GEN_9532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9534 = 10'h1bc == r_count_12_io_out ? io_r_444_b : _GEN_9533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9535 = 10'h1bd == r_count_12_io_out ? io_r_445_b : _GEN_9534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9536 = 10'h1be == r_count_12_io_out ? io_r_446_b : _GEN_9535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9537 = 10'h1bf == r_count_12_io_out ? io_r_447_b : _GEN_9536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9538 = 10'h1c0 == r_count_12_io_out ? io_r_448_b : _GEN_9537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9539 = 10'h1c1 == r_count_12_io_out ? io_r_449_b : _GEN_9538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9540 = 10'h1c2 == r_count_12_io_out ? io_r_450_b : _GEN_9539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9541 = 10'h1c3 == r_count_12_io_out ? io_r_451_b : _GEN_9540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9542 = 10'h1c4 == r_count_12_io_out ? io_r_452_b : _GEN_9541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9543 = 10'h1c5 == r_count_12_io_out ? io_r_453_b : _GEN_9542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9544 = 10'h1c6 == r_count_12_io_out ? io_r_454_b : _GEN_9543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9545 = 10'h1c7 == r_count_12_io_out ? io_r_455_b : _GEN_9544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9546 = 10'h1c8 == r_count_12_io_out ? io_r_456_b : _GEN_9545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9547 = 10'h1c9 == r_count_12_io_out ? io_r_457_b : _GEN_9546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9548 = 10'h1ca == r_count_12_io_out ? io_r_458_b : _GEN_9547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9549 = 10'h1cb == r_count_12_io_out ? io_r_459_b : _GEN_9548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9550 = 10'h1cc == r_count_12_io_out ? io_r_460_b : _GEN_9549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9551 = 10'h1cd == r_count_12_io_out ? io_r_461_b : _GEN_9550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9552 = 10'h1ce == r_count_12_io_out ? io_r_462_b : _GEN_9551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9553 = 10'h1cf == r_count_12_io_out ? io_r_463_b : _GEN_9552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9554 = 10'h1d0 == r_count_12_io_out ? io_r_464_b : _GEN_9553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9555 = 10'h1d1 == r_count_12_io_out ? io_r_465_b : _GEN_9554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9556 = 10'h1d2 == r_count_12_io_out ? io_r_466_b : _GEN_9555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9557 = 10'h1d3 == r_count_12_io_out ? io_r_467_b : _GEN_9556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9558 = 10'h1d4 == r_count_12_io_out ? io_r_468_b : _GEN_9557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9559 = 10'h1d5 == r_count_12_io_out ? io_r_469_b : _GEN_9558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9560 = 10'h1d6 == r_count_12_io_out ? io_r_470_b : _GEN_9559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9561 = 10'h1d7 == r_count_12_io_out ? io_r_471_b : _GEN_9560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9562 = 10'h1d8 == r_count_12_io_out ? io_r_472_b : _GEN_9561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9563 = 10'h1d9 == r_count_12_io_out ? io_r_473_b : _GEN_9562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9564 = 10'h1da == r_count_12_io_out ? io_r_474_b : _GEN_9563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9565 = 10'h1db == r_count_12_io_out ? io_r_475_b : _GEN_9564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9566 = 10'h1dc == r_count_12_io_out ? io_r_476_b : _GEN_9565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9567 = 10'h1dd == r_count_12_io_out ? io_r_477_b : _GEN_9566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9568 = 10'h1de == r_count_12_io_out ? io_r_478_b : _GEN_9567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9569 = 10'h1df == r_count_12_io_out ? io_r_479_b : _GEN_9568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9570 = 10'h1e0 == r_count_12_io_out ? io_r_480_b : _GEN_9569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9571 = 10'h1e1 == r_count_12_io_out ? io_r_481_b : _GEN_9570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9572 = 10'h1e2 == r_count_12_io_out ? io_r_482_b : _GEN_9571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9573 = 10'h1e3 == r_count_12_io_out ? io_r_483_b : _GEN_9572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9574 = 10'h1e4 == r_count_12_io_out ? io_r_484_b : _GEN_9573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9575 = 10'h1e5 == r_count_12_io_out ? io_r_485_b : _GEN_9574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9576 = 10'h1e6 == r_count_12_io_out ? io_r_486_b : _GEN_9575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9577 = 10'h1e7 == r_count_12_io_out ? io_r_487_b : _GEN_9576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9578 = 10'h1e8 == r_count_12_io_out ? io_r_488_b : _GEN_9577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9579 = 10'h1e9 == r_count_12_io_out ? io_r_489_b : _GEN_9578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9580 = 10'h1ea == r_count_12_io_out ? io_r_490_b : _GEN_9579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9581 = 10'h1eb == r_count_12_io_out ? io_r_491_b : _GEN_9580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9582 = 10'h1ec == r_count_12_io_out ? io_r_492_b : _GEN_9581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9583 = 10'h1ed == r_count_12_io_out ? io_r_493_b : _GEN_9582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9584 = 10'h1ee == r_count_12_io_out ? io_r_494_b : _GEN_9583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9585 = 10'h1ef == r_count_12_io_out ? io_r_495_b : _GEN_9584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9586 = 10'h1f0 == r_count_12_io_out ? io_r_496_b : _GEN_9585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9587 = 10'h1f1 == r_count_12_io_out ? io_r_497_b : _GEN_9586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9588 = 10'h1f2 == r_count_12_io_out ? io_r_498_b : _GEN_9587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9589 = 10'h1f3 == r_count_12_io_out ? io_r_499_b : _GEN_9588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9590 = 10'h1f4 == r_count_12_io_out ? io_r_500_b : _GEN_9589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9591 = 10'h1f5 == r_count_12_io_out ? io_r_501_b : _GEN_9590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9592 = 10'h1f6 == r_count_12_io_out ? io_r_502_b : _GEN_9591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9593 = 10'h1f7 == r_count_12_io_out ? io_r_503_b : _GEN_9592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9594 = 10'h1f8 == r_count_12_io_out ? io_r_504_b : _GEN_9593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9595 = 10'h1f9 == r_count_12_io_out ? io_r_505_b : _GEN_9594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9596 = 10'h1fa == r_count_12_io_out ? io_r_506_b : _GEN_9595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9597 = 10'h1fb == r_count_12_io_out ? io_r_507_b : _GEN_9596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9598 = 10'h1fc == r_count_12_io_out ? io_r_508_b : _GEN_9597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9599 = 10'h1fd == r_count_12_io_out ? io_r_509_b : _GEN_9598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9600 = 10'h1fe == r_count_12_io_out ? io_r_510_b : _GEN_9599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9601 = 10'h1ff == r_count_12_io_out ? io_r_511_b : _GEN_9600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9602 = 10'h200 == r_count_12_io_out ? io_r_512_b : _GEN_9601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9603 = 10'h201 == r_count_12_io_out ? io_r_513_b : _GEN_9602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9604 = 10'h202 == r_count_12_io_out ? io_r_514_b : _GEN_9603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9605 = 10'h203 == r_count_12_io_out ? io_r_515_b : _GEN_9604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9606 = 10'h204 == r_count_12_io_out ? io_r_516_b : _GEN_9605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9607 = 10'h205 == r_count_12_io_out ? io_r_517_b : _GEN_9606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9608 = 10'h206 == r_count_12_io_out ? io_r_518_b : _GEN_9607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9609 = 10'h207 == r_count_12_io_out ? io_r_519_b : _GEN_9608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9610 = 10'h208 == r_count_12_io_out ? io_r_520_b : _GEN_9609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9611 = 10'h209 == r_count_12_io_out ? io_r_521_b : _GEN_9610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9612 = 10'h20a == r_count_12_io_out ? io_r_522_b : _GEN_9611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9613 = 10'h20b == r_count_12_io_out ? io_r_523_b : _GEN_9612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9614 = 10'h20c == r_count_12_io_out ? io_r_524_b : _GEN_9613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9615 = 10'h20d == r_count_12_io_out ? io_r_525_b : _GEN_9614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9616 = 10'h20e == r_count_12_io_out ? io_r_526_b : _GEN_9615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9617 = 10'h20f == r_count_12_io_out ? io_r_527_b : _GEN_9616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9618 = 10'h210 == r_count_12_io_out ? io_r_528_b : _GEN_9617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9619 = 10'h211 == r_count_12_io_out ? io_r_529_b : _GEN_9618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9620 = 10'h212 == r_count_12_io_out ? io_r_530_b : _GEN_9619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9621 = 10'h213 == r_count_12_io_out ? io_r_531_b : _GEN_9620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9622 = 10'h214 == r_count_12_io_out ? io_r_532_b : _GEN_9621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9623 = 10'h215 == r_count_12_io_out ? io_r_533_b : _GEN_9622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9624 = 10'h216 == r_count_12_io_out ? io_r_534_b : _GEN_9623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9625 = 10'h217 == r_count_12_io_out ? io_r_535_b : _GEN_9624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9626 = 10'h218 == r_count_12_io_out ? io_r_536_b : _GEN_9625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9627 = 10'h219 == r_count_12_io_out ? io_r_537_b : _GEN_9626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9628 = 10'h21a == r_count_12_io_out ? io_r_538_b : _GEN_9627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9629 = 10'h21b == r_count_12_io_out ? io_r_539_b : _GEN_9628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9630 = 10'h21c == r_count_12_io_out ? io_r_540_b : _GEN_9629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9631 = 10'h21d == r_count_12_io_out ? io_r_541_b : _GEN_9630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9632 = 10'h21e == r_count_12_io_out ? io_r_542_b : _GEN_9631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9633 = 10'h21f == r_count_12_io_out ? io_r_543_b : _GEN_9632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9634 = 10'h220 == r_count_12_io_out ? io_r_544_b : _GEN_9633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9635 = 10'h221 == r_count_12_io_out ? io_r_545_b : _GEN_9634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9636 = 10'h222 == r_count_12_io_out ? io_r_546_b : _GEN_9635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9637 = 10'h223 == r_count_12_io_out ? io_r_547_b : _GEN_9636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9638 = 10'h224 == r_count_12_io_out ? io_r_548_b : _GEN_9637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9639 = 10'h225 == r_count_12_io_out ? io_r_549_b : _GEN_9638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9640 = 10'h226 == r_count_12_io_out ? io_r_550_b : _GEN_9639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9641 = 10'h227 == r_count_12_io_out ? io_r_551_b : _GEN_9640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9642 = 10'h228 == r_count_12_io_out ? io_r_552_b : _GEN_9641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9643 = 10'h229 == r_count_12_io_out ? io_r_553_b : _GEN_9642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9644 = 10'h22a == r_count_12_io_out ? io_r_554_b : _GEN_9643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9645 = 10'h22b == r_count_12_io_out ? io_r_555_b : _GEN_9644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9646 = 10'h22c == r_count_12_io_out ? io_r_556_b : _GEN_9645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9647 = 10'h22d == r_count_12_io_out ? io_r_557_b : _GEN_9646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9648 = 10'h22e == r_count_12_io_out ? io_r_558_b : _GEN_9647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9649 = 10'h22f == r_count_12_io_out ? io_r_559_b : _GEN_9648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9650 = 10'h230 == r_count_12_io_out ? io_r_560_b : _GEN_9649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9651 = 10'h231 == r_count_12_io_out ? io_r_561_b : _GEN_9650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9652 = 10'h232 == r_count_12_io_out ? io_r_562_b : _GEN_9651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9653 = 10'h233 == r_count_12_io_out ? io_r_563_b : _GEN_9652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9654 = 10'h234 == r_count_12_io_out ? io_r_564_b : _GEN_9653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9655 = 10'h235 == r_count_12_io_out ? io_r_565_b : _GEN_9654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9656 = 10'h236 == r_count_12_io_out ? io_r_566_b : _GEN_9655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9657 = 10'h237 == r_count_12_io_out ? io_r_567_b : _GEN_9656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9658 = 10'h238 == r_count_12_io_out ? io_r_568_b : _GEN_9657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9659 = 10'h239 == r_count_12_io_out ? io_r_569_b : _GEN_9658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9660 = 10'h23a == r_count_12_io_out ? io_r_570_b : _GEN_9659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9661 = 10'h23b == r_count_12_io_out ? io_r_571_b : _GEN_9660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9662 = 10'h23c == r_count_12_io_out ? io_r_572_b : _GEN_9661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9663 = 10'h23d == r_count_12_io_out ? io_r_573_b : _GEN_9662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9664 = 10'h23e == r_count_12_io_out ? io_r_574_b : _GEN_9663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9665 = 10'h23f == r_count_12_io_out ? io_r_575_b : _GEN_9664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9666 = 10'h240 == r_count_12_io_out ? io_r_576_b : _GEN_9665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9667 = 10'h241 == r_count_12_io_out ? io_r_577_b : _GEN_9666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9668 = 10'h242 == r_count_12_io_out ? io_r_578_b : _GEN_9667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9669 = 10'h243 == r_count_12_io_out ? io_r_579_b : _GEN_9668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9670 = 10'h244 == r_count_12_io_out ? io_r_580_b : _GEN_9669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9671 = 10'h245 == r_count_12_io_out ? io_r_581_b : _GEN_9670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9672 = 10'h246 == r_count_12_io_out ? io_r_582_b : _GEN_9671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9673 = 10'h247 == r_count_12_io_out ? io_r_583_b : _GEN_9672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9674 = 10'h248 == r_count_12_io_out ? io_r_584_b : _GEN_9673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9675 = 10'h249 == r_count_12_io_out ? io_r_585_b : _GEN_9674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9676 = 10'h24a == r_count_12_io_out ? io_r_586_b : _GEN_9675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9677 = 10'h24b == r_count_12_io_out ? io_r_587_b : _GEN_9676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9678 = 10'h24c == r_count_12_io_out ? io_r_588_b : _GEN_9677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9679 = 10'h24d == r_count_12_io_out ? io_r_589_b : _GEN_9678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9680 = 10'h24e == r_count_12_io_out ? io_r_590_b : _GEN_9679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9681 = 10'h24f == r_count_12_io_out ? io_r_591_b : _GEN_9680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9682 = 10'h250 == r_count_12_io_out ? io_r_592_b : _GEN_9681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9683 = 10'h251 == r_count_12_io_out ? io_r_593_b : _GEN_9682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9684 = 10'h252 == r_count_12_io_out ? io_r_594_b : _GEN_9683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9685 = 10'h253 == r_count_12_io_out ? io_r_595_b : _GEN_9684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9686 = 10'h254 == r_count_12_io_out ? io_r_596_b : _GEN_9685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9687 = 10'h255 == r_count_12_io_out ? io_r_597_b : _GEN_9686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9688 = 10'h256 == r_count_12_io_out ? io_r_598_b : _GEN_9687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9689 = 10'h257 == r_count_12_io_out ? io_r_599_b : _GEN_9688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9690 = 10'h258 == r_count_12_io_out ? io_r_600_b : _GEN_9689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9691 = 10'h259 == r_count_12_io_out ? io_r_601_b : _GEN_9690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9692 = 10'h25a == r_count_12_io_out ? io_r_602_b : _GEN_9691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9693 = 10'h25b == r_count_12_io_out ? io_r_603_b : _GEN_9692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9694 = 10'h25c == r_count_12_io_out ? io_r_604_b : _GEN_9693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9695 = 10'h25d == r_count_12_io_out ? io_r_605_b : _GEN_9694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9696 = 10'h25e == r_count_12_io_out ? io_r_606_b : _GEN_9695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9697 = 10'h25f == r_count_12_io_out ? io_r_607_b : _GEN_9696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9698 = 10'h260 == r_count_12_io_out ? io_r_608_b : _GEN_9697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9699 = 10'h261 == r_count_12_io_out ? io_r_609_b : _GEN_9698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9700 = 10'h262 == r_count_12_io_out ? io_r_610_b : _GEN_9699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9701 = 10'h263 == r_count_12_io_out ? io_r_611_b : _GEN_9700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9702 = 10'h264 == r_count_12_io_out ? io_r_612_b : _GEN_9701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9703 = 10'h265 == r_count_12_io_out ? io_r_613_b : _GEN_9702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9704 = 10'h266 == r_count_12_io_out ? io_r_614_b : _GEN_9703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9705 = 10'h267 == r_count_12_io_out ? io_r_615_b : _GEN_9704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9706 = 10'h268 == r_count_12_io_out ? io_r_616_b : _GEN_9705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9707 = 10'h269 == r_count_12_io_out ? io_r_617_b : _GEN_9706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9708 = 10'h26a == r_count_12_io_out ? io_r_618_b : _GEN_9707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9709 = 10'h26b == r_count_12_io_out ? io_r_619_b : _GEN_9708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9710 = 10'h26c == r_count_12_io_out ? io_r_620_b : _GEN_9709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9711 = 10'h26d == r_count_12_io_out ? io_r_621_b : _GEN_9710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9712 = 10'h26e == r_count_12_io_out ? io_r_622_b : _GEN_9711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9713 = 10'h26f == r_count_12_io_out ? io_r_623_b : _GEN_9712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9714 = 10'h270 == r_count_12_io_out ? io_r_624_b : _GEN_9713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9715 = 10'h271 == r_count_12_io_out ? io_r_625_b : _GEN_9714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9716 = 10'h272 == r_count_12_io_out ? io_r_626_b : _GEN_9715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9717 = 10'h273 == r_count_12_io_out ? io_r_627_b : _GEN_9716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9718 = 10'h274 == r_count_12_io_out ? io_r_628_b : _GEN_9717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9719 = 10'h275 == r_count_12_io_out ? io_r_629_b : _GEN_9718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9720 = 10'h276 == r_count_12_io_out ? io_r_630_b : _GEN_9719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9721 = 10'h277 == r_count_12_io_out ? io_r_631_b : _GEN_9720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9722 = 10'h278 == r_count_12_io_out ? io_r_632_b : _GEN_9721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9723 = 10'h279 == r_count_12_io_out ? io_r_633_b : _GEN_9722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9724 = 10'h27a == r_count_12_io_out ? io_r_634_b : _GEN_9723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9725 = 10'h27b == r_count_12_io_out ? io_r_635_b : _GEN_9724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9726 = 10'h27c == r_count_12_io_out ? io_r_636_b : _GEN_9725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9727 = 10'h27d == r_count_12_io_out ? io_r_637_b : _GEN_9726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9728 = 10'h27e == r_count_12_io_out ? io_r_638_b : _GEN_9727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9729 = 10'h27f == r_count_12_io_out ? io_r_639_b : _GEN_9728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9730 = 10'h280 == r_count_12_io_out ? io_r_640_b : _GEN_9729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9731 = 10'h281 == r_count_12_io_out ? io_r_641_b : _GEN_9730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9732 = 10'h282 == r_count_12_io_out ? io_r_642_b : _GEN_9731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9733 = 10'h283 == r_count_12_io_out ? io_r_643_b : _GEN_9732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9734 = 10'h284 == r_count_12_io_out ? io_r_644_b : _GEN_9733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9735 = 10'h285 == r_count_12_io_out ? io_r_645_b : _GEN_9734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9736 = 10'h286 == r_count_12_io_out ? io_r_646_b : _GEN_9735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9737 = 10'h287 == r_count_12_io_out ? io_r_647_b : _GEN_9736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9738 = 10'h288 == r_count_12_io_out ? io_r_648_b : _GEN_9737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9739 = 10'h289 == r_count_12_io_out ? io_r_649_b : _GEN_9738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9740 = 10'h28a == r_count_12_io_out ? io_r_650_b : _GEN_9739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9741 = 10'h28b == r_count_12_io_out ? io_r_651_b : _GEN_9740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9742 = 10'h28c == r_count_12_io_out ? io_r_652_b : _GEN_9741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9743 = 10'h28d == r_count_12_io_out ? io_r_653_b : _GEN_9742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9744 = 10'h28e == r_count_12_io_out ? io_r_654_b : _GEN_9743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9745 = 10'h28f == r_count_12_io_out ? io_r_655_b : _GEN_9744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9746 = 10'h290 == r_count_12_io_out ? io_r_656_b : _GEN_9745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9747 = 10'h291 == r_count_12_io_out ? io_r_657_b : _GEN_9746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9748 = 10'h292 == r_count_12_io_out ? io_r_658_b : _GEN_9747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9749 = 10'h293 == r_count_12_io_out ? io_r_659_b : _GEN_9748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9750 = 10'h294 == r_count_12_io_out ? io_r_660_b : _GEN_9749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9751 = 10'h295 == r_count_12_io_out ? io_r_661_b : _GEN_9750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9752 = 10'h296 == r_count_12_io_out ? io_r_662_b : _GEN_9751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9753 = 10'h297 == r_count_12_io_out ? io_r_663_b : _GEN_9752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9754 = 10'h298 == r_count_12_io_out ? io_r_664_b : _GEN_9753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9755 = 10'h299 == r_count_12_io_out ? io_r_665_b : _GEN_9754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9756 = 10'h29a == r_count_12_io_out ? io_r_666_b : _GEN_9755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9757 = 10'h29b == r_count_12_io_out ? io_r_667_b : _GEN_9756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9758 = 10'h29c == r_count_12_io_out ? io_r_668_b : _GEN_9757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9759 = 10'h29d == r_count_12_io_out ? io_r_669_b : _GEN_9758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9760 = 10'h29e == r_count_12_io_out ? io_r_670_b : _GEN_9759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9761 = 10'h29f == r_count_12_io_out ? io_r_671_b : _GEN_9760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9762 = 10'h2a0 == r_count_12_io_out ? io_r_672_b : _GEN_9761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9763 = 10'h2a1 == r_count_12_io_out ? io_r_673_b : _GEN_9762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9764 = 10'h2a2 == r_count_12_io_out ? io_r_674_b : _GEN_9763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9765 = 10'h2a3 == r_count_12_io_out ? io_r_675_b : _GEN_9764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9766 = 10'h2a4 == r_count_12_io_out ? io_r_676_b : _GEN_9765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9767 = 10'h2a5 == r_count_12_io_out ? io_r_677_b : _GEN_9766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9768 = 10'h2a6 == r_count_12_io_out ? io_r_678_b : _GEN_9767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9769 = 10'h2a7 == r_count_12_io_out ? io_r_679_b : _GEN_9768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9770 = 10'h2a8 == r_count_12_io_out ? io_r_680_b : _GEN_9769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9771 = 10'h2a9 == r_count_12_io_out ? io_r_681_b : _GEN_9770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9772 = 10'h2aa == r_count_12_io_out ? io_r_682_b : _GEN_9771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9773 = 10'h2ab == r_count_12_io_out ? io_r_683_b : _GEN_9772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9774 = 10'h2ac == r_count_12_io_out ? io_r_684_b : _GEN_9773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9775 = 10'h2ad == r_count_12_io_out ? io_r_685_b : _GEN_9774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9776 = 10'h2ae == r_count_12_io_out ? io_r_686_b : _GEN_9775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9777 = 10'h2af == r_count_12_io_out ? io_r_687_b : _GEN_9776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9778 = 10'h2b0 == r_count_12_io_out ? io_r_688_b : _GEN_9777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9779 = 10'h2b1 == r_count_12_io_out ? io_r_689_b : _GEN_9778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9780 = 10'h2b2 == r_count_12_io_out ? io_r_690_b : _GEN_9779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9781 = 10'h2b3 == r_count_12_io_out ? io_r_691_b : _GEN_9780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9782 = 10'h2b4 == r_count_12_io_out ? io_r_692_b : _GEN_9781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9783 = 10'h2b5 == r_count_12_io_out ? io_r_693_b : _GEN_9782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9784 = 10'h2b6 == r_count_12_io_out ? io_r_694_b : _GEN_9783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9785 = 10'h2b7 == r_count_12_io_out ? io_r_695_b : _GEN_9784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9786 = 10'h2b8 == r_count_12_io_out ? io_r_696_b : _GEN_9785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9787 = 10'h2b9 == r_count_12_io_out ? io_r_697_b : _GEN_9786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9788 = 10'h2ba == r_count_12_io_out ? io_r_698_b : _GEN_9787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9789 = 10'h2bb == r_count_12_io_out ? io_r_699_b : _GEN_9788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9790 = 10'h2bc == r_count_12_io_out ? io_r_700_b : _GEN_9789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9791 = 10'h2bd == r_count_12_io_out ? io_r_701_b : _GEN_9790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9792 = 10'h2be == r_count_12_io_out ? io_r_702_b : _GEN_9791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9793 = 10'h2bf == r_count_12_io_out ? io_r_703_b : _GEN_9792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9794 = 10'h2c0 == r_count_12_io_out ? io_r_704_b : _GEN_9793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9795 = 10'h2c1 == r_count_12_io_out ? io_r_705_b : _GEN_9794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9796 = 10'h2c2 == r_count_12_io_out ? io_r_706_b : _GEN_9795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9797 = 10'h2c3 == r_count_12_io_out ? io_r_707_b : _GEN_9796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9798 = 10'h2c4 == r_count_12_io_out ? io_r_708_b : _GEN_9797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9799 = 10'h2c5 == r_count_12_io_out ? io_r_709_b : _GEN_9798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9800 = 10'h2c6 == r_count_12_io_out ? io_r_710_b : _GEN_9799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9801 = 10'h2c7 == r_count_12_io_out ? io_r_711_b : _GEN_9800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9802 = 10'h2c8 == r_count_12_io_out ? io_r_712_b : _GEN_9801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9803 = 10'h2c9 == r_count_12_io_out ? io_r_713_b : _GEN_9802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9804 = 10'h2ca == r_count_12_io_out ? io_r_714_b : _GEN_9803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9805 = 10'h2cb == r_count_12_io_out ? io_r_715_b : _GEN_9804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9806 = 10'h2cc == r_count_12_io_out ? io_r_716_b : _GEN_9805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9807 = 10'h2cd == r_count_12_io_out ? io_r_717_b : _GEN_9806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9808 = 10'h2ce == r_count_12_io_out ? io_r_718_b : _GEN_9807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9809 = 10'h2cf == r_count_12_io_out ? io_r_719_b : _GEN_9808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9810 = 10'h2d0 == r_count_12_io_out ? io_r_720_b : _GEN_9809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9811 = 10'h2d1 == r_count_12_io_out ? io_r_721_b : _GEN_9810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9812 = 10'h2d2 == r_count_12_io_out ? io_r_722_b : _GEN_9811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9813 = 10'h2d3 == r_count_12_io_out ? io_r_723_b : _GEN_9812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9814 = 10'h2d4 == r_count_12_io_out ? io_r_724_b : _GEN_9813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9815 = 10'h2d5 == r_count_12_io_out ? io_r_725_b : _GEN_9814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9816 = 10'h2d6 == r_count_12_io_out ? io_r_726_b : _GEN_9815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9817 = 10'h2d7 == r_count_12_io_out ? io_r_727_b : _GEN_9816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9818 = 10'h2d8 == r_count_12_io_out ? io_r_728_b : _GEN_9817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9819 = 10'h2d9 == r_count_12_io_out ? io_r_729_b : _GEN_9818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9820 = 10'h2da == r_count_12_io_out ? io_r_730_b : _GEN_9819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9821 = 10'h2db == r_count_12_io_out ? io_r_731_b : _GEN_9820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9822 = 10'h2dc == r_count_12_io_out ? io_r_732_b : _GEN_9821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9823 = 10'h2dd == r_count_12_io_out ? io_r_733_b : _GEN_9822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9824 = 10'h2de == r_count_12_io_out ? io_r_734_b : _GEN_9823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9825 = 10'h2df == r_count_12_io_out ? io_r_735_b : _GEN_9824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9826 = 10'h2e0 == r_count_12_io_out ? io_r_736_b : _GEN_9825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9827 = 10'h2e1 == r_count_12_io_out ? io_r_737_b : _GEN_9826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9828 = 10'h2e2 == r_count_12_io_out ? io_r_738_b : _GEN_9827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9829 = 10'h2e3 == r_count_12_io_out ? io_r_739_b : _GEN_9828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9830 = 10'h2e4 == r_count_12_io_out ? io_r_740_b : _GEN_9829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9831 = 10'h2e5 == r_count_12_io_out ? io_r_741_b : _GEN_9830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9832 = 10'h2e6 == r_count_12_io_out ? io_r_742_b : _GEN_9831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9833 = 10'h2e7 == r_count_12_io_out ? io_r_743_b : _GEN_9832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9834 = 10'h2e8 == r_count_12_io_out ? io_r_744_b : _GEN_9833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9835 = 10'h2e9 == r_count_12_io_out ? io_r_745_b : _GEN_9834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9836 = 10'h2ea == r_count_12_io_out ? io_r_746_b : _GEN_9835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9837 = 10'h2eb == r_count_12_io_out ? io_r_747_b : _GEN_9836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9838 = 10'h2ec == r_count_12_io_out ? io_r_748_b : _GEN_9837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9841 = 10'h1 == r_count_13_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9842 = 10'h2 == r_count_13_io_out ? io_r_2_b : _GEN_9841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9843 = 10'h3 == r_count_13_io_out ? io_r_3_b : _GEN_9842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9844 = 10'h4 == r_count_13_io_out ? io_r_4_b : _GEN_9843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9845 = 10'h5 == r_count_13_io_out ? io_r_5_b : _GEN_9844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9846 = 10'h6 == r_count_13_io_out ? io_r_6_b : _GEN_9845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9847 = 10'h7 == r_count_13_io_out ? io_r_7_b : _GEN_9846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9848 = 10'h8 == r_count_13_io_out ? io_r_8_b : _GEN_9847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9849 = 10'h9 == r_count_13_io_out ? io_r_9_b : _GEN_9848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9850 = 10'ha == r_count_13_io_out ? io_r_10_b : _GEN_9849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9851 = 10'hb == r_count_13_io_out ? io_r_11_b : _GEN_9850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9852 = 10'hc == r_count_13_io_out ? io_r_12_b : _GEN_9851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9853 = 10'hd == r_count_13_io_out ? io_r_13_b : _GEN_9852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9854 = 10'he == r_count_13_io_out ? io_r_14_b : _GEN_9853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9855 = 10'hf == r_count_13_io_out ? io_r_15_b : _GEN_9854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9856 = 10'h10 == r_count_13_io_out ? io_r_16_b : _GEN_9855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9857 = 10'h11 == r_count_13_io_out ? io_r_17_b : _GEN_9856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9858 = 10'h12 == r_count_13_io_out ? io_r_18_b : _GEN_9857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9859 = 10'h13 == r_count_13_io_out ? io_r_19_b : _GEN_9858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9860 = 10'h14 == r_count_13_io_out ? io_r_20_b : _GEN_9859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9861 = 10'h15 == r_count_13_io_out ? io_r_21_b : _GEN_9860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9862 = 10'h16 == r_count_13_io_out ? io_r_22_b : _GEN_9861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9863 = 10'h17 == r_count_13_io_out ? io_r_23_b : _GEN_9862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9864 = 10'h18 == r_count_13_io_out ? io_r_24_b : _GEN_9863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9865 = 10'h19 == r_count_13_io_out ? io_r_25_b : _GEN_9864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9866 = 10'h1a == r_count_13_io_out ? io_r_26_b : _GEN_9865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9867 = 10'h1b == r_count_13_io_out ? io_r_27_b : _GEN_9866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9868 = 10'h1c == r_count_13_io_out ? io_r_28_b : _GEN_9867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9869 = 10'h1d == r_count_13_io_out ? io_r_29_b : _GEN_9868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9870 = 10'h1e == r_count_13_io_out ? io_r_30_b : _GEN_9869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9871 = 10'h1f == r_count_13_io_out ? io_r_31_b : _GEN_9870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9872 = 10'h20 == r_count_13_io_out ? io_r_32_b : _GEN_9871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9873 = 10'h21 == r_count_13_io_out ? io_r_33_b : _GEN_9872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9874 = 10'h22 == r_count_13_io_out ? io_r_34_b : _GEN_9873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9875 = 10'h23 == r_count_13_io_out ? io_r_35_b : _GEN_9874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9876 = 10'h24 == r_count_13_io_out ? io_r_36_b : _GEN_9875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9877 = 10'h25 == r_count_13_io_out ? io_r_37_b : _GEN_9876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9878 = 10'h26 == r_count_13_io_out ? io_r_38_b : _GEN_9877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9879 = 10'h27 == r_count_13_io_out ? io_r_39_b : _GEN_9878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9880 = 10'h28 == r_count_13_io_out ? io_r_40_b : _GEN_9879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9881 = 10'h29 == r_count_13_io_out ? io_r_41_b : _GEN_9880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9882 = 10'h2a == r_count_13_io_out ? io_r_42_b : _GEN_9881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9883 = 10'h2b == r_count_13_io_out ? io_r_43_b : _GEN_9882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9884 = 10'h2c == r_count_13_io_out ? io_r_44_b : _GEN_9883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9885 = 10'h2d == r_count_13_io_out ? io_r_45_b : _GEN_9884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9886 = 10'h2e == r_count_13_io_out ? io_r_46_b : _GEN_9885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9887 = 10'h2f == r_count_13_io_out ? io_r_47_b : _GEN_9886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9888 = 10'h30 == r_count_13_io_out ? io_r_48_b : _GEN_9887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9889 = 10'h31 == r_count_13_io_out ? io_r_49_b : _GEN_9888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9890 = 10'h32 == r_count_13_io_out ? io_r_50_b : _GEN_9889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9891 = 10'h33 == r_count_13_io_out ? io_r_51_b : _GEN_9890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9892 = 10'h34 == r_count_13_io_out ? io_r_52_b : _GEN_9891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9893 = 10'h35 == r_count_13_io_out ? io_r_53_b : _GEN_9892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9894 = 10'h36 == r_count_13_io_out ? io_r_54_b : _GEN_9893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9895 = 10'h37 == r_count_13_io_out ? io_r_55_b : _GEN_9894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9896 = 10'h38 == r_count_13_io_out ? io_r_56_b : _GEN_9895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9897 = 10'h39 == r_count_13_io_out ? io_r_57_b : _GEN_9896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9898 = 10'h3a == r_count_13_io_out ? io_r_58_b : _GEN_9897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9899 = 10'h3b == r_count_13_io_out ? io_r_59_b : _GEN_9898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9900 = 10'h3c == r_count_13_io_out ? io_r_60_b : _GEN_9899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9901 = 10'h3d == r_count_13_io_out ? io_r_61_b : _GEN_9900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9902 = 10'h3e == r_count_13_io_out ? io_r_62_b : _GEN_9901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9903 = 10'h3f == r_count_13_io_out ? io_r_63_b : _GEN_9902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9904 = 10'h40 == r_count_13_io_out ? io_r_64_b : _GEN_9903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9905 = 10'h41 == r_count_13_io_out ? io_r_65_b : _GEN_9904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9906 = 10'h42 == r_count_13_io_out ? io_r_66_b : _GEN_9905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9907 = 10'h43 == r_count_13_io_out ? io_r_67_b : _GEN_9906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9908 = 10'h44 == r_count_13_io_out ? io_r_68_b : _GEN_9907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9909 = 10'h45 == r_count_13_io_out ? io_r_69_b : _GEN_9908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9910 = 10'h46 == r_count_13_io_out ? io_r_70_b : _GEN_9909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9911 = 10'h47 == r_count_13_io_out ? io_r_71_b : _GEN_9910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9912 = 10'h48 == r_count_13_io_out ? io_r_72_b : _GEN_9911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9913 = 10'h49 == r_count_13_io_out ? io_r_73_b : _GEN_9912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9914 = 10'h4a == r_count_13_io_out ? io_r_74_b : _GEN_9913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9915 = 10'h4b == r_count_13_io_out ? io_r_75_b : _GEN_9914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9916 = 10'h4c == r_count_13_io_out ? io_r_76_b : _GEN_9915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9917 = 10'h4d == r_count_13_io_out ? io_r_77_b : _GEN_9916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9918 = 10'h4e == r_count_13_io_out ? io_r_78_b : _GEN_9917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9919 = 10'h4f == r_count_13_io_out ? io_r_79_b : _GEN_9918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9920 = 10'h50 == r_count_13_io_out ? io_r_80_b : _GEN_9919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9921 = 10'h51 == r_count_13_io_out ? io_r_81_b : _GEN_9920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9922 = 10'h52 == r_count_13_io_out ? io_r_82_b : _GEN_9921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9923 = 10'h53 == r_count_13_io_out ? io_r_83_b : _GEN_9922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9924 = 10'h54 == r_count_13_io_out ? io_r_84_b : _GEN_9923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9925 = 10'h55 == r_count_13_io_out ? io_r_85_b : _GEN_9924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9926 = 10'h56 == r_count_13_io_out ? io_r_86_b : _GEN_9925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9927 = 10'h57 == r_count_13_io_out ? io_r_87_b : _GEN_9926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9928 = 10'h58 == r_count_13_io_out ? io_r_88_b : _GEN_9927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9929 = 10'h59 == r_count_13_io_out ? io_r_89_b : _GEN_9928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9930 = 10'h5a == r_count_13_io_out ? io_r_90_b : _GEN_9929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9931 = 10'h5b == r_count_13_io_out ? io_r_91_b : _GEN_9930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9932 = 10'h5c == r_count_13_io_out ? io_r_92_b : _GEN_9931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9933 = 10'h5d == r_count_13_io_out ? io_r_93_b : _GEN_9932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9934 = 10'h5e == r_count_13_io_out ? io_r_94_b : _GEN_9933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9935 = 10'h5f == r_count_13_io_out ? io_r_95_b : _GEN_9934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9936 = 10'h60 == r_count_13_io_out ? io_r_96_b : _GEN_9935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9937 = 10'h61 == r_count_13_io_out ? io_r_97_b : _GEN_9936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9938 = 10'h62 == r_count_13_io_out ? io_r_98_b : _GEN_9937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9939 = 10'h63 == r_count_13_io_out ? io_r_99_b : _GEN_9938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9940 = 10'h64 == r_count_13_io_out ? io_r_100_b : _GEN_9939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9941 = 10'h65 == r_count_13_io_out ? io_r_101_b : _GEN_9940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9942 = 10'h66 == r_count_13_io_out ? io_r_102_b : _GEN_9941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9943 = 10'h67 == r_count_13_io_out ? io_r_103_b : _GEN_9942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9944 = 10'h68 == r_count_13_io_out ? io_r_104_b : _GEN_9943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9945 = 10'h69 == r_count_13_io_out ? io_r_105_b : _GEN_9944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9946 = 10'h6a == r_count_13_io_out ? io_r_106_b : _GEN_9945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9947 = 10'h6b == r_count_13_io_out ? io_r_107_b : _GEN_9946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9948 = 10'h6c == r_count_13_io_out ? io_r_108_b : _GEN_9947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9949 = 10'h6d == r_count_13_io_out ? io_r_109_b : _GEN_9948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9950 = 10'h6e == r_count_13_io_out ? io_r_110_b : _GEN_9949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9951 = 10'h6f == r_count_13_io_out ? io_r_111_b : _GEN_9950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9952 = 10'h70 == r_count_13_io_out ? io_r_112_b : _GEN_9951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9953 = 10'h71 == r_count_13_io_out ? io_r_113_b : _GEN_9952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9954 = 10'h72 == r_count_13_io_out ? io_r_114_b : _GEN_9953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9955 = 10'h73 == r_count_13_io_out ? io_r_115_b : _GEN_9954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9956 = 10'h74 == r_count_13_io_out ? io_r_116_b : _GEN_9955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9957 = 10'h75 == r_count_13_io_out ? io_r_117_b : _GEN_9956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9958 = 10'h76 == r_count_13_io_out ? io_r_118_b : _GEN_9957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9959 = 10'h77 == r_count_13_io_out ? io_r_119_b : _GEN_9958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9960 = 10'h78 == r_count_13_io_out ? io_r_120_b : _GEN_9959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9961 = 10'h79 == r_count_13_io_out ? io_r_121_b : _GEN_9960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9962 = 10'h7a == r_count_13_io_out ? io_r_122_b : _GEN_9961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9963 = 10'h7b == r_count_13_io_out ? io_r_123_b : _GEN_9962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9964 = 10'h7c == r_count_13_io_out ? io_r_124_b : _GEN_9963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9965 = 10'h7d == r_count_13_io_out ? io_r_125_b : _GEN_9964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9966 = 10'h7e == r_count_13_io_out ? io_r_126_b : _GEN_9965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9967 = 10'h7f == r_count_13_io_out ? io_r_127_b : _GEN_9966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9968 = 10'h80 == r_count_13_io_out ? io_r_128_b : _GEN_9967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9969 = 10'h81 == r_count_13_io_out ? io_r_129_b : _GEN_9968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9970 = 10'h82 == r_count_13_io_out ? io_r_130_b : _GEN_9969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9971 = 10'h83 == r_count_13_io_out ? io_r_131_b : _GEN_9970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9972 = 10'h84 == r_count_13_io_out ? io_r_132_b : _GEN_9971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9973 = 10'h85 == r_count_13_io_out ? io_r_133_b : _GEN_9972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9974 = 10'h86 == r_count_13_io_out ? io_r_134_b : _GEN_9973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9975 = 10'h87 == r_count_13_io_out ? io_r_135_b : _GEN_9974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9976 = 10'h88 == r_count_13_io_out ? io_r_136_b : _GEN_9975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9977 = 10'h89 == r_count_13_io_out ? io_r_137_b : _GEN_9976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9978 = 10'h8a == r_count_13_io_out ? io_r_138_b : _GEN_9977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9979 = 10'h8b == r_count_13_io_out ? io_r_139_b : _GEN_9978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9980 = 10'h8c == r_count_13_io_out ? io_r_140_b : _GEN_9979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9981 = 10'h8d == r_count_13_io_out ? io_r_141_b : _GEN_9980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9982 = 10'h8e == r_count_13_io_out ? io_r_142_b : _GEN_9981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9983 = 10'h8f == r_count_13_io_out ? io_r_143_b : _GEN_9982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9984 = 10'h90 == r_count_13_io_out ? io_r_144_b : _GEN_9983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9985 = 10'h91 == r_count_13_io_out ? io_r_145_b : _GEN_9984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9986 = 10'h92 == r_count_13_io_out ? io_r_146_b : _GEN_9985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9987 = 10'h93 == r_count_13_io_out ? io_r_147_b : _GEN_9986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9988 = 10'h94 == r_count_13_io_out ? io_r_148_b : _GEN_9987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9989 = 10'h95 == r_count_13_io_out ? io_r_149_b : _GEN_9988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9990 = 10'h96 == r_count_13_io_out ? io_r_150_b : _GEN_9989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9991 = 10'h97 == r_count_13_io_out ? io_r_151_b : _GEN_9990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9992 = 10'h98 == r_count_13_io_out ? io_r_152_b : _GEN_9991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9993 = 10'h99 == r_count_13_io_out ? io_r_153_b : _GEN_9992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9994 = 10'h9a == r_count_13_io_out ? io_r_154_b : _GEN_9993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9995 = 10'h9b == r_count_13_io_out ? io_r_155_b : _GEN_9994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9996 = 10'h9c == r_count_13_io_out ? io_r_156_b : _GEN_9995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9997 = 10'h9d == r_count_13_io_out ? io_r_157_b : _GEN_9996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9998 = 10'h9e == r_count_13_io_out ? io_r_158_b : _GEN_9997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9999 = 10'h9f == r_count_13_io_out ? io_r_159_b : _GEN_9998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10000 = 10'ha0 == r_count_13_io_out ? io_r_160_b : _GEN_9999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10001 = 10'ha1 == r_count_13_io_out ? io_r_161_b : _GEN_10000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10002 = 10'ha2 == r_count_13_io_out ? io_r_162_b : _GEN_10001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10003 = 10'ha3 == r_count_13_io_out ? io_r_163_b : _GEN_10002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10004 = 10'ha4 == r_count_13_io_out ? io_r_164_b : _GEN_10003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10005 = 10'ha5 == r_count_13_io_out ? io_r_165_b : _GEN_10004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10006 = 10'ha6 == r_count_13_io_out ? io_r_166_b : _GEN_10005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10007 = 10'ha7 == r_count_13_io_out ? io_r_167_b : _GEN_10006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10008 = 10'ha8 == r_count_13_io_out ? io_r_168_b : _GEN_10007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10009 = 10'ha9 == r_count_13_io_out ? io_r_169_b : _GEN_10008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10010 = 10'haa == r_count_13_io_out ? io_r_170_b : _GEN_10009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10011 = 10'hab == r_count_13_io_out ? io_r_171_b : _GEN_10010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10012 = 10'hac == r_count_13_io_out ? io_r_172_b : _GEN_10011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10013 = 10'had == r_count_13_io_out ? io_r_173_b : _GEN_10012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10014 = 10'hae == r_count_13_io_out ? io_r_174_b : _GEN_10013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10015 = 10'haf == r_count_13_io_out ? io_r_175_b : _GEN_10014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10016 = 10'hb0 == r_count_13_io_out ? io_r_176_b : _GEN_10015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10017 = 10'hb1 == r_count_13_io_out ? io_r_177_b : _GEN_10016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10018 = 10'hb2 == r_count_13_io_out ? io_r_178_b : _GEN_10017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10019 = 10'hb3 == r_count_13_io_out ? io_r_179_b : _GEN_10018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10020 = 10'hb4 == r_count_13_io_out ? io_r_180_b : _GEN_10019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10021 = 10'hb5 == r_count_13_io_out ? io_r_181_b : _GEN_10020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10022 = 10'hb6 == r_count_13_io_out ? io_r_182_b : _GEN_10021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10023 = 10'hb7 == r_count_13_io_out ? io_r_183_b : _GEN_10022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10024 = 10'hb8 == r_count_13_io_out ? io_r_184_b : _GEN_10023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10025 = 10'hb9 == r_count_13_io_out ? io_r_185_b : _GEN_10024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10026 = 10'hba == r_count_13_io_out ? io_r_186_b : _GEN_10025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10027 = 10'hbb == r_count_13_io_out ? io_r_187_b : _GEN_10026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10028 = 10'hbc == r_count_13_io_out ? io_r_188_b : _GEN_10027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10029 = 10'hbd == r_count_13_io_out ? io_r_189_b : _GEN_10028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10030 = 10'hbe == r_count_13_io_out ? io_r_190_b : _GEN_10029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10031 = 10'hbf == r_count_13_io_out ? io_r_191_b : _GEN_10030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10032 = 10'hc0 == r_count_13_io_out ? io_r_192_b : _GEN_10031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10033 = 10'hc1 == r_count_13_io_out ? io_r_193_b : _GEN_10032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10034 = 10'hc2 == r_count_13_io_out ? io_r_194_b : _GEN_10033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10035 = 10'hc3 == r_count_13_io_out ? io_r_195_b : _GEN_10034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10036 = 10'hc4 == r_count_13_io_out ? io_r_196_b : _GEN_10035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10037 = 10'hc5 == r_count_13_io_out ? io_r_197_b : _GEN_10036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10038 = 10'hc6 == r_count_13_io_out ? io_r_198_b : _GEN_10037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10039 = 10'hc7 == r_count_13_io_out ? io_r_199_b : _GEN_10038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10040 = 10'hc8 == r_count_13_io_out ? io_r_200_b : _GEN_10039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10041 = 10'hc9 == r_count_13_io_out ? io_r_201_b : _GEN_10040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10042 = 10'hca == r_count_13_io_out ? io_r_202_b : _GEN_10041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10043 = 10'hcb == r_count_13_io_out ? io_r_203_b : _GEN_10042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10044 = 10'hcc == r_count_13_io_out ? io_r_204_b : _GEN_10043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10045 = 10'hcd == r_count_13_io_out ? io_r_205_b : _GEN_10044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10046 = 10'hce == r_count_13_io_out ? io_r_206_b : _GEN_10045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10047 = 10'hcf == r_count_13_io_out ? io_r_207_b : _GEN_10046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10048 = 10'hd0 == r_count_13_io_out ? io_r_208_b : _GEN_10047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10049 = 10'hd1 == r_count_13_io_out ? io_r_209_b : _GEN_10048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10050 = 10'hd2 == r_count_13_io_out ? io_r_210_b : _GEN_10049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10051 = 10'hd3 == r_count_13_io_out ? io_r_211_b : _GEN_10050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10052 = 10'hd4 == r_count_13_io_out ? io_r_212_b : _GEN_10051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10053 = 10'hd5 == r_count_13_io_out ? io_r_213_b : _GEN_10052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10054 = 10'hd6 == r_count_13_io_out ? io_r_214_b : _GEN_10053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10055 = 10'hd7 == r_count_13_io_out ? io_r_215_b : _GEN_10054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10056 = 10'hd8 == r_count_13_io_out ? io_r_216_b : _GEN_10055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10057 = 10'hd9 == r_count_13_io_out ? io_r_217_b : _GEN_10056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10058 = 10'hda == r_count_13_io_out ? io_r_218_b : _GEN_10057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10059 = 10'hdb == r_count_13_io_out ? io_r_219_b : _GEN_10058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10060 = 10'hdc == r_count_13_io_out ? io_r_220_b : _GEN_10059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10061 = 10'hdd == r_count_13_io_out ? io_r_221_b : _GEN_10060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10062 = 10'hde == r_count_13_io_out ? io_r_222_b : _GEN_10061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10063 = 10'hdf == r_count_13_io_out ? io_r_223_b : _GEN_10062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10064 = 10'he0 == r_count_13_io_out ? io_r_224_b : _GEN_10063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10065 = 10'he1 == r_count_13_io_out ? io_r_225_b : _GEN_10064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10066 = 10'he2 == r_count_13_io_out ? io_r_226_b : _GEN_10065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10067 = 10'he3 == r_count_13_io_out ? io_r_227_b : _GEN_10066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10068 = 10'he4 == r_count_13_io_out ? io_r_228_b : _GEN_10067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10069 = 10'he5 == r_count_13_io_out ? io_r_229_b : _GEN_10068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10070 = 10'he6 == r_count_13_io_out ? io_r_230_b : _GEN_10069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10071 = 10'he7 == r_count_13_io_out ? io_r_231_b : _GEN_10070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10072 = 10'he8 == r_count_13_io_out ? io_r_232_b : _GEN_10071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10073 = 10'he9 == r_count_13_io_out ? io_r_233_b : _GEN_10072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10074 = 10'hea == r_count_13_io_out ? io_r_234_b : _GEN_10073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10075 = 10'heb == r_count_13_io_out ? io_r_235_b : _GEN_10074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10076 = 10'hec == r_count_13_io_out ? io_r_236_b : _GEN_10075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10077 = 10'hed == r_count_13_io_out ? io_r_237_b : _GEN_10076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10078 = 10'hee == r_count_13_io_out ? io_r_238_b : _GEN_10077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10079 = 10'hef == r_count_13_io_out ? io_r_239_b : _GEN_10078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10080 = 10'hf0 == r_count_13_io_out ? io_r_240_b : _GEN_10079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10081 = 10'hf1 == r_count_13_io_out ? io_r_241_b : _GEN_10080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10082 = 10'hf2 == r_count_13_io_out ? io_r_242_b : _GEN_10081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10083 = 10'hf3 == r_count_13_io_out ? io_r_243_b : _GEN_10082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10084 = 10'hf4 == r_count_13_io_out ? io_r_244_b : _GEN_10083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10085 = 10'hf5 == r_count_13_io_out ? io_r_245_b : _GEN_10084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10086 = 10'hf6 == r_count_13_io_out ? io_r_246_b : _GEN_10085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10087 = 10'hf7 == r_count_13_io_out ? io_r_247_b : _GEN_10086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10088 = 10'hf8 == r_count_13_io_out ? io_r_248_b : _GEN_10087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10089 = 10'hf9 == r_count_13_io_out ? io_r_249_b : _GEN_10088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10090 = 10'hfa == r_count_13_io_out ? io_r_250_b : _GEN_10089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10091 = 10'hfb == r_count_13_io_out ? io_r_251_b : _GEN_10090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10092 = 10'hfc == r_count_13_io_out ? io_r_252_b : _GEN_10091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10093 = 10'hfd == r_count_13_io_out ? io_r_253_b : _GEN_10092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10094 = 10'hfe == r_count_13_io_out ? io_r_254_b : _GEN_10093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10095 = 10'hff == r_count_13_io_out ? io_r_255_b : _GEN_10094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10096 = 10'h100 == r_count_13_io_out ? io_r_256_b : _GEN_10095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10097 = 10'h101 == r_count_13_io_out ? io_r_257_b : _GEN_10096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10098 = 10'h102 == r_count_13_io_out ? io_r_258_b : _GEN_10097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10099 = 10'h103 == r_count_13_io_out ? io_r_259_b : _GEN_10098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10100 = 10'h104 == r_count_13_io_out ? io_r_260_b : _GEN_10099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10101 = 10'h105 == r_count_13_io_out ? io_r_261_b : _GEN_10100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10102 = 10'h106 == r_count_13_io_out ? io_r_262_b : _GEN_10101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10103 = 10'h107 == r_count_13_io_out ? io_r_263_b : _GEN_10102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10104 = 10'h108 == r_count_13_io_out ? io_r_264_b : _GEN_10103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10105 = 10'h109 == r_count_13_io_out ? io_r_265_b : _GEN_10104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10106 = 10'h10a == r_count_13_io_out ? io_r_266_b : _GEN_10105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10107 = 10'h10b == r_count_13_io_out ? io_r_267_b : _GEN_10106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10108 = 10'h10c == r_count_13_io_out ? io_r_268_b : _GEN_10107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10109 = 10'h10d == r_count_13_io_out ? io_r_269_b : _GEN_10108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10110 = 10'h10e == r_count_13_io_out ? io_r_270_b : _GEN_10109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10111 = 10'h10f == r_count_13_io_out ? io_r_271_b : _GEN_10110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10112 = 10'h110 == r_count_13_io_out ? io_r_272_b : _GEN_10111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10113 = 10'h111 == r_count_13_io_out ? io_r_273_b : _GEN_10112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10114 = 10'h112 == r_count_13_io_out ? io_r_274_b : _GEN_10113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10115 = 10'h113 == r_count_13_io_out ? io_r_275_b : _GEN_10114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10116 = 10'h114 == r_count_13_io_out ? io_r_276_b : _GEN_10115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10117 = 10'h115 == r_count_13_io_out ? io_r_277_b : _GEN_10116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10118 = 10'h116 == r_count_13_io_out ? io_r_278_b : _GEN_10117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10119 = 10'h117 == r_count_13_io_out ? io_r_279_b : _GEN_10118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10120 = 10'h118 == r_count_13_io_out ? io_r_280_b : _GEN_10119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10121 = 10'h119 == r_count_13_io_out ? io_r_281_b : _GEN_10120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10122 = 10'h11a == r_count_13_io_out ? io_r_282_b : _GEN_10121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10123 = 10'h11b == r_count_13_io_out ? io_r_283_b : _GEN_10122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10124 = 10'h11c == r_count_13_io_out ? io_r_284_b : _GEN_10123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10125 = 10'h11d == r_count_13_io_out ? io_r_285_b : _GEN_10124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10126 = 10'h11e == r_count_13_io_out ? io_r_286_b : _GEN_10125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10127 = 10'h11f == r_count_13_io_out ? io_r_287_b : _GEN_10126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10128 = 10'h120 == r_count_13_io_out ? io_r_288_b : _GEN_10127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10129 = 10'h121 == r_count_13_io_out ? io_r_289_b : _GEN_10128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10130 = 10'h122 == r_count_13_io_out ? io_r_290_b : _GEN_10129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10131 = 10'h123 == r_count_13_io_out ? io_r_291_b : _GEN_10130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10132 = 10'h124 == r_count_13_io_out ? io_r_292_b : _GEN_10131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10133 = 10'h125 == r_count_13_io_out ? io_r_293_b : _GEN_10132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10134 = 10'h126 == r_count_13_io_out ? io_r_294_b : _GEN_10133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10135 = 10'h127 == r_count_13_io_out ? io_r_295_b : _GEN_10134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10136 = 10'h128 == r_count_13_io_out ? io_r_296_b : _GEN_10135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10137 = 10'h129 == r_count_13_io_out ? io_r_297_b : _GEN_10136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10138 = 10'h12a == r_count_13_io_out ? io_r_298_b : _GEN_10137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10139 = 10'h12b == r_count_13_io_out ? io_r_299_b : _GEN_10138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10140 = 10'h12c == r_count_13_io_out ? io_r_300_b : _GEN_10139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10141 = 10'h12d == r_count_13_io_out ? io_r_301_b : _GEN_10140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10142 = 10'h12e == r_count_13_io_out ? io_r_302_b : _GEN_10141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10143 = 10'h12f == r_count_13_io_out ? io_r_303_b : _GEN_10142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10144 = 10'h130 == r_count_13_io_out ? io_r_304_b : _GEN_10143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10145 = 10'h131 == r_count_13_io_out ? io_r_305_b : _GEN_10144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10146 = 10'h132 == r_count_13_io_out ? io_r_306_b : _GEN_10145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10147 = 10'h133 == r_count_13_io_out ? io_r_307_b : _GEN_10146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10148 = 10'h134 == r_count_13_io_out ? io_r_308_b : _GEN_10147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10149 = 10'h135 == r_count_13_io_out ? io_r_309_b : _GEN_10148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10150 = 10'h136 == r_count_13_io_out ? io_r_310_b : _GEN_10149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10151 = 10'h137 == r_count_13_io_out ? io_r_311_b : _GEN_10150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10152 = 10'h138 == r_count_13_io_out ? io_r_312_b : _GEN_10151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10153 = 10'h139 == r_count_13_io_out ? io_r_313_b : _GEN_10152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10154 = 10'h13a == r_count_13_io_out ? io_r_314_b : _GEN_10153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10155 = 10'h13b == r_count_13_io_out ? io_r_315_b : _GEN_10154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10156 = 10'h13c == r_count_13_io_out ? io_r_316_b : _GEN_10155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10157 = 10'h13d == r_count_13_io_out ? io_r_317_b : _GEN_10156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10158 = 10'h13e == r_count_13_io_out ? io_r_318_b : _GEN_10157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10159 = 10'h13f == r_count_13_io_out ? io_r_319_b : _GEN_10158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10160 = 10'h140 == r_count_13_io_out ? io_r_320_b : _GEN_10159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10161 = 10'h141 == r_count_13_io_out ? io_r_321_b : _GEN_10160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10162 = 10'h142 == r_count_13_io_out ? io_r_322_b : _GEN_10161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10163 = 10'h143 == r_count_13_io_out ? io_r_323_b : _GEN_10162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10164 = 10'h144 == r_count_13_io_out ? io_r_324_b : _GEN_10163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10165 = 10'h145 == r_count_13_io_out ? io_r_325_b : _GEN_10164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10166 = 10'h146 == r_count_13_io_out ? io_r_326_b : _GEN_10165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10167 = 10'h147 == r_count_13_io_out ? io_r_327_b : _GEN_10166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10168 = 10'h148 == r_count_13_io_out ? io_r_328_b : _GEN_10167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10169 = 10'h149 == r_count_13_io_out ? io_r_329_b : _GEN_10168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10170 = 10'h14a == r_count_13_io_out ? io_r_330_b : _GEN_10169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10171 = 10'h14b == r_count_13_io_out ? io_r_331_b : _GEN_10170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10172 = 10'h14c == r_count_13_io_out ? io_r_332_b : _GEN_10171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10173 = 10'h14d == r_count_13_io_out ? io_r_333_b : _GEN_10172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10174 = 10'h14e == r_count_13_io_out ? io_r_334_b : _GEN_10173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10175 = 10'h14f == r_count_13_io_out ? io_r_335_b : _GEN_10174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10176 = 10'h150 == r_count_13_io_out ? io_r_336_b : _GEN_10175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10177 = 10'h151 == r_count_13_io_out ? io_r_337_b : _GEN_10176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10178 = 10'h152 == r_count_13_io_out ? io_r_338_b : _GEN_10177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10179 = 10'h153 == r_count_13_io_out ? io_r_339_b : _GEN_10178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10180 = 10'h154 == r_count_13_io_out ? io_r_340_b : _GEN_10179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10181 = 10'h155 == r_count_13_io_out ? io_r_341_b : _GEN_10180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10182 = 10'h156 == r_count_13_io_out ? io_r_342_b : _GEN_10181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10183 = 10'h157 == r_count_13_io_out ? io_r_343_b : _GEN_10182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10184 = 10'h158 == r_count_13_io_out ? io_r_344_b : _GEN_10183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10185 = 10'h159 == r_count_13_io_out ? io_r_345_b : _GEN_10184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10186 = 10'h15a == r_count_13_io_out ? io_r_346_b : _GEN_10185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10187 = 10'h15b == r_count_13_io_out ? io_r_347_b : _GEN_10186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10188 = 10'h15c == r_count_13_io_out ? io_r_348_b : _GEN_10187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10189 = 10'h15d == r_count_13_io_out ? io_r_349_b : _GEN_10188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10190 = 10'h15e == r_count_13_io_out ? io_r_350_b : _GEN_10189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10191 = 10'h15f == r_count_13_io_out ? io_r_351_b : _GEN_10190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10192 = 10'h160 == r_count_13_io_out ? io_r_352_b : _GEN_10191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10193 = 10'h161 == r_count_13_io_out ? io_r_353_b : _GEN_10192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10194 = 10'h162 == r_count_13_io_out ? io_r_354_b : _GEN_10193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10195 = 10'h163 == r_count_13_io_out ? io_r_355_b : _GEN_10194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10196 = 10'h164 == r_count_13_io_out ? io_r_356_b : _GEN_10195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10197 = 10'h165 == r_count_13_io_out ? io_r_357_b : _GEN_10196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10198 = 10'h166 == r_count_13_io_out ? io_r_358_b : _GEN_10197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10199 = 10'h167 == r_count_13_io_out ? io_r_359_b : _GEN_10198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10200 = 10'h168 == r_count_13_io_out ? io_r_360_b : _GEN_10199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10201 = 10'h169 == r_count_13_io_out ? io_r_361_b : _GEN_10200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10202 = 10'h16a == r_count_13_io_out ? io_r_362_b : _GEN_10201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10203 = 10'h16b == r_count_13_io_out ? io_r_363_b : _GEN_10202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10204 = 10'h16c == r_count_13_io_out ? io_r_364_b : _GEN_10203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10205 = 10'h16d == r_count_13_io_out ? io_r_365_b : _GEN_10204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10206 = 10'h16e == r_count_13_io_out ? io_r_366_b : _GEN_10205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10207 = 10'h16f == r_count_13_io_out ? io_r_367_b : _GEN_10206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10208 = 10'h170 == r_count_13_io_out ? io_r_368_b : _GEN_10207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10209 = 10'h171 == r_count_13_io_out ? io_r_369_b : _GEN_10208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10210 = 10'h172 == r_count_13_io_out ? io_r_370_b : _GEN_10209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10211 = 10'h173 == r_count_13_io_out ? io_r_371_b : _GEN_10210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10212 = 10'h174 == r_count_13_io_out ? io_r_372_b : _GEN_10211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10213 = 10'h175 == r_count_13_io_out ? io_r_373_b : _GEN_10212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10214 = 10'h176 == r_count_13_io_out ? io_r_374_b : _GEN_10213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10215 = 10'h177 == r_count_13_io_out ? io_r_375_b : _GEN_10214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10216 = 10'h178 == r_count_13_io_out ? io_r_376_b : _GEN_10215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10217 = 10'h179 == r_count_13_io_out ? io_r_377_b : _GEN_10216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10218 = 10'h17a == r_count_13_io_out ? io_r_378_b : _GEN_10217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10219 = 10'h17b == r_count_13_io_out ? io_r_379_b : _GEN_10218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10220 = 10'h17c == r_count_13_io_out ? io_r_380_b : _GEN_10219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10221 = 10'h17d == r_count_13_io_out ? io_r_381_b : _GEN_10220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10222 = 10'h17e == r_count_13_io_out ? io_r_382_b : _GEN_10221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10223 = 10'h17f == r_count_13_io_out ? io_r_383_b : _GEN_10222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10224 = 10'h180 == r_count_13_io_out ? io_r_384_b : _GEN_10223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10225 = 10'h181 == r_count_13_io_out ? io_r_385_b : _GEN_10224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10226 = 10'h182 == r_count_13_io_out ? io_r_386_b : _GEN_10225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10227 = 10'h183 == r_count_13_io_out ? io_r_387_b : _GEN_10226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10228 = 10'h184 == r_count_13_io_out ? io_r_388_b : _GEN_10227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10229 = 10'h185 == r_count_13_io_out ? io_r_389_b : _GEN_10228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10230 = 10'h186 == r_count_13_io_out ? io_r_390_b : _GEN_10229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10231 = 10'h187 == r_count_13_io_out ? io_r_391_b : _GEN_10230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10232 = 10'h188 == r_count_13_io_out ? io_r_392_b : _GEN_10231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10233 = 10'h189 == r_count_13_io_out ? io_r_393_b : _GEN_10232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10234 = 10'h18a == r_count_13_io_out ? io_r_394_b : _GEN_10233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10235 = 10'h18b == r_count_13_io_out ? io_r_395_b : _GEN_10234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10236 = 10'h18c == r_count_13_io_out ? io_r_396_b : _GEN_10235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10237 = 10'h18d == r_count_13_io_out ? io_r_397_b : _GEN_10236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10238 = 10'h18e == r_count_13_io_out ? io_r_398_b : _GEN_10237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10239 = 10'h18f == r_count_13_io_out ? io_r_399_b : _GEN_10238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10240 = 10'h190 == r_count_13_io_out ? io_r_400_b : _GEN_10239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10241 = 10'h191 == r_count_13_io_out ? io_r_401_b : _GEN_10240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10242 = 10'h192 == r_count_13_io_out ? io_r_402_b : _GEN_10241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10243 = 10'h193 == r_count_13_io_out ? io_r_403_b : _GEN_10242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10244 = 10'h194 == r_count_13_io_out ? io_r_404_b : _GEN_10243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10245 = 10'h195 == r_count_13_io_out ? io_r_405_b : _GEN_10244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10246 = 10'h196 == r_count_13_io_out ? io_r_406_b : _GEN_10245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10247 = 10'h197 == r_count_13_io_out ? io_r_407_b : _GEN_10246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10248 = 10'h198 == r_count_13_io_out ? io_r_408_b : _GEN_10247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10249 = 10'h199 == r_count_13_io_out ? io_r_409_b : _GEN_10248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10250 = 10'h19a == r_count_13_io_out ? io_r_410_b : _GEN_10249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10251 = 10'h19b == r_count_13_io_out ? io_r_411_b : _GEN_10250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10252 = 10'h19c == r_count_13_io_out ? io_r_412_b : _GEN_10251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10253 = 10'h19d == r_count_13_io_out ? io_r_413_b : _GEN_10252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10254 = 10'h19e == r_count_13_io_out ? io_r_414_b : _GEN_10253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10255 = 10'h19f == r_count_13_io_out ? io_r_415_b : _GEN_10254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10256 = 10'h1a0 == r_count_13_io_out ? io_r_416_b : _GEN_10255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10257 = 10'h1a1 == r_count_13_io_out ? io_r_417_b : _GEN_10256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10258 = 10'h1a2 == r_count_13_io_out ? io_r_418_b : _GEN_10257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10259 = 10'h1a3 == r_count_13_io_out ? io_r_419_b : _GEN_10258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10260 = 10'h1a4 == r_count_13_io_out ? io_r_420_b : _GEN_10259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10261 = 10'h1a5 == r_count_13_io_out ? io_r_421_b : _GEN_10260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10262 = 10'h1a6 == r_count_13_io_out ? io_r_422_b : _GEN_10261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10263 = 10'h1a7 == r_count_13_io_out ? io_r_423_b : _GEN_10262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10264 = 10'h1a8 == r_count_13_io_out ? io_r_424_b : _GEN_10263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10265 = 10'h1a9 == r_count_13_io_out ? io_r_425_b : _GEN_10264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10266 = 10'h1aa == r_count_13_io_out ? io_r_426_b : _GEN_10265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10267 = 10'h1ab == r_count_13_io_out ? io_r_427_b : _GEN_10266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10268 = 10'h1ac == r_count_13_io_out ? io_r_428_b : _GEN_10267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10269 = 10'h1ad == r_count_13_io_out ? io_r_429_b : _GEN_10268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10270 = 10'h1ae == r_count_13_io_out ? io_r_430_b : _GEN_10269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10271 = 10'h1af == r_count_13_io_out ? io_r_431_b : _GEN_10270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10272 = 10'h1b0 == r_count_13_io_out ? io_r_432_b : _GEN_10271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10273 = 10'h1b1 == r_count_13_io_out ? io_r_433_b : _GEN_10272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10274 = 10'h1b2 == r_count_13_io_out ? io_r_434_b : _GEN_10273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10275 = 10'h1b3 == r_count_13_io_out ? io_r_435_b : _GEN_10274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10276 = 10'h1b4 == r_count_13_io_out ? io_r_436_b : _GEN_10275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10277 = 10'h1b5 == r_count_13_io_out ? io_r_437_b : _GEN_10276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10278 = 10'h1b6 == r_count_13_io_out ? io_r_438_b : _GEN_10277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10279 = 10'h1b7 == r_count_13_io_out ? io_r_439_b : _GEN_10278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10280 = 10'h1b8 == r_count_13_io_out ? io_r_440_b : _GEN_10279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10281 = 10'h1b9 == r_count_13_io_out ? io_r_441_b : _GEN_10280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10282 = 10'h1ba == r_count_13_io_out ? io_r_442_b : _GEN_10281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10283 = 10'h1bb == r_count_13_io_out ? io_r_443_b : _GEN_10282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10284 = 10'h1bc == r_count_13_io_out ? io_r_444_b : _GEN_10283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10285 = 10'h1bd == r_count_13_io_out ? io_r_445_b : _GEN_10284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10286 = 10'h1be == r_count_13_io_out ? io_r_446_b : _GEN_10285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10287 = 10'h1bf == r_count_13_io_out ? io_r_447_b : _GEN_10286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10288 = 10'h1c0 == r_count_13_io_out ? io_r_448_b : _GEN_10287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10289 = 10'h1c1 == r_count_13_io_out ? io_r_449_b : _GEN_10288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10290 = 10'h1c2 == r_count_13_io_out ? io_r_450_b : _GEN_10289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10291 = 10'h1c3 == r_count_13_io_out ? io_r_451_b : _GEN_10290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10292 = 10'h1c4 == r_count_13_io_out ? io_r_452_b : _GEN_10291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10293 = 10'h1c5 == r_count_13_io_out ? io_r_453_b : _GEN_10292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10294 = 10'h1c6 == r_count_13_io_out ? io_r_454_b : _GEN_10293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10295 = 10'h1c7 == r_count_13_io_out ? io_r_455_b : _GEN_10294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10296 = 10'h1c8 == r_count_13_io_out ? io_r_456_b : _GEN_10295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10297 = 10'h1c9 == r_count_13_io_out ? io_r_457_b : _GEN_10296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10298 = 10'h1ca == r_count_13_io_out ? io_r_458_b : _GEN_10297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10299 = 10'h1cb == r_count_13_io_out ? io_r_459_b : _GEN_10298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10300 = 10'h1cc == r_count_13_io_out ? io_r_460_b : _GEN_10299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10301 = 10'h1cd == r_count_13_io_out ? io_r_461_b : _GEN_10300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10302 = 10'h1ce == r_count_13_io_out ? io_r_462_b : _GEN_10301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10303 = 10'h1cf == r_count_13_io_out ? io_r_463_b : _GEN_10302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10304 = 10'h1d0 == r_count_13_io_out ? io_r_464_b : _GEN_10303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10305 = 10'h1d1 == r_count_13_io_out ? io_r_465_b : _GEN_10304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10306 = 10'h1d2 == r_count_13_io_out ? io_r_466_b : _GEN_10305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10307 = 10'h1d3 == r_count_13_io_out ? io_r_467_b : _GEN_10306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10308 = 10'h1d4 == r_count_13_io_out ? io_r_468_b : _GEN_10307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10309 = 10'h1d5 == r_count_13_io_out ? io_r_469_b : _GEN_10308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10310 = 10'h1d6 == r_count_13_io_out ? io_r_470_b : _GEN_10309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10311 = 10'h1d7 == r_count_13_io_out ? io_r_471_b : _GEN_10310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10312 = 10'h1d8 == r_count_13_io_out ? io_r_472_b : _GEN_10311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10313 = 10'h1d9 == r_count_13_io_out ? io_r_473_b : _GEN_10312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10314 = 10'h1da == r_count_13_io_out ? io_r_474_b : _GEN_10313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10315 = 10'h1db == r_count_13_io_out ? io_r_475_b : _GEN_10314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10316 = 10'h1dc == r_count_13_io_out ? io_r_476_b : _GEN_10315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10317 = 10'h1dd == r_count_13_io_out ? io_r_477_b : _GEN_10316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10318 = 10'h1de == r_count_13_io_out ? io_r_478_b : _GEN_10317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10319 = 10'h1df == r_count_13_io_out ? io_r_479_b : _GEN_10318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10320 = 10'h1e0 == r_count_13_io_out ? io_r_480_b : _GEN_10319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10321 = 10'h1e1 == r_count_13_io_out ? io_r_481_b : _GEN_10320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10322 = 10'h1e2 == r_count_13_io_out ? io_r_482_b : _GEN_10321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10323 = 10'h1e3 == r_count_13_io_out ? io_r_483_b : _GEN_10322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10324 = 10'h1e4 == r_count_13_io_out ? io_r_484_b : _GEN_10323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10325 = 10'h1e5 == r_count_13_io_out ? io_r_485_b : _GEN_10324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10326 = 10'h1e6 == r_count_13_io_out ? io_r_486_b : _GEN_10325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10327 = 10'h1e7 == r_count_13_io_out ? io_r_487_b : _GEN_10326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10328 = 10'h1e8 == r_count_13_io_out ? io_r_488_b : _GEN_10327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10329 = 10'h1e9 == r_count_13_io_out ? io_r_489_b : _GEN_10328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10330 = 10'h1ea == r_count_13_io_out ? io_r_490_b : _GEN_10329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10331 = 10'h1eb == r_count_13_io_out ? io_r_491_b : _GEN_10330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10332 = 10'h1ec == r_count_13_io_out ? io_r_492_b : _GEN_10331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10333 = 10'h1ed == r_count_13_io_out ? io_r_493_b : _GEN_10332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10334 = 10'h1ee == r_count_13_io_out ? io_r_494_b : _GEN_10333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10335 = 10'h1ef == r_count_13_io_out ? io_r_495_b : _GEN_10334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10336 = 10'h1f0 == r_count_13_io_out ? io_r_496_b : _GEN_10335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10337 = 10'h1f1 == r_count_13_io_out ? io_r_497_b : _GEN_10336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10338 = 10'h1f2 == r_count_13_io_out ? io_r_498_b : _GEN_10337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10339 = 10'h1f3 == r_count_13_io_out ? io_r_499_b : _GEN_10338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10340 = 10'h1f4 == r_count_13_io_out ? io_r_500_b : _GEN_10339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10341 = 10'h1f5 == r_count_13_io_out ? io_r_501_b : _GEN_10340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10342 = 10'h1f6 == r_count_13_io_out ? io_r_502_b : _GEN_10341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10343 = 10'h1f7 == r_count_13_io_out ? io_r_503_b : _GEN_10342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10344 = 10'h1f8 == r_count_13_io_out ? io_r_504_b : _GEN_10343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10345 = 10'h1f9 == r_count_13_io_out ? io_r_505_b : _GEN_10344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10346 = 10'h1fa == r_count_13_io_out ? io_r_506_b : _GEN_10345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10347 = 10'h1fb == r_count_13_io_out ? io_r_507_b : _GEN_10346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10348 = 10'h1fc == r_count_13_io_out ? io_r_508_b : _GEN_10347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10349 = 10'h1fd == r_count_13_io_out ? io_r_509_b : _GEN_10348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10350 = 10'h1fe == r_count_13_io_out ? io_r_510_b : _GEN_10349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10351 = 10'h1ff == r_count_13_io_out ? io_r_511_b : _GEN_10350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10352 = 10'h200 == r_count_13_io_out ? io_r_512_b : _GEN_10351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10353 = 10'h201 == r_count_13_io_out ? io_r_513_b : _GEN_10352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10354 = 10'h202 == r_count_13_io_out ? io_r_514_b : _GEN_10353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10355 = 10'h203 == r_count_13_io_out ? io_r_515_b : _GEN_10354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10356 = 10'h204 == r_count_13_io_out ? io_r_516_b : _GEN_10355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10357 = 10'h205 == r_count_13_io_out ? io_r_517_b : _GEN_10356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10358 = 10'h206 == r_count_13_io_out ? io_r_518_b : _GEN_10357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10359 = 10'h207 == r_count_13_io_out ? io_r_519_b : _GEN_10358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10360 = 10'h208 == r_count_13_io_out ? io_r_520_b : _GEN_10359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10361 = 10'h209 == r_count_13_io_out ? io_r_521_b : _GEN_10360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10362 = 10'h20a == r_count_13_io_out ? io_r_522_b : _GEN_10361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10363 = 10'h20b == r_count_13_io_out ? io_r_523_b : _GEN_10362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10364 = 10'h20c == r_count_13_io_out ? io_r_524_b : _GEN_10363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10365 = 10'h20d == r_count_13_io_out ? io_r_525_b : _GEN_10364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10366 = 10'h20e == r_count_13_io_out ? io_r_526_b : _GEN_10365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10367 = 10'h20f == r_count_13_io_out ? io_r_527_b : _GEN_10366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10368 = 10'h210 == r_count_13_io_out ? io_r_528_b : _GEN_10367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10369 = 10'h211 == r_count_13_io_out ? io_r_529_b : _GEN_10368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10370 = 10'h212 == r_count_13_io_out ? io_r_530_b : _GEN_10369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10371 = 10'h213 == r_count_13_io_out ? io_r_531_b : _GEN_10370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10372 = 10'h214 == r_count_13_io_out ? io_r_532_b : _GEN_10371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10373 = 10'h215 == r_count_13_io_out ? io_r_533_b : _GEN_10372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10374 = 10'h216 == r_count_13_io_out ? io_r_534_b : _GEN_10373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10375 = 10'h217 == r_count_13_io_out ? io_r_535_b : _GEN_10374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10376 = 10'h218 == r_count_13_io_out ? io_r_536_b : _GEN_10375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10377 = 10'h219 == r_count_13_io_out ? io_r_537_b : _GEN_10376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10378 = 10'h21a == r_count_13_io_out ? io_r_538_b : _GEN_10377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10379 = 10'h21b == r_count_13_io_out ? io_r_539_b : _GEN_10378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10380 = 10'h21c == r_count_13_io_out ? io_r_540_b : _GEN_10379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10381 = 10'h21d == r_count_13_io_out ? io_r_541_b : _GEN_10380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10382 = 10'h21e == r_count_13_io_out ? io_r_542_b : _GEN_10381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10383 = 10'h21f == r_count_13_io_out ? io_r_543_b : _GEN_10382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10384 = 10'h220 == r_count_13_io_out ? io_r_544_b : _GEN_10383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10385 = 10'h221 == r_count_13_io_out ? io_r_545_b : _GEN_10384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10386 = 10'h222 == r_count_13_io_out ? io_r_546_b : _GEN_10385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10387 = 10'h223 == r_count_13_io_out ? io_r_547_b : _GEN_10386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10388 = 10'h224 == r_count_13_io_out ? io_r_548_b : _GEN_10387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10389 = 10'h225 == r_count_13_io_out ? io_r_549_b : _GEN_10388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10390 = 10'h226 == r_count_13_io_out ? io_r_550_b : _GEN_10389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10391 = 10'h227 == r_count_13_io_out ? io_r_551_b : _GEN_10390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10392 = 10'h228 == r_count_13_io_out ? io_r_552_b : _GEN_10391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10393 = 10'h229 == r_count_13_io_out ? io_r_553_b : _GEN_10392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10394 = 10'h22a == r_count_13_io_out ? io_r_554_b : _GEN_10393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10395 = 10'h22b == r_count_13_io_out ? io_r_555_b : _GEN_10394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10396 = 10'h22c == r_count_13_io_out ? io_r_556_b : _GEN_10395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10397 = 10'h22d == r_count_13_io_out ? io_r_557_b : _GEN_10396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10398 = 10'h22e == r_count_13_io_out ? io_r_558_b : _GEN_10397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10399 = 10'h22f == r_count_13_io_out ? io_r_559_b : _GEN_10398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10400 = 10'h230 == r_count_13_io_out ? io_r_560_b : _GEN_10399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10401 = 10'h231 == r_count_13_io_out ? io_r_561_b : _GEN_10400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10402 = 10'h232 == r_count_13_io_out ? io_r_562_b : _GEN_10401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10403 = 10'h233 == r_count_13_io_out ? io_r_563_b : _GEN_10402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10404 = 10'h234 == r_count_13_io_out ? io_r_564_b : _GEN_10403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10405 = 10'h235 == r_count_13_io_out ? io_r_565_b : _GEN_10404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10406 = 10'h236 == r_count_13_io_out ? io_r_566_b : _GEN_10405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10407 = 10'h237 == r_count_13_io_out ? io_r_567_b : _GEN_10406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10408 = 10'h238 == r_count_13_io_out ? io_r_568_b : _GEN_10407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10409 = 10'h239 == r_count_13_io_out ? io_r_569_b : _GEN_10408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10410 = 10'h23a == r_count_13_io_out ? io_r_570_b : _GEN_10409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10411 = 10'h23b == r_count_13_io_out ? io_r_571_b : _GEN_10410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10412 = 10'h23c == r_count_13_io_out ? io_r_572_b : _GEN_10411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10413 = 10'h23d == r_count_13_io_out ? io_r_573_b : _GEN_10412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10414 = 10'h23e == r_count_13_io_out ? io_r_574_b : _GEN_10413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10415 = 10'h23f == r_count_13_io_out ? io_r_575_b : _GEN_10414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10416 = 10'h240 == r_count_13_io_out ? io_r_576_b : _GEN_10415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10417 = 10'h241 == r_count_13_io_out ? io_r_577_b : _GEN_10416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10418 = 10'h242 == r_count_13_io_out ? io_r_578_b : _GEN_10417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10419 = 10'h243 == r_count_13_io_out ? io_r_579_b : _GEN_10418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10420 = 10'h244 == r_count_13_io_out ? io_r_580_b : _GEN_10419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10421 = 10'h245 == r_count_13_io_out ? io_r_581_b : _GEN_10420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10422 = 10'h246 == r_count_13_io_out ? io_r_582_b : _GEN_10421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10423 = 10'h247 == r_count_13_io_out ? io_r_583_b : _GEN_10422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10424 = 10'h248 == r_count_13_io_out ? io_r_584_b : _GEN_10423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10425 = 10'h249 == r_count_13_io_out ? io_r_585_b : _GEN_10424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10426 = 10'h24a == r_count_13_io_out ? io_r_586_b : _GEN_10425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10427 = 10'h24b == r_count_13_io_out ? io_r_587_b : _GEN_10426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10428 = 10'h24c == r_count_13_io_out ? io_r_588_b : _GEN_10427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10429 = 10'h24d == r_count_13_io_out ? io_r_589_b : _GEN_10428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10430 = 10'h24e == r_count_13_io_out ? io_r_590_b : _GEN_10429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10431 = 10'h24f == r_count_13_io_out ? io_r_591_b : _GEN_10430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10432 = 10'h250 == r_count_13_io_out ? io_r_592_b : _GEN_10431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10433 = 10'h251 == r_count_13_io_out ? io_r_593_b : _GEN_10432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10434 = 10'h252 == r_count_13_io_out ? io_r_594_b : _GEN_10433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10435 = 10'h253 == r_count_13_io_out ? io_r_595_b : _GEN_10434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10436 = 10'h254 == r_count_13_io_out ? io_r_596_b : _GEN_10435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10437 = 10'h255 == r_count_13_io_out ? io_r_597_b : _GEN_10436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10438 = 10'h256 == r_count_13_io_out ? io_r_598_b : _GEN_10437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10439 = 10'h257 == r_count_13_io_out ? io_r_599_b : _GEN_10438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10440 = 10'h258 == r_count_13_io_out ? io_r_600_b : _GEN_10439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10441 = 10'h259 == r_count_13_io_out ? io_r_601_b : _GEN_10440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10442 = 10'h25a == r_count_13_io_out ? io_r_602_b : _GEN_10441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10443 = 10'h25b == r_count_13_io_out ? io_r_603_b : _GEN_10442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10444 = 10'h25c == r_count_13_io_out ? io_r_604_b : _GEN_10443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10445 = 10'h25d == r_count_13_io_out ? io_r_605_b : _GEN_10444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10446 = 10'h25e == r_count_13_io_out ? io_r_606_b : _GEN_10445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10447 = 10'h25f == r_count_13_io_out ? io_r_607_b : _GEN_10446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10448 = 10'h260 == r_count_13_io_out ? io_r_608_b : _GEN_10447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10449 = 10'h261 == r_count_13_io_out ? io_r_609_b : _GEN_10448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10450 = 10'h262 == r_count_13_io_out ? io_r_610_b : _GEN_10449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10451 = 10'h263 == r_count_13_io_out ? io_r_611_b : _GEN_10450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10452 = 10'h264 == r_count_13_io_out ? io_r_612_b : _GEN_10451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10453 = 10'h265 == r_count_13_io_out ? io_r_613_b : _GEN_10452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10454 = 10'h266 == r_count_13_io_out ? io_r_614_b : _GEN_10453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10455 = 10'h267 == r_count_13_io_out ? io_r_615_b : _GEN_10454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10456 = 10'h268 == r_count_13_io_out ? io_r_616_b : _GEN_10455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10457 = 10'h269 == r_count_13_io_out ? io_r_617_b : _GEN_10456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10458 = 10'h26a == r_count_13_io_out ? io_r_618_b : _GEN_10457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10459 = 10'h26b == r_count_13_io_out ? io_r_619_b : _GEN_10458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10460 = 10'h26c == r_count_13_io_out ? io_r_620_b : _GEN_10459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10461 = 10'h26d == r_count_13_io_out ? io_r_621_b : _GEN_10460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10462 = 10'h26e == r_count_13_io_out ? io_r_622_b : _GEN_10461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10463 = 10'h26f == r_count_13_io_out ? io_r_623_b : _GEN_10462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10464 = 10'h270 == r_count_13_io_out ? io_r_624_b : _GEN_10463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10465 = 10'h271 == r_count_13_io_out ? io_r_625_b : _GEN_10464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10466 = 10'h272 == r_count_13_io_out ? io_r_626_b : _GEN_10465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10467 = 10'h273 == r_count_13_io_out ? io_r_627_b : _GEN_10466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10468 = 10'h274 == r_count_13_io_out ? io_r_628_b : _GEN_10467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10469 = 10'h275 == r_count_13_io_out ? io_r_629_b : _GEN_10468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10470 = 10'h276 == r_count_13_io_out ? io_r_630_b : _GEN_10469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10471 = 10'h277 == r_count_13_io_out ? io_r_631_b : _GEN_10470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10472 = 10'h278 == r_count_13_io_out ? io_r_632_b : _GEN_10471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10473 = 10'h279 == r_count_13_io_out ? io_r_633_b : _GEN_10472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10474 = 10'h27a == r_count_13_io_out ? io_r_634_b : _GEN_10473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10475 = 10'h27b == r_count_13_io_out ? io_r_635_b : _GEN_10474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10476 = 10'h27c == r_count_13_io_out ? io_r_636_b : _GEN_10475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10477 = 10'h27d == r_count_13_io_out ? io_r_637_b : _GEN_10476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10478 = 10'h27e == r_count_13_io_out ? io_r_638_b : _GEN_10477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10479 = 10'h27f == r_count_13_io_out ? io_r_639_b : _GEN_10478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10480 = 10'h280 == r_count_13_io_out ? io_r_640_b : _GEN_10479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10481 = 10'h281 == r_count_13_io_out ? io_r_641_b : _GEN_10480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10482 = 10'h282 == r_count_13_io_out ? io_r_642_b : _GEN_10481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10483 = 10'h283 == r_count_13_io_out ? io_r_643_b : _GEN_10482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10484 = 10'h284 == r_count_13_io_out ? io_r_644_b : _GEN_10483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10485 = 10'h285 == r_count_13_io_out ? io_r_645_b : _GEN_10484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10486 = 10'h286 == r_count_13_io_out ? io_r_646_b : _GEN_10485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10487 = 10'h287 == r_count_13_io_out ? io_r_647_b : _GEN_10486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10488 = 10'h288 == r_count_13_io_out ? io_r_648_b : _GEN_10487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10489 = 10'h289 == r_count_13_io_out ? io_r_649_b : _GEN_10488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10490 = 10'h28a == r_count_13_io_out ? io_r_650_b : _GEN_10489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10491 = 10'h28b == r_count_13_io_out ? io_r_651_b : _GEN_10490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10492 = 10'h28c == r_count_13_io_out ? io_r_652_b : _GEN_10491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10493 = 10'h28d == r_count_13_io_out ? io_r_653_b : _GEN_10492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10494 = 10'h28e == r_count_13_io_out ? io_r_654_b : _GEN_10493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10495 = 10'h28f == r_count_13_io_out ? io_r_655_b : _GEN_10494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10496 = 10'h290 == r_count_13_io_out ? io_r_656_b : _GEN_10495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10497 = 10'h291 == r_count_13_io_out ? io_r_657_b : _GEN_10496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10498 = 10'h292 == r_count_13_io_out ? io_r_658_b : _GEN_10497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10499 = 10'h293 == r_count_13_io_out ? io_r_659_b : _GEN_10498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10500 = 10'h294 == r_count_13_io_out ? io_r_660_b : _GEN_10499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10501 = 10'h295 == r_count_13_io_out ? io_r_661_b : _GEN_10500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10502 = 10'h296 == r_count_13_io_out ? io_r_662_b : _GEN_10501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10503 = 10'h297 == r_count_13_io_out ? io_r_663_b : _GEN_10502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10504 = 10'h298 == r_count_13_io_out ? io_r_664_b : _GEN_10503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10505 = 10'h299 == r_count_13_io_out ? io_r_665_b : _GEN_10504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10506 = 10'h29a == r_count_13_io_out ? io_r_666_b : _GEN_10505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10507 = 10'h29b == r_count_13_io_out ? io_r_667_b : _GEN_10506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10508 = 10'h29c == r_count_13_io_out ? io_r_668_b : _GEN_10507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10509 = 10'h29d == r_count_13_io_out ? io_r_669_b : _GEN_10508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10510 = 10'h29e == r_count_13_io_out ? io_r_670_b : _GEN_10509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10511 = 10'h29f == r_count_13_io_out ? io_r_671_b : _GEN_10510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10512 = 10'h2a0 == r_count_13_io_out ? io_r_672_b : _GEN_10511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10513 = 10'h2a1 == r_count_13_io_out ? io_r_673_b : _GEN_10512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10514 = 10'h2a2 == r_count_13_io_out ? io_r_674_b : _GEN_10513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10515 = 10'h2a3 == r_count_13_io_out ? io_r_675_b : _GEN_10514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10516 = 10'h2a4 == r_count_13_io_out ? io_r_676_b : _GEN_10515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10517 = 10'h2a5 == r_count_13_io_out ? io_r_677_b : _GEN_10516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10518 = 10'h2a6 == r_count_13_io_out ? io_r_678_b : _GEN_10517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10519 = 10'h2a7 == r_count_13_io_out ? io_r_679_b : _GEN_10518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10520 = 10'h2a8 == r_count_13_io_out ? io_r_680_b : _GEN_10519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10521 = 10'h2a9 == r_count_13_io_out ? io_r_681_b : _GEN_10520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10522 = 10'h2aa == r_count_13_io_out ? io_r_682_b : _GEN_10521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10523 = 10'h2ab == r_count_13_io_out ? io_r_683_b : _GEN_10522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10524 = 10'h2ac == r_count_13_io_out ? io_r_684_b : _GEN_10523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10525 = 10'h2ad == r_count_13_io_out ? io_r_685_b : _GEN_10524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10526 = 10'h2ae == r_count_13_io_out ? io_r_686_b : _GEN_10525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10527 = 10'h2af == r_count_13_io_out ? io_r_687_b : _GEN_10526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10528 = 10'h2b0 == r_count_13_io_out ? io_r_688_b : _GEN_10527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10529 = 10'h2b1 == r_count_13_io_out ? io_r_689_b : _GEN_10528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10530 = 10'h2b2 == r_count_13_io_out ? io_r_690_b : _GEN_10529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10531 = 10'h2b3 == r_count_13_io_out ? io_r_691_b : _GEN_10530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10532 = 10'h2b4 == r_count_13_io_out ? io_r_692_b : _GEN_10531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10533 = 10'h2b5 == r_count_13_io_out ? io_r_693_b : _GEN_10532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10534 = 10'h2b6 == r_count_13_io_out ? io_r_694_b : _GEN_10533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10535 = 10'h2b7 == r_count_13_io_out ? io_r_695_b : _GEN_10534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10536 = 10'h2b8 == r_count_13_io_out ? io_r_696_b : _GEN_10535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10537 = 10'h2b9 == r_count_13_io_out ? io_r_697_b : _GEN_10536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10538 = 10'h2ba == r_count_13_io_out ? io_r_698_b : _GEN_10537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10539 = 10'h2bb == r_count_13_io_out ? io_r_699_b : _GEN_10538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10540 = 10'h2bc == r_count_13_io_out ? io_r_700_b : _GEN_10539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10541 = 10'h2bd == r_count_13_io_out ? io_r_701_b : _GEN_10540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10542 = 10'h2be == r_count_13_io_out ? io_r_702_b : _GEN_10541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10543 = 10'h2bf == r_count_13_io_out ? io_r_703_b : _GEN_10542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10544 = 10'h2c0 == r_count_13_io_out ? io_r_704_b : _GEN_10543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10545 = 10'h2c1 == r_count_13_io_out ? io_r_705_b : _GEN_10544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10546 = 10'h2c2 == r_count_13_io_out ? io_r_706_b : _GEN_10545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10547 = 10'h2c3 == r_count_13_io_out ? io_r_707_b : _GEN_10546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10548 = 10'h2c4 == r_count_13_io_out ? io_r_708_b : _GEN_10547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10549 = 10'h2c5 == r_count_13_io_out ? io_r_709_b : _GEN_10548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10550 = 10'h2c6 == r_count_13_io_out ? io_r_710_b : _GEN_10549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10551 = 10'h2c7 == r_count_13_io_out ? io_r_711_b : _GEN_10550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10552 = 10'h2c8 == r_count_13_io_out ? io_r_712_b : _GEN_10551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10553 = 10'h2c9 == r_count_13_io_out ? io_r_713_b : _GEN_10552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10554 = 10'h2ca == r_count_13_io_out ? io_r_714_b : _GEN_10553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10555 = 10'h2cb == r_count_13_io_out ? io_r_715_b : _GEN_10554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10556 = 10'h2cc == r_count_13_io_out ? io_r_716_b : _GEN_10555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10557 = 10'h2cd == r_count_13_io_out ? io_r_717_b : _GEN_10556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10558 = 10'h2ce == r_count_13_io_out ? io_r_718_b : _GEN_10557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10559 = 10'h2cf == r_count_13_io_out ? io_r_719_b : _GEN_10558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10560 = 10'h2d0 == r_count_13_io_out ? io_r_720_b : _GEN_10559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10561 = 10'h2d1 == r_count_13_io_out ? io_r_721_b : _GEN_10560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10562 = 10'h2d2 == r_count_13_io_out ? io_r_722_b : _GEN_10561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10563 = 10'h2d3 == r_count_13_io_out ? io_r_723_b : _GEN_10562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10564 = 10'h2d4 == r_count_13_io_out ? io_r_724_b : _GEN_10563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10565 = 10'h2d5 == r_count_13_io_out ? io_r_725_b : _GEN_10564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10566 = 10'h2d6 == r_count_13_io_out ? io_r_726_b : _GEN_10565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10567 = 10'h2d7 == r_count_13_io_out ? io_r_727_b : _GEN_10566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10568 = 10'h2d8 == r_count_13_io_out ? io_r_728_b : _GEN_10567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10569 = 10'h2d9 == r_count_13_io_out ? io_r_729_b : _GEN_10568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10570 = 10'h2da == r_count_13_io_out ? io_r_730_b : _GEN_10569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10571 = 10'h2db == r_count_13_io_out ? io_r_731_b : _GEN_10570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10572 = 10'h2dc == r_count_13_io_out ? io_r_732_b : _GEN_10571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10573 = 10'h2dd == r_count_13_io_out ? io_r_733_b : _GEN_10572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10574 = 10'h2de == r_count_13_io_out ? io_r_734_b : _GEN_10573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10575 = 10'h2df == r_count_13_io_out ? io_r_735_b : _GEN_10574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10576 = 10'h2e0 == r_count_13_io_out ? io_r_736_b : _GEN_10575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10577 = 10'h2e1 == r_count_13_io_out ? io_r_737_b : _GEN_10576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10578 = 10'h2e2 == r_count_13_io_out ? io_r_738_b : _GEN_10577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10579 = 10'h2e3 == r_count_13_io_out ? io_r_739_b : _GEN_10578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10580 = 10'h2e4 == r_count_13_io_out ? io_r_740_b : _GEN_10579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10581 = 10'h2e5 == r_count_13_io_out ? io_r_741_b : _GEN_10580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10582 = 10'h2e6 == r_count_13_io_out ? io_r_742_b : _GEN_10581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10583 = 10'h2e7 == r_count_13_io_out ? io_r_743_b : _GEN_10582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10584 = 10'h2e8 == r_count_13_io_out ? io_r_744_b : _GEN_10583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10585 = 10'h2e9 == r_count_13_io_out ? io_r_745_b : _GEN_10584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10586 = 10'h2ea == r_count_13_io_out ? io_r_746_b : _GEN_10585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10587 = 10'h2eb == r_count_13_io_out ? io_r_747_b : _GEN_10586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10588 = 10'h2ec == r_count_13_io_out ? io_r_748_b : _GEN_10587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10591 = 10'h1 == r_count_14_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10592 = 10'h2 == r_count_14_io_out ? io_r_2_b : _GEN_10591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10593 = 10'h3 == r_count_14_io_out ? io_r_3_b : _GEN_10592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10594 = 10'h4 == r_count_14_io_out ? io_r_4_b : _GEN_10593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10595 = 10'h5 == r_count_14_io_out ? io_r_5_b : _GEN_10594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10596 = 10'h6 == r_count_14_io_out ? io_r_6_b : _GEN_10595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10597 = 10'h7 == r_count_14_io_out ? io_r_7_b : _GEN_10596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10598 = 10'h8 == r_count_14_io_out ? io_r_8_b : _GEN_10597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10599 = 10'h9 == r_count_14_io_out ? io_r_9_b : _GEN_10598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10600 = 10'ha == r_count_14_io_out ? io_r_10_b : _GEN_10599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10601 = 10'hb == r_count_14_io_out ? io_r_11_b : _GEN_10600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10602 = 10'hc == r_count_14_io_out ? io_r_12_b : _GEN_10601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10603 = 10'hd == r_count_14_io_out ? io_r_13_b : _GEN_10602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10604 = 10'he == r_count_14_io_out ? io_r_14_b : _GEN_10603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10605 = 10'hf == r_count_14_io_out ? io_r_15_b : _GEN_10604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10606 = 10'h10 == r_count_14_io_out ? io_r_16_b : _GEN_10605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10607 = 10'h11 == r_count_14_io_out ? io_r_17_b : _GEN_10606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10608 = 10'h12 == r_count_14_io_out ? io_r_18_b : _GEN_10607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10609 = 10'h13 == r_count_14_io_out ? io_r_19_b : _GEN_10608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10610 = 10'h14 == r_count_14_io_out ? io_r_20_b : _GEN_10609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10611 = 10'h15 == r_count_14_io_out ? io_r_21_b : _GEN_10610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10612 = 10'h16 == r_count_14_io_out ? io_r_22_b : _GEN_10611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10613 = 10'h17 == r_count_14_io_out ? io_r_23_b : _GEN_10612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10614 = 10'h18 == r_count_14_io_out ? io_r_24_b : _GEN_10613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10615 = 10'h19 == r_count_14_io_out ? io_r_25_b : _GEN_10614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10616 = 10'h1a == r_count_14_io_out ? io_r_26_b : _GEN_10615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10617 = 10'h1b == r_count_14_io_out ? io_r_27_b : _GEN_10616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10618 = 10'h1c == r_count_14_io_out ? io_r_28_b : _GEN_10617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10619 = 10'h1d == r_count_14_io_out ? io_r_29_b : _GEN_10618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10620 = 10'h1e == r_count_14_io_out ? io_r_30_b : _GEN_10619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10621 = 10'h1f == r_count_14_io_out ? io_r_31_b : _GEN_10620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10622 = 10'h20 == r_count_14_io_out ? io_r_32_b : _GEN_10621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10623 = 10'h21 == r_count_14_io_out ? io_r_33_b : _GEN_10622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10624 = 10'h22 == r_count_14_io_out ? io_r_34_b : _GEN_10623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10625 = 10'h23 == r_count_14_io_out ? io_r_35_b : _GEN_10624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10626 = 10'h24 == r_count_14_io_out ? io_r_36_b : _GEN_10625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10627 = 10'h25 == r_count_14_io_out ? io_r_37_b : _GEN_10626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10628 = 10'h26 == r_count_14_io_out ? io_r_38_b : _GEN_10627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10629 = 10'h27 == r_count_14_io_out ? io_r_39_b : _GEN_10628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10630 = 10'h28 == r_count_14_io_out ? io_r_40_b : _GEN_10629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10631 = 10'h29 == r_count_14_io_out ? io_r_41_b : _GEN_10630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10632 = 10'h2a == r_count_14_io_out ? io_r_42_b : _GEN_10631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10633 = 10'h2b == r_count_14_io_out ? io_r_43_b : _GEN_10632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10634 = 10'h2c == r_count_14_io_out ? io_r_44_b : _GEN_10633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10635 = 10'h2d == r_count_14_io_out ? io_r_45_b : _GEN_10634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10636 = 10'h2e == r_count_14_io_out ? io_r_46_b : _GEN_10635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10637 = 10'h2f == r_count_14_io_out ? io_r_47_b : _GEN_10636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10638 = 10'h30 == r_count_14_io_out ? io_r_48_b : _GEN_10637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10639 = 10'h31 == r_count_14_io_out ? io_r_49_b : _GEN_10638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10640 = 10'h32 == r_count_14_io_out ? io_r_50_b : _GEN_10639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10641 = 10'h33 == r_count_14_io_out ? io_r_51_b : _GEN_10640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10642 = 10'h34 == r_count_14_io_out ? io_r_52_b : _GEN_10641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10643 = 10'h35 == r_count_14_io_out ? io_r_53_b : _GEN_10642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10644 = 10'h36 == r_count_14_io_out ? io_r_54_b : _GEN_10643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10645 = 10'h37 == r_count_14_io_out ? io_r_55_b : _GEN_10644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10646 = 10'h38 == r_count_14_io_out ? io_r_56_b : _GEN_10645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10647 = 10'h39 == r_count_14_io_out ? io_r_57_b : _GEN_10646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10648 = 10'h3a == r_count_14_io_out ? io_r_58_b : _GEN_10647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10649 = 10'h3b == r_count_14_io_out ? io_r_59_b : _GEN_10648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10650 = 10'h3c == r_count_14_io_out ? io_r_60_b : _GEN_10649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10651 = 10'h3d == r_count_14_io_out ? io_r_61_b : _GEN_10650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10652 = 10'h3e == r_count_14_io_out ? io_r_62_b : _GEN_10651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10653 = 10'h3f == r_count_14_io_out ? io_r_63_b : _GEN_10652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10654 = 10'h40 == r_count_14_io_out ? io_r_64_b : _GEN_10653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10655 = 10'h41 == r_count_14_io_out ? io_r_65_b : _GEN_10654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10656 = 10'h42 == r_count_14_io_out ? io_r_66_b : _GEN_10655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10657 = 10'h43 == r_count_14_io_out ? io_r_67_b : _GEN_10656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10658 = 10'h44 == r_count_14_io_out ? io_r_68_b : _GEN_10657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10659 = 10'h45 == r_count_14_io_out ? io_r_69_b : _GEN_10658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10660 = 10'h46 == r_count_14_io_out ? io_r_70_b : _GEN_10659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10661 = 10'h47 == r_count_14_io_out ? io_r_71_b : _GEN_10660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10662 = 10'h48 == r_count_14_io_out ? io_r_72_b : _GEN_10661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10663 = 10'h49 == r_count_14_io_out ? io_r_73_b : _GEN_10662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10664 = 10'h4a == r_count_14_io_out ? io_r_74_b : _GEN_10663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10665 = 10'h4b == r_count_14_io_out ? io_r_75_b : _GEN_10664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10666 = 10'h4c == r_count_14_io_out ? io_r_76_b : _GEN_10665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10667 = 10'h4d == r_count_14_io_out ? io_r_77_b : _GEN_10666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10668 = 10'h4e == r_count_14_io_out ? io_r_78_b : _GEN_10667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10669 = 10'h4f == r_count_14_io_out ? io_r_79_b : _GEN_10668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10670 = 10'h50 == r_count_14_io_out ? io_r_80_b : _GEN_10669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10671 = 10'h51 == r_count_14_io_out ? io_r_81_b : _GEN_10670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10672 = 10'h52 == r_count_14_io_out ? io_r_82_b : _GEN_10671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10673 = 10'h53 == r_count_14_io_out ? io_r_83_b : _GEN_10672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10674 = 10'h54 == r_count_14_io_out ? io_r_84_b : _GEN_10673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10675 = 10'h55 == r_count_14_io_out ? io_r_85_b : _GEN_10674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10676 = 10'h56 == r_count_14_io_out ? io_r_86_b : _GEN_10675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10677 = 10'h57 == r_count_14_io_out ? io_r_87_b : _GEN_10676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10678 = 10'h58 == r_count_14_io_out ? io_r_88_b : _GEN_10677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10679 = 10'h59 == r_count_14_io_out ? io_r_89_b : _GEN_10678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10680 = 10'h5a == r_count_14_io_out ? io_r_90_b : _GEN_10679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10681 = 10'h5b == r_count_14_io_out ? io_r_91_b : _GEN_10680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10682 = 10'h5c == r_count_14_io_out ? io_r_92_b : _GEN_10681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10683 = 10'h5d == r_count_14_io_out ? io_r_93_b : _GEN_10682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10684 = 10'h5e == r_count_14_io_out ? io_r_94_b : _GEN_10683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10685 = 10'h5f == r_count_14_io_out ? io_r_95_b : _GEN_10684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10686 = 10'h60 == r_count_14_io_out ? io_r_96_b : _GEN_10685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10687 = 10'h61 == r_count_14_io_out ? io_r_97_b : _GEN_10686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10688 = 10'h62 == r_count_14_io_out ? io_r_98_b : _GEN_10687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10689 = 10'h63 == r_count_14_io_out ? io_r_99_b : _GEN_10688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10690 = 10'h64 == r_count_14_io_out ? io_r_100_b : _GEN_10689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10691 = 10'h65 == r_count_14_io_out ? io_r_101_b : _GEN_10690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10692 = 10'h66 == r_count_14_io_out ? io_r_102_b : _GEN_10691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10693 = 10'h67 == r_count_14_io_out ? io_r_103_b : _GEN_10692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10694 = 10'h68 == r_count_14_io_out ? io_r_104_b : _GEN_10693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10695 = 10'h69 == r_count_14_io_out ? io_r_105_b : _GEN_10694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10696 = 10'h6a == r_count_14_io_out ? io_r_106_b : _GEN_10695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10697 = 10'h6b == r_count_14_io_out ? io_r_107_b : _GEN_10696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10698 = 10'h6c == r_count_14_io_out ? io_r_108_b : _GEN_10697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10699 = 10'h6d == r_count_14_io_out ? io_r_109_b : _GEN_10698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10700 = 10'h6e == r_count_14_io_out ? io_r_110_b : _GEN_10699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10701 = 10'h6f == r_count_14_io_out ? io_r_111_b : _GEN_10700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10702 = 10'h70 == r_count_14_io_out ? io_r_112_b : _GEN_10701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10703 = 10'h71 == r_count_14_io_out ? io_r_113_b : _GEN_10702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10704 = 10'h72 == r_count_14_io_out ? io_r_114_b : _GEN_10703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10705 = 10'h73 == r_count_14_io_out ? io_r_115_b : _GEN_10704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10706 = 10'h74 == r_count_14_io_out ? io_r_116_b : _GEN_10705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10707 = 10'h75 == r_count_14_io_out ? io_r_117_b : _GEN_10706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10708 = 10'h76 == r_count_14_io_out ? io_r_118_b : _GEN_10707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10709 = 10'h77 == r_count_14_io_out ? io_r_119_b : _GEN_10708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10710 = 10'h78 == r_count_14_io_out ? io_r_120_b : _GEN_10709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10711 = 10'h79 == r_count_14_io_out ? io_r_121_b : _GEN_10710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10712 = 10'h7a == r_count_14_io_out ? io_r_122_b : _GEN_10711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10713 = 10'h7b == r_count_14_io_out ? io_r_123_b : _GEN_10712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10714 = 10'h7c == r_count_14_io_out ? io_r_124_b : _GEN_10713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10715 = 10'h7d == r_count_14_io_out ? io_r_125_b : _GEN_10714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10716 = 10'h7e == r_count_14_io_out ? io_r_126_b : _GEN_10715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10717 = 10'h7f == r_count_14_io_out ? io_r_127_b : _GEN_10716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10718 = 10'h80 == r_count_14_io_out ? io_r_128_b : _GEN_10717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10719 = 10'h81 == r_count_14_io_out ? io_r_129_b : _GEN_10718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10720 = 10'h82 == r_count_14_io_out ? io_r_130_b : _GEN_10719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10721 = 10'h83 == r_count_14_io_out ? io_r_131_b : _GEN_10720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10722 = 10'h84 == r_count_14_io_out ? io_r_132_b : _GEN_10721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10723 = 10'h85 == r_count_14_io_out ? io_r_133_b : _GEN_10722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10724 = 10'h86 == r_count_14_io_out ? io_r_134_b : _GEN_10723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10725 = 10'h87 == r_count_14_io_out ? io_r_135_b : _GEN_10724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10726 = 10'h88 == r_count_14_io_out ? io_r_136_b : _GEN_10725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10727 = 10'h89 == r_count_14_io_out ? io_r_137_b : _GEN_10726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10728 = 10'h8a == r_count_14_io_out ? io_r_138_b : _GEN_10727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10729 = 10'h8b == r_count_14_io_out ? io_r_139_b : _GEN_10728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10730 = 10'h8c == r_count_14_io_out ? io_r_140_b : _GEN_10729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10731 = 10'h8d == r_count_14_io_out ? io_r_141_b : _GEN_10730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10732 = 10'h8e == r_count_14_io_out ? io_r_142_b : _GEN_10731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10733 = 10'h8f == r_count_14_io_out ? io_r_143_b : _GEN_10732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10734 = 10'h90 == r_count_14_io_out ? io_r_144_b : _GEN_10733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10735 = 10'h91 == r_count_14_io_out ? io_r_145_b : _GEN_10734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10736 = 10'h92 == r_count_14_io_out ? io_r_146_b : _GEN_10735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10737 = 10'h93 == r_count_14_io_out ? io_r_147_b : _GEN_10736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10738 = 10'h94 == r_count_14_io_out ? io_r_148_b : _GEN_10737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10739 = 10'h95 == r_count_14_io_out ? io_r_149_b : _GEN_10738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10740 = 10'h96 == r_count_14_io_out ? io_r_150_b : _GEN_10739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10741 = 10'h97 == r_count_14_io_out ? io_r_151_b : _GEN_10740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10742 = 10'h98 == r_count_14_io_out ? io_r_152_b : _GEN_10741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10743 = 10'h99 == r_count_14_io_out ? io_r_153_b : _GEN_10742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10744 = 10'h9a == r_count_14_io_out ? io_r_154_b : _GEN_10743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10745 = 10'h9b == r_count_14_io_out ? io_r_155_b : _GEN_10744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10746 = 10'h9c == r_count_14_io_out ? io_r_156_b : _GEN_10745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10747 = 10'h9d == r_count_14_io_out ? io_r_157_b : _GEN_10746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10748 = 10'h9e == r_count_14_io_out ? io_r_158_b : _GEN_10747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10749 = 10'h9f == r_count_14_io_out ? io_r_159_b : _GEN_10748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10750 = 10'ha0 == r_count_14_io_out ? io_r_160_b : _GEN_10749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10751 = 10'ha1 == r_count_14_io_out ? io_r_161_b : _GEN_10750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10752 = 10'ha2 == r_count_14_io_out ? io_r_162_b : _GEN_10751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10753 = 10'ha3 == r_count_14_io_out ? io_r_163_b : _GEN_10752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10754 = 10'ha4 == r_count_14_io_out ? io_r_164_b : _GEN_10753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10755 = 10'ha5 == r_count_14_io_out ? io_r_165_b : _GEN_10754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10756 = 10'ha6 == r_count_14_io_out ? io_r_166_b : _GEN_10755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10757 = 10'ha7 == r_count_14_io_out ? io_r_167_b : _GEN_10756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10758 = 10'ha8 == r_count_14_io_out ? io_r_168_b : _GEN_10757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10759 = 10'ha9 == r_count_14_io_out ? io_r_169_b : _GEN_10758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10760 = 10'haa == r_count_14_io_out ? io_r_170_b : _GEN_10759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10761 = 10'hab == r_count_14_io_out ? io_r_171_b : _GEN_10760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10762 = 10'hac == r_count_14_io_out ? io_r_172_b : _GEN_10761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10763 = 10'had == r_count_14_io_out ? io_r_173_b : _GEN_10762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10764 = 10'hae == r_count_14_io_out ? io_r_174_b : _GEN_10763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10765 = 10'haf == r_count_14_io_out ? io_r_175_b : _GEN_10764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10766 = 10'hb0 == r_count_14_io_out ? io_r_176_b : _GEN_10765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10767 = 10'hb1 == r_count_14_io_out ? io_r_177_b : _GEN_10766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10768 = 10'hb2 == r_count_14_io_out ? io_r_178_b : _GEN_10767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10769 = 10'hb3 == r_count_14_io_out ? io_r_179_b : _GEN_10768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10770 = 10'hb4 == r_count_14_io_out ? io_r_180_b : _GEN_10769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10771 = 10'hb5 == r_count_14_io_out ? io_r_181_b : _GEN_10770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10772 = 10'hb6 == r_count_14_io_out ? io_r_182_b : _GEN_10771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10773 = 10'hb7 == r_count_14_io_out ? io_r_183_b : _GEN_10772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10774 = 10'hb8 == r_count_14_io_out ? io_r_184_b : _GEN_10773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10775 = 10'hb9 == r_count_14_io_out ? io_r_185_b : _GEN_10774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10776 = 10'hba == r_count_14_io_out ? io_r_186_b : _GEN_10775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10777 = 10'hbb == r_count_14_io_out ? io_r_187_b : _GEN_10776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10778 = 10'hbc == r_count_14_io_out ? io_r_188_b : _GEN_10777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10779 = 10'hbd == r_count_14_io_out ? io_r_189_b : _GEN_10778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10780 = 10'hbe == r_count_14_io_out ? io_r_190_b : _GEN_10779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10781 = 10'hbf == r_count_14_io_out ? io_r_191_b : _GEN_10780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10782 = 10'hc0 == r_count_14_io_out ? io_r_192_b : _GEN_10781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10783 = 10'hc1 == r_count_14_io_out ? io_r_193_b : _GEN_10782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10784 = 10'hc2 == r_count_14_io_out ? io_r_194_b : _GEN_10783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10785 = 10'hc3 == r_count_14_io_out ? io_r_195_b : _GEN_10784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10786 = 10'hc4 == r_count_14_io_out ? io_r_196_b : _GEN_10785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10787 = 10'hc5 == r_count_14_io_out ? io_r_197_b : _GEN_10786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10788 = 10'hc6 == r_count_14_io_out ? io_r_198_b : _GEN_10787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10789 = 10'hc7 == r_count_14_io_out ? io_r_199_b : _GEN_10788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10790 = 10'hc8 == r_count_14_io_out ? io_r_200_b : _GEN_10789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10791 = 10'hc9 == r_count_14_io_out ? io_r_201_b : _GEN_10790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10792 = 10'hca == r_count_14_io_out ? io_r_202_b : _GEN_10791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10793 = 10'hcb == r_count_14_io_out ? io_r_203_b : _GEN_10792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10794 = 10'hcc == r_count_14_io_out ? io_r_204_b : _GEN_10793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10795 = 10'hcd == r_count_14_io_out ? io_r_205_b : _GEN_10794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10796 = 10'hce == r_count_14_io_out ? io_r_206_b : _GEN_10795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10797 = 10'hcf == r_count_14_io_out ? io_r_207_b : _GEN_10796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10798 = 10'hd0 == r_count_14_io_out ? io_r_208_b : _GEN_10797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10799 = 10'hd1 == r_count_14_io_out ? io_r_209_b : _GEN_10798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10800 = 10'hd2 == r_count_14_io_out ? io_r_210_b : _GEN_10799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10801 = 10'hd3 == r_count_14_io_out ? io_r_211_b : _GEN_10800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10802 = 10'hd4 == r_count_14_io_out ? io_r_212_b : _GEN_10801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10803 = 10'hd5 == r_count_14_io_out ? io_r_213_b : _GEN_10802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10804 = 10'hd6 == r_count_14_io_out ? io_r_214_b : _GEN_10803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10805 = 10'hd7 == r_count_14_io_out ? io_r_215_b : _GEN_10804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10806 = 10'hd8 == r_count_14_io_out ? io_r_216_b : _GEN_10805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10807 = 10'hd9 == r_count_14_io_out ? io_r_217_b : _GEN_10806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10808 = 10'hda == r_count_14_io_out ? io_r_218_b : _GEN_10807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10809 = 10'hdb == r_count_14_io_out ? io_r_219_b : _GEN_10808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10810 = 10'hdc == r_count_14_io_out ? io_r_220_b : _GEN_10809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10811 = 10'hdd == r_count_14_io_out ? io_r_221_b : _GEN_10810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10812 = 10'hde == r_count_14_io_out ? io_r_222_b : _GEN_10811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10813 = 10'hdf == r_count_14_io_out ? io_r_223_b : _GEN_10812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10814 = 10'he0 == r_count_14_io_out ? io_r_224_b : _GEN_10813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10815 = 10'he1 == r_count_14_io_out ? io_r_225_b : _GEN_10814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10816 = 10'he2 == r_count_14_io_out ? io_r_226_b : _GEN_10815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10817 = 10'he3 == r_count_14_io_out ? io_r_227_b : _GEN_10816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10818 = 10'he4 == r_count_14_io_out ? io_r_228_b : _GEN_10817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10819 = 10'he5 == r_count_14_io_out ? io_r_229_b : _GEN_10818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10820 = 10'he6 == r_count_14_io_out ? io_r_230_b : _GEN_10819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10821 = 10'he7 == r_count_14_io_out ? io_r_231_b : _GEN_10820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10822 = 10'he8 == r_count_14_io_out ? io_r_232_b : _GEN_10821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10823 = 10'he9 == r_count_14_io_out ? io_r_233_b : _GEN_10822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10824 = 10'hea == r_count_14_io_out ? io_r_234_b : _GEN_10823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10825 = 10'heb == r_count_14_io_out ? io_r_235_b : _GEN_10824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10826 = 10'hec == r_count_14_io_out ? io_r_236_b : _GEN_10825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10827 = 10'hed == r_count_14_io_out ? io_r_237_b : _GEN_10826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10828 = 10'hee == r_count_14_io_out ? io_r_238_b : _GEN_10827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10829 = 10'hef == r_count_14_io_out ? io_r_239_b : _GEN_10828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10830 = 10'hf0 == r_count_14_io_out ? io_r_240_b : _GEN_10829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10831 = 10'hf1 == r_count_14_io_out ? io_r_241_b : _GEN_10830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10832 = 10'hf2 == r_count_14_io_out ? io_r_242_b : _GEN_10831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10833 = 10'hf3 == r_count_14_io_out ? io_r_243_b : _GEN_10832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10834 = 10'hf4 == r_count_14_io_out ? io_r_244_b : _GEN_10833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10835 = 10'hf5 == r_count_14_io_out ? io_r_245_b : _GEN_10834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10836 = 10'hf6 == r_count_14_io_out ? io_r_246_b : _GEN_10835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10837 = 10'hf7 == r_count_14_io_out ? io_r_247_b : _GEN_10836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10838 = 10'hf8 == r_count_14_io_out ? io_r_248_b : _GEN_10837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10839 = 10'hf9 == r_count_14_io_out ? io_r_249_b : _GEN_10838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10840 = 10'hfa == r_count_14_io_out ? io_r_250_b : _GEN_10839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10841 = 10'hfb == r_count_14_io_out ? io_r_251_b : _GEN_10840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10842 = 10'hfc == r_count_14_io_out ? io_r_252_b : _GEN_10841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10843 = 10'hfd == r_count_14_io_out ? io_r_253_b : _GEN_10842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10844 = 10'hfe == r_count_14_io_out ? io_r_254_b : _GEN_10843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10845 = 10'hff == r_count_14_io_out ? io_r_255_b : _GEN_10844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10846 = 10'h100 == r_count_14_io_out ? io_r_256_b : _GEN_10845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10847 = 10'h101 == r_count_14_io_out ? io_r_257_b : _GEN_10846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10848 = 10'h102 == r_count_14_io_out ? io_r_258_b : _GEN_10847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10849 = 10'h103 == r_count_14_io_out ? io_r_259_b : _GEN_10848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10850 = 10'h104 == r_count_14_io_out ? io_r_260_b : _GEN_10849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10851 = 10'h105 == r_count_14_io_out ? io_r_261_b : _GEN_10850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10852 = 10'h106 == r_count_14_io_out ? io_r_262_b : _GEN_10851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10853 = 10'h107 == r_count_14_io_out ? io_r_263_b : _GEN_10852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10854 = 10'h108 == r_count_14_io_out ? io_r_264_b : _GEN_10853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10855 = 10'h109 == r_count_14_io_out ? io_r_265_b : _GEN_10854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10856 = 10'h10a == r_count_14_io_out ? io_r_266_b : _GEN_10855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10857 = 10'h10b == r_count_14_io_out ? io_r_267_b : _GEN_10856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10858 = 10'h10c == r_count_14_io_out ? io_r_268_b : _GEN_10857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10859 = 10'h10d == r_count_14_io_out ? io_r_269_b : _GEN_10858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10860 = 10'h10e == r_count_14_io_out ? io_r_270_b : _GEN_10859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10861 = 10'h10f == r_count_14_io_out ? io_r_271_b : _GEN_10860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10862 = 10'h110 == r_count_14_io_out ? io_r_272_b : _GEN_10861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10863 = 10'h111 == r_count_14_io_out ? io_r_273_b : _GEN_10862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10864 = 10'h112 == r_count_14_io_out ? io_r_274_b : _GEN_10863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10865 = 10'h113 == r_count_14_io_out ? io_r_275_b : _GEN_10864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10866 = 10'h114 == r_count_14_io_out ? io_r_276_b : _GEN_10865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10867 = 10'h115 == r_count_14_io_out ? io_r_277_b : _GEN_10866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10868 = 10'h116 == r_count_14_io_out ? io_r_278_b : _GEN_10867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10869 = 10'h117 == r_count_14_io_out ? io_r_279_b : _GEN_10868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10870 = 10'h118 == r_count_14_io_out ? io_r_280_b : _GEN_10869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10871 = 10'h119 == r_count_14_io_out ? io_r_281_b : _GEN_10870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10872 = 10'h11a == r_count_14_io_out ? io_r_282_b : _GEN_10871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10873 = 10'h11b == r_count_14_io_out ? io_r_283_b : _GEN_10872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10874 = 10'h11c == r_count_14_io_out ? io_r_284_b : _GEN_10873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10875 = 10'h11d == r_count_14_io_out ? io_r_285_b : _GEN_10874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10876 = 10'h11e == r_count_14_io_out ? io_r_286_b : _GEN_10875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10877 = 10'h11f == r_count_14_io_out ? io_r_287_b : _GEN_10876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10878 = 10'h120 == r_count_14_io_out ? io_r_288_b : _GEN_10877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10879 = 10'h121 == r_count_14_io_out ? io_r_289_b : _GEN_10878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10880 = 10'h122 == r_count_14_io_out ? io_r_290_b : _GEN_10879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10881 = 10'h123 == r_count_14_io_out ? io_r_291_b : _GEN_10880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10882 = 10'h124 == r_count_14_io_out ? io_r_292_b : _GEN_10881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10883 = 10'h125 == r_count_14_io_out ? io_r_293_b : _GEN_10882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10884 = 10'h126 == r_count_14_io_out ? io_r_294_b : _GEN_10883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10885 = 10'h127 == r_count_14_io_out ? io_r_295_b : _GEN_10884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10886 = 10'h128 == r_count_14_io_out ? io_r_296_b : _GEN_10885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10887 = 10'h129 == r_count_14_io_out ? io_r_297_b : _GEN_10886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10888 = 10'h12a == r_count_14_io_out ? io_r_298_b : _GEN_10887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10889 = 10'h12b == r_count_14_io_out ? io_r_299_b : _GEN_10888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10890 = 10'h12c == r_count_14_io_out ? io_r_300_b : _GEN_10889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10891 = 10'h12d == r_count_14_io_out ? io_r_301_b : _GEN_10890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10892 = 10'h12e == r_count_14_io_out ? io_r_302_b : _GEN_10891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10893 = 10'h12f == r_count_14_io_out ? io_r_303_b : _GEN_10892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10894 = 10'h130 == r_count_14_io_out ? io_r_304_b : _GEN_10893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10895 = 10'h131 == r_count_14_io_out ? io_r_305_b : _GEN_10894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10896 = 10'h132 == r_count_14_io_out ? io_r_306_b : _GEN_10895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10897 = 10'h133 == r_count_14_io_out ? io_r_307_b : _GEN_10896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10898 = 10'h134 == r_count_14_io_out ? io_r_308_b : _GEN_10897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10899 = 10'h135 == r_count_14_io_out ? io_r_309_b : _GEN_10898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10900 = 10'h136 == r_count_14_io_out ? io_r_310_b : _GEN_10899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10901 = 10'h137 == r_count_14_io_out ? io_r_311_b : _GEN_10900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10902 = 10'h138 == r_count_14_io_out ? io_r_312_b : _GEN_10901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10903 = 10'h139 == r_count_14_io_out ? io_r_313_b : _GEN_10902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10904 = 10'h13a == r_count_14_io_out ? io_r_314_b : _GEN_10903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10905 = 10'h13b == r_count_14_io_out ? io_r_315_b : _GEN_10904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10906 = 10'h13c == r_count_14_io_out ? io_r_316_b : _GEN_10905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10907 = 10'h13d == r_count_14_io_out ? io_r_317_b : _GEN_10906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10908 = 10'h13e == r_count_14_io_out ? io_r_318_b : _GEN_10907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10909 = 10'h13f == r_count_14_io_out ? io_r_319_b : _GEN_10908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10910 = 10'h140 == r_count_14_io_out ? io_r_320_b : _GEN_10909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10911 = 10'h141 == r_count_14_io_out ? io_r_321_b : _GEN_10910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10912 = 10'h142 == r_count_14_io_out ? io_r_322_b : _GEN_10911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10913 = 10'h143 == r_count_14_io_out ? io_r_323_b : _GEN_10912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10914 = 10'h144 == r_count_14_io_out ? io_r_324_b : _GEN_10913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10915 = 10'h145 == r_count_14_io_out ? io_r_325_b : _GEN_10914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10916 = 10'h146 == r_count_14_io_out ? io_r_326_b : _GEN_10915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10917 = 10'h147 == r_count_14_io_out ? io_r_327_b : _GEN_10916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10918 = 10'h148 == r_count_14_io_out ? io_r_328_b : _GEN_10917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10919 = 10'h149 == r_count_14_io_out ? io_r_329_b : _GEN_10918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10920 = 10'h14a == r_count_14_io_out ? io_r_330_b : _GEN_10919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10921 = 10'h14b == r_count_14_io_out ? io_r_331_b : _GEN_10920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10922 = 10'h14c == r_count_14_io_out ? io_r_332_b : _GEN_10921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10923 = 10'h14d == r_count_14_io_out ? io_r_333_b : _GEN_10922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10924 = 10'h14e == r_count_14_io_out ? io_r_334_b : _GEN_10923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10925 = 10'h14f == r_count_14_io_out ? io_r_335_b : _GEN_10924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10926 = 10'h150 == r_count_14_io_out ? io_r_336_b : _GEN_10925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10927 = 10'h151 == r_count_14_io_out ? io_r_337_b : _GEN_10926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10928 = 10'h152 == r_count_14_io_out ? io_r_338_b : _GEN_10927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10929 = 10'h153 == r_count_14_io_out ? io_r_339_b : _GEN_10928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10930 = 10'h154 == r_count_14_io_out ? io_r_340_b : _GEN_10929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10931 = 10'h155 == r_count_14_io_out ? io_r_341_b : _GEN_10930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10932 = 10'h156 == r_count_14_io_out ? io_r_342_b : _GEN_10931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10933 = 10'h157 == r_count_14_io_out ? io_r_343_b : _GEN_10932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10934 = 10'h158 == r_count_14_io_out ? io_r_344_b : _GEN_10933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10935 = 10'h159 == r_count_14_io_out ? io_r_345_b : _GEN_10934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10936 = 10'h15a == r_count_14_io_out ? io_r_346_b : _GEN_10935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10937 = 10'h15b == r_count_14_io_out ? io_r_347_b : _GEN_10936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10938 = 10'h15c == r_count_14_io_out ? io_r_348_b : _GEN_10937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10939 = 10'h15d == r_count_14_io_out ? io_r_349_b : _GEN_10938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10940 = 10'h15e == r_count_14_io_out ? io_r_350_b : _GEN_10939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10941 = 10'h15f == r_count_14_io_out ? io_r_351_b : _GEN_10940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10942 = 10'h160 == r_count_14_io_out ? io_r_352_b : _GEN_10941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10943 = 10'h161 == r_count_14_io_out ? io_r_353_b : _GEN_10942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10944 = 10'h162 == r_count_14_io_out ? io_r_354_b : _GEN_10943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10945 = 10'h163 == r_count_14_io_out ? io_r_355_b : _GEN_10944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10946 = 10'h164 == r_count_14_io_out ? io_r_356_b : _GEN_10945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10947 = 10'h165 == r_count_14_io_out ? io_r_357_b : _GEN_10946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10948 = 10'h166 == r_count_14_io_out ? io_r_358_b : _GEN_10947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10949 = 10'h167 == r_count_14_io_out ? io_r_359_b : _GEN_10948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10950 = 10'h168 == r_count_14_io_out ? io_r_360_b : _GEN_10949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10951 = 10'h169 == r_count_14_io_out ? io_r_361_b : _GEN_10950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10952 = 10'h16a == r_count_14_io_out ? io_r_362_b : _GEN_10951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10953 = 10'h16b == r_count_14_io_out ? io_r_363_b : _GEN_10952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10954 = 10'h16c == r_count_14_io_out ? io_r_364_b : _GEN_10953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10955 = 10'h16d == r_count_14_io_out ? io_r_365_b : _GEN_10954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10956 = 10'h16e == r_count_14_io_out ? io_r_366_b : _GEN_10955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10957 = 10'h16f == r_count_14_io_out ? io_r_367_b : _GEN_10956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10958 = 10'h170 == r_count_14_io_out ? io_r_368_b : _GEN_10957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10959 = 10'h171 == r_count_14_io_out ? io_r_369_b : _GEN_10958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10960 = 10'h172 == r_count_14_io_out ? io_r_370_b : _GEN_10959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10961 = 10'h173 == r_count_14_io_out ? io_r_371_b : _GEN_10960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10962 = 10'h174 == r_count_14_io_out ? io_r_372_b : _GEN_10961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10963 = 10'h175 == r_count_14_io_out ? io_r_373_b : _GEN_10962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10964 = 10'h176 == r_count_14_io_out ? io_r_374_b : _GEN_10963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10965 = 10'h177 == r_count_14_io_out ? io_r_375_b : _GEN_10964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10966 = 10'h178 == r_count_14_io_out ? io_r_376_b : _GEN_10965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10967 = 10'h179 == r_count_14_io_out ? io_r_377_b : _GEN_10966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10968 = 10'h17a == r_count_14_io_out ? io_r_378_b : _GEN_10967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10969 = 10'h17b == r_count_14_io_out ? io_r_379_b : _GEN_10968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10970 = 10'h17c == r_count_14_io_out ? io_r_380_b : _GEN_10969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10971 = 10'h17d == r_count_14_io_out ? io_r_381_b : _GEN_10970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10972 = 10'h17e == r_count_14_io_out ? io_r_382_b : _GEN_10971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10973 = 10'h17f == r_count_14_io_out ? io_r_383_b : _GEN_10972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10974 = 10'h180 == r_count_14_io_out ? io_r_384_b : _GEN_10973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10975 = 10'h181 == r_count_14_io_out ? io_r_385_b : _GEN_10974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10976 = 10'h182 == r_count_14_io_out ? io_r_386_b : _GEN_10975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10977 = 10'h183 == r_count_14_io_out ? io_r_387_b : _GEN_10976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10978 = 10'h184 == r_count_14_io_out ? io_r_388_b : _GEN_10977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10979 = 10'h185 == r_count_14_io_out ? io_r_389_b : _GEN_10978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10980 = 10'h186 == r_count_14_io_out ? io_r_390_b : _GEN_10979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10981 = 10'h187 == r_count_14_io_out ? io_r_391_b : _GEN_10980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10982 = 10'h188 == r_count_14_io_out ? io_r_392_b : _GEN_10981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10983 = 10'h189 == r_count_14_io_out ? io_r_393_b : _GEN_10982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10984 = 10'h18a == r_count_14_io_out ? io_r_394_b : _GEN_10983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10985 = 10'h18b == r_count_14_io_out ? io_r_395_b : _GEN_10984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10986 = 10'h18c == r_count_14_io_out ? io_r_396_b : _GEN_10985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10987 = 10'h18d == r_count_14_io_out ? io_r_397_b : _GEN_10986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10988 = 10'h18e == r_count_14_io_out ? io_r_398_b : _GEN_10987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10989 = 10'h18f == r_count_14_io_out ? io_r_399_b : _GEN_10988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10990 = 10'h190 == r_count_14_io_out ? io_r_400_b : _GEN_10989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10991 = 10'h191 == r_count_14_io_out ? io_r_401_b : _GEN_10990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10992 = 10'h192 == r_count_14_io_out ? io_r_402_b : _GEN_10991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10993 = 10'h193 == r_count_14_io_out ? io_r_403_b : _GEN_10992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10994 = 10'h194 == r_count_14_io_out ? io_r_404_b : _GEN_10993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10995 = 10'h195 == r_count_14_io_out ? io_r_405_b : _GEN_10994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10996 = 10'h196 == r_count_14_io_out ? io_r_406_b : _GEN_10995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10997 = 10'h197 == r_count_14_io_out ? io_r_407_b : _GEN_10996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10998 = 10'h198 == r_count_14_io_out ? io_r_408_b : _GEN_10997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10999 = 10'h199 == r_count_14_io_out ? io_r_409_b : _GEN_10998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11000 = 10'h19a == r_count_14_io_out ? io_r_410_b : _GEN_10999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11001 = 10'h19b == r_count_14_io_out ? io_r_411_b : _GEN_11000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11002 = 10'h19c == r_count_14_io_out ? io_r_412_b : _GEN_11001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11003 = 10'h19d == r_count_14_io_out ? io_r_413_b : _GEN_11002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11004 = 10'h19e == r_count_14_io_out ? io_r_414_b : _GEN_11003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11005 = 10'h19f == r_count_14_io_out ? io_r_415_b : _GEN_11004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11006 = 10'h1a0 == r_count_14_io_out ? io_r_416_b : _GEN_11005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11007 = 10'h1a1 == r_count_14_io_out ? io_r_417_b : _GEN_11006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11008 = 10'h1a2 == r_count_14_io_out ? io_r_418_b : _GEN_11007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11009 = 10'h1a3 == r_count_14_io_out ? io_r_419_b : _GEN_11008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11010 = 10'h1a4 == r_count_14_io_out ? io_r_420_b : _GEN_11009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11011 = 10'h1a5 == r_count_14_io_out ? io_r_421_b : _GEN_11010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11012 = 10'h1a6 == r_count_14_io_out ? io_r_422_b : _GEN_11011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11013 = 10'h1a7 == r_count_14_io_out ? io_r_423_b : _GEN_11012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11014 = 10'h1a8 == r_count_14_io_out ? io_r_424_b : _GEN_11013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11015 = 10'h1a9 == r_count_14_io_out ? io_r_425_b : _GEN_11014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11016 = 10'h1aa == r_count_14_io_out ? io_r_426_b : _GEN_11015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11017 = 10'h1ab == r_count_14_io_out ? io_r_427_b : _GEN_11016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11018 = 10'h1ac == r_count_14_io_out ? io_r_428_b : _GEN_11017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11019 = 10'h1ad == r_count_14_io_out ? io_r_429_b : _GEN_11018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11020 = 10'h1ae == r_count_14_io_out ? io_r_430_b : _GEN_11019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11021 = 10'h1af == r_count_14_io_out ? io_r_431_b : _GEN_11020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11022 = 10'h1b0 == r_count_14_io_out ? io_r_432_b : _GEN_11021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11023 = 10'h1b1 == r_count_14_io_out ? io_r_433_b : _GEN_11022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11024 = 10'h1b2 == r_count_14_io_out ? io_r_434_b : _GEN_11023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11025 = 10'h1b3 == r_count_14_io_out ? io_r_435_b : _GEN_11024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11026 = 10'h1b4 == r_count_14_io_out ? io_r_436_b : _GEN_11025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11027 = 10'h1b5 == r_count_14_io_out ? io_r_437_b : _GEN_11026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11028 = 10'h1b6 == r_count_14_io_out ? io_r_438_b : _GEN_11027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11029 = 10'h1b7 == r_count_14_io_out ? io_r_439_b : _GEN_11028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11030 = 10'h1b8 == r_count_14_io_out ? io_r_440_b : _GEN_11029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11031 = 10'h1b9 == r_count_14_io_out ? io_r_441_b : _GEN_11030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11032 = 10'h1ba == r_count_14_io_out ? io_r_442_b : _GEN_11031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11033 = 10'h1bb == r_count_14_io_out ? io_r_443_b : _GEN_11032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11034 = 10'h1bc == r_count_14_io_out ? io_r_444_b : _GEN_11033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11035 = 10'h1bd == r_count_14_io_out ? io_r_445_b : _GEN_11034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11036 = 10'h1be == r_count_14_io_out ? io_r_446_b : _GEN_11035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11037 = 10'h1bf == r_count_14_io_out ? io_r_447_b : _GEN_11036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11038 = 10'h1c0 == r_count_14_io_out ? io_r_448_b : _GEN_11037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11039 = 10'h1c1 == r_count_14_io_out ? io_r_449_b : _GEN_11038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11040 = 10'h1c2 == r_count_14_io_out ? io_r_450_b : _GEN_11039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11041 = 10'h1c3 == r_count_14_io_out ? io_r_451_b : _GEN_11040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11042 = 10'h1c4 == r_count_14_io_out ? io_r_452_b : _GEN_11041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11043 = 10'h1c5 == r_count_14_io_out ? io_r_453_b : _GEN_11042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11044 = 10'h1c6 == r_count_14_io_out ? io_r_454_b : _GEN_11043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11045 = 10'h1c7 == r_count_14_io_out ? io_r_455_b : _GEN_11044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11046 = 10'h1c8 == r_count_14_io_out ? io_r_456_b : _GEN_11045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11047 = 10'h1c9 == r_count_14_io_out ? io_r_457_b : _GEN_11046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11048 = 10'h1ca == r_count_14_io_out ? io_r_458_b : _GEN_11047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11049 = 10'h1cb == r_count_14_io_out ? io_r_459_b : _GEN_11048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11050 = 10'h1cc == r_count_14_io_out ? io_r_460_b : _GEN_11049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11051 = 10'h1cd == r_count_14_io_out ? io_r_461_b : _GEN_11050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11052 = 10'h1ce == r_count_14_io_out ? io_r_462_b : _GEN_11051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11053 = 10'h1cf == r_count_14_io_out ? io_r_463_b : _GEN_11052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11054 = 10'h1d0 == r_count_14_io_out ? io_r_464_b : _GEN_11053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11055 = 10'h1d1 == r_count_14_io_out ? io_r_465_b : _GEN_11054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11056 = 10'h1d2 == r_count_14_io_out ? io_r_466_b : _GEN_11055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11057 = 10'h1d3 == r_count_14_io_out ? io_r_467_b : _GEN_11056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11058 = 10'h1d4 == r_count_14_io_out ? io_r_468_b : _GEN_11057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11059 = 10'h1d5 == r_count_14_io_out ? io_r_469_b : _GEN_11058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11060 = 10'h1d6 == r_count_14_io_out ? io_r_470_b : _GEN_11059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11061 = 10'h1d7 == r_count_14_io_out ? io_r_471_b : _GEN_11060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11062 = 10'h1d8 == r_count_14_io_out ? io_r_472_b : _GEN_11061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11063 = 10'h1d9 == r_count_14_io_out ? io_r_473_b : _GEN_11062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11064 = 10'h1da == r_count_14_io_out ? io_r_474_b : _GEN_11063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11065 = 10'h1db == r_count_14_io_out ? io_r_475_b : _GEN_11064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11066 = 10'h1dc == r_count_14_io_out ? io_r_476_b : _GEN_11065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11067 = 10'h1dd == r_count_14_io_out ? io_r_477_b : _GEN_11066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11068 = 10'h1de == r_count_14_io_out ? io_r_478_b : _GEN_11067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11069 = 10'h1df == r_count_14_io_out ? io_r_479_b : _GEN_11068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11070 = 10'h1e0 == r_count_14_io_out ? io_r_480_b : _GEN_11069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11071 = 10'h1e1 == r_count_14_io_out ? io_r_481_b : _GEN_11070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11072 = 10'h1e2 == r_count_14_io_out ? io_r_482_b : _GEN_11071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11073 = 10'h1e3 == r_count_14_io_out ? io_r_483_b : _GEN_11072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11074 = 10'h1e4 == r_count_14_io_out ? io_r_484_b : _GEN_11073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11075 = 10'h1e5 == r_count_14_io_out ? io_r_485_b : _GEN_11074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11076 = 10'h1e6 == r_count_14_io_out ? io_r_486_b : _GEN_11075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11077 = 10'h1e7 == r_count_14_io_out ? io_r_487_b : _GEN_11076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11078 = 10'h1e8 == r_count_14_io_out ? io_r_488_b : _GEN_11077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11079 = 10'h1e9 == r_count_14_io_out ? io_r_489_b : _GEN_11078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11080 = 10'h1ea == r_count_14_io_out ? io_r_490_b : _GEN_11079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11081 = 10'h1eb == r_count_14_io_out ? io_r_491_b : _GEN_11080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11082 = 10'h1ec == r_count_14_io_out ? io_r_492_b : _GEN_11081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11083 = 10'h1ed == r_count_14_io_out ? io_r_493_b : _GEN_11082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11084 = 10'h1ee == r_count_14_io_out ? io_r_494_b : _GEN_11083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11085 = 10'h1ef == r_count_14_io_out ? io_r_495_b : _GEN_11084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11086 = 10'h1f0 == r_count_14_io_out ? io_r_496_b : _GEN_11085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11087 = 10'h1f1 == r_count_14_io_out ? io_r_497_b : _GEN_11086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11088 = 10'h1f2 == r_count_14_io_out ? io_r_498_b : _GEN_11087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11089 = 10'h1f3 == r_count_14_io_out ? io_r_499_b : _GEN_11088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11090 = 10'h1f4 == r_count_14_io_out ? io_r_500_b : _GEN_11089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11091 = 10'h1f5 == r_count_14_io_out ? io_r_501_b : _GEN_11090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11092 = 10'h1f6 == r_count_14_io_out ? io_r_502_b : _GEN_11091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11093 = 10'h1f7 == r_count_14_io_out ? io_r_503_b : _GEN_11092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11094 = 10'h1f8 == r_count_14_io_out ? io_r_504_b : _GEN_11093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11095 = 10'h1f9 == r_count_14_io_out ? io_r_505_b : _GEN_11094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11096 = 10'h1fa == r_count_14_io_out ? io_r_506_b : _GEN_11095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11097 = 10'h1fb == r_count_14_io_out ? io_r_507_b : _GEN_11096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11098 = 10'h1fc == r_count_14_io_out ? io_r_508_b : _GEN_11097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11099 = 10'h1fd == r_count_14_io_out ? io_r_509_b : _GEN_11098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11100 = 10'h1fe == r_count_14_io_out ? io_r_510_b : _GEN_11099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11101 = 10'h1ff == r_count_14_io_out ? io_r_511_b : _GEN_11100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11102 = 10'h200 == r_count_14_io_out ? io_r_512_b : _GEN_11101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11103 = 10'h201 == r_count_14_io_out ? io_r_513_b : _GEN_11102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11104 = 10'h202 == r_count_14_io_out ? io_r_514_b : _GEN_11103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11105 = 10'h203 == r_count_14_io_out ? io_r_515_b : _GEN_11104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11106 = 10'h204 == r_count_14_io_out ? io_r_516_b : _GEN_11105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11107 = 10'h205 == r_count_14_io_out ? io_r_517_b : _GEN_11106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11108 = 10'h206 == r_count_14_io_out ? io_r_518_b : _GEN_11107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11109 = 10'h207 == r_count_14_io_out ? io_r_519_b : _GEN_11108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11110 = 10'h208 == r_count_14_io_out ? io_r_520_b : _GEN_11109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11111 = 10'h209 == r_count_14_io_out ? io_r_521_b : _GEN_11110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11112 = 10'h20a == r_count_14_io_out ? io_r_522_b : _GEN_11111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11113 = 10'h20b == r_count_14_io_out ? io_r_523_b : _GEN_11112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11114 = 10'h20c == r_count_14_io_out ? io_r_524_b : _GEN_11113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11115 = 10'h20d == r_count_14_io_out ? io_r_525_b : _GEN_11114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11116 = 10'h20e == r_count_14_io_out ? io_r_526_b : _GEN_11115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11117 = 10'h20f == r_count_14_io_out ? io_r_527_b : _GEN_11116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11118 = 10'h210 == r_count_14_io_out ? io_r_528_b : _GEN_11117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11119 = 10'h211 == r_count_14_io_out ? io_r_529_b : _GEN_11118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11120 = 10'h212 == r_count_14_io_out ? io_r_530_b : _GEN_11119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11121 = 10'h213 == r_count_14_io_out ? io_r_531_b : _GEN_11120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11122 = 10'h214 == r_count_14_io_out ? io_r_532_b : _GEN_11121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11123 = 10'h215 == r_count_14_io_out ? io_r_533_b : _GEN_11122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11124 = 10'h216 == r_count_14_io_out ? io_r_534_b : _GEN_11123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11125 = 10'h217 == r_count_14_io_out ? io_r_535_b : _GEN_11124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11126 = 10'h218 == r_count_14_io_out ? io_r_536_b : _GEN_11125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11127 = 10'h219 == r_count_14_io_out ? io_r_537_b : _GEN_11126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11128 = 10'h21a == r_count_14_io_out ? io_r_538_b : _GEN_11127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11129 = 10'h21b == r_count_14_io_out ? io_r_539_b : _GEN_11128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11130 = 10'h21c == r_count_14_io_out ? io_r_540_b : _GEN_11129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11131 = 10'h21d == r_count_14_io_out ? io_r_541_b : _GEN_11130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11132 = 10'h21e == r_count_14_io_out ? io_r_542_b : _GEN_11131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11133 = 10'h21f == r_count_14_io_out ? io_r_543_b : _GEN_11132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11134 = 10'h220 == r_count_14_io_out ? io_r_544_b : _GEN_11133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11135 = 10'h221 == r_count_14_io_out ? io_r_545_b : _GEN_11134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11136 = 10'h222 == r_count_14_io_out ? io_r_546_b : _GEN_11135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11137 = 10'h223 == r_count_14_io_out ? io_r_547_b : _GEN_11136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11138 = 10'h224 == r_count_14_io_out ? io_r_548_b : _GEN_11137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11139 = 10'h225 == r_count_14_io_out ? io_r_549_b : _GEN_11138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11140 = 10'h226 == r_count_14_io_out ? io_r_550_b : _GEN_11139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11141 = 10'h227 == r_count_14_io_out ? io_r_551_b : _GEN_11140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11142 = 10'h228 == r_count_14_io_out ? io_r_552_b : _GEN_11141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11143 = 10'h229 == r_count_14_io_out ? io_r_553_b : _GEN_11142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11144 = 10'h22a == r_count_14_io_out ? io_r_554_b : _GEN_11143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11145 = 10'h22b == r_count_14_io_out ? io_r_555_b : _GEN_11144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11146 = 10'h22c == r_count_14_io_out ? io_r_556_b : _GEN_11145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11147 = 10'h22d == r_count_14_io_out ? io_r_557_b : _GEN_11146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11148 = 10'h22e == r_count_14_io_out ? io_r_558_b : _GEN_11147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11149 = 10'h22f == r_count_14_io_out ? io_r_559_b : _GEN_11148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11150 = 10'h230 == r_count_14_io_out ? io_r_560_b : _GEN_11149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11151 = 10'h231 == r_count_14_io_out ? io_r_561_b : _GEN_11150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11152 = 10'h232 == r_count_14_io_out ? io_r_562_b : _GEN_11151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11153 = 10'h233 == r_count_14_io_out ? io_r_563_b : _GEN_11152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11154 = 10'h234 == r_count_14_io_out ? io_r_564_b : _GEN_11153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11155 = 10'h235 == r_count_14_io_out ? io_r_565_b : _GEN_11154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11156 = 10'h236 == r_count_14_io_out ? io_r_566_b : _GEN_11155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11157 = 10'h237 == r_count_14_io_out ? io_r_567_b : _GEN_11156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11158 = 10'h238 == r_count_14_io_out ? io_r_568_b : _GEN_11157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11159 = 10'h239 == r_count_14_io_out ? io_r_569_b : _GEN_11158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11160 = 10'h23a == r_count_14_io_out ? io_r_570_b : _GEN_11159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11161 = 10'h23b == r_count_14_io_out ? io_r_571_b : _GEN_11160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11162 = 10'h23c == r_count_14_io_out ? io_r_572_b : _GEN_11161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11163 = 10'h23d == r_count_14_io_out ? io_r_573_b : _GEN_11162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11164 = 10'h23e == r_count_14_io_out ? io_r_574_b : _GEN_11163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11165 = 10'h23f == r_count_14_io_out ? io_r_575_b : _GEN_11164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11166 = 10'h240 == r_count_14_io_out ? io_r_576_b : _GEN_11165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11167 = 10'h241 == r_count_14_io_out ? io_r_577_b : _GEN_11166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11168 = 10'h242 == r_count_14_io_out ? io_r_578_b : _GEN_11167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11169 = 10'h243 == r_count_14_io_out ? io_r_579_b : _GEN_11168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11170 = 10'h244 == r_count_14_io_out ? io_r_580_b : _GEN_11169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11171 = 10'h245 == r_count_14_io_out ? io_r_581_b : _GEN_11170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11172 = 10'h246 == r_count_14_io_out ? io_r_582_b : _GEN_11171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11173 = 10'h247 == r_count_14_io_out ? io_r_583_b : _GEN_11172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11174 = 10'h248 == r_count_14_io_out ? io_r_584_b : _GEN_11173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11175 = 10'h249 == r_count_14_io_out ? io_r_585_b : _GEN_11174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11176 = 10'h24a == r_count_14_io_out ? io_r_586_b : _GEN_11175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11177 = 10'h24b == r_count_14_io_out ? io_r_587_b : _GEN_11176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11178 = 10'h24c == r_count_14_io_out ? io_r_588_b : _GEN_11177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11179 = 10'h24d == r_count_14_io_out ? io_r_589_b : _GEN_11178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11180 = 10'h24e == r_count_14_io_out ? io_r_590_b : _GEN_11179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11181 = 10'h24f == r_count_14_io_out ? io_r_591_b : _GEN_11180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11182 = 10'h250 == r_count_14_io_out ? io_r_592_b : _GEN_11181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11183 = 10'h251 == r_count_14_io_out ? io_r_593_b : _GEN_11182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11184 = 10'h252 == r_count_14_io_out ? io_r_594_b : _GEN_11183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11185 = 10'h253 == r_count_14_io_out ? io_r_595_b : _GEN_11184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11186 = 10'h254 == r_count_14_io_out ? io_r_596_b : _GEN_11185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11187 = 10'h255 == r_count_14_io_out ? io_r_597_b : _GEN_11186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11188 = 10'h256 == r_count_14_io_out ? io_r_598_b : _GEN_11187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11189 = 10'h257 == r_count_14_io_out ? io_r_599_b : _GEN_11188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11190 = 10'h258 == r_count_14_io_out ? io_r_600_b : _GEN_11189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11191 = 10'h259 == r_count_14_io_out ? io_r_601_b : _GEN_11190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11192 = 10'h25a == r_count_14_io_out ? io_r_602_b : _GEN_11191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11193 = 10'h25b == r_count_14_io_out ? io_r_603_b : _GEN_11192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11194 = 10'h25c == r_count_14_io_out ? io_r_604_b : _GEN_11193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11195 = 10'h25d == r_count_14_io_out ? io_r_605_b : _GEN_11194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11196 = 10'h25e == r_count_14_io_out ? io_r_606_b : _GEN_11195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11197 = 10'h25f == r_count_14_io_out ? io_r_607_b : _GEN_11196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11198 = 10'h260 == r_count_14_io_out ? io_r_608_b : _GEN_11197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11199 = 10'h261 == r_count_14_io_out ? io_r_609_b : _GEN_11198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11200 = 10'h262 == r_count_14_io_out ? io_r_610_b : _GEN_11199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11201 = 10'h263 == r_count_14_io_out ? io_r_611_b : _GEN_11200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11202 = 10'h264 == r_count_14_io_out ? io_r_612_b : _GEN_11201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11203 = 10'h265 == r_count_14_io_out ? io_r_613_b : _GEN_11202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11204 = 10'h266 == r_count_14_io_out ? io_r_614_b : _GEN_11203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11205 = 10'h267 == r_count_14_io_out ? io_r_615_b : _GEN_11204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11206 = 10'h268 == r_count_14_io_out ? io_r_616_b : _GEN_11205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11207 = 10'h269 == r_count_14_io_out ? io_r_617_b : _GEN_11206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11208 = 10'h26a == r_count_14_io_out ? io_r_618_b : _GEN_11207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11209 = 10'h26b == r_count_14_io_out ? io_r_619_b : _GEN_11208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11210 = 10'h26c == r_count_14_io_out ? io_r_620_b : _GEN_11209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11211 = 10'h26d == r_count_14_io_out ? io_r_621_b : _GEN_11210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11212 = 10'h26e == r_count_14_io_out ? io_r_622_b : _GEN_11211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11213 = 10'h26f == r_count_14_io_out ? io_r_623_b : _GEN_11212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11214 = 10'h270 == r_count_14_io_out ? io_r_624_b : _GEN_11213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11215 = 10'h271 == r_count_14_io_out ? io_r_625_b : _GEN_11214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11216 = 10'h272 == r_count_14_io_out ? io_r_626_b : _GEN_11215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11217 = 10'h273 == r_count_14_io_out ? io_r_627_b : _GEN_11216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11218 = 10'h274 == r_count_14_io_out ? io_r_628_b : _GEN_11217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11219 = 10'h275 == r_count_14_io_out ? io_r_629_b : _GEN_11218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11220 = 10'h276 == r_count_14_io_out ? io_r_630_b : _GEN_11219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11221 = 10'h277 == r_count_14_io_out ? io_r_631_b : _GEN_11220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11222 = 10'h278 == r_count_14_io_out ? io_r_632_b : _GEN_11221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11223 = 10'h279 == r_count_14_io_out ? io_r_633_b : _GEN_11222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11224 = 10'h27a == r_count_14_io_out ? io_r_634_b : _GEN_11223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11225 = 10'h27b == r_count_14_io_out ? io_r_635_b : _GEN_11224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11226 = 10'h27c == r_count_14_io_out ? io_r_636_b : _GEN_11225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11227 = 10'h27d == r_count_14_io_out ? io_r_637_b : _GEN_11226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11228 = 10'h27e == r_count_14_io_out ? io_r_638_b : _GEN_11227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11229 = 10'h27f == r_count_14_io_out ? io_r_639_b : _GEN_11228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11230 = 10'h280 == r_count_14_io_out ? io_r_640_b : _GEN_11229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11231 = 10'h281 == r_count_14_io_out ? io_r_641_b : _GEN_11230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11232 = 10'h282 == r_count_14_io_out ? io_r_642_b : _GEN_11231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11233 = 10'h283 == r_count_14_io_out ? io_r_643_b : _GEN_11232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11234 = 10'h284 == r_count_14_io_out ? io_r_644_b : _GEN_11233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11235 = 10'h285 == r_count_14_io_out ? io_r_645_b : _GEN_11234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11236 = 10'h286 == r_count_14_io_out ? io_r_646_b : _GEN_11235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11237 = 10'h287 == r_count_14_io_out ? io_r_647_b : _GEN_11236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11238 = 10'h288 == r_count_14_io_out ? io_r_648_b : _GEN_11237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11239 = 10'h289 == r_count_14_io_out ? io_r_649_b : _GEN_11238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11240 = 10'h28a == r_count_14_io_out ? io_r_650_b : _GEN_11239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11241 = 10'h28b == r_count_14_io_out ? io_r_651_b : _GEN_11240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11242 = 10'h28c == r_count_14_io_out ? io_r_652_b : _GEN_11241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11243 = 10'h28d == r_count_14_io_out ? io_r_653_b : _GEN_11242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11244 = 10'h28e == r_count_14_io_out ? io_r_654_b : _GEN_11243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11245 = 10'h28f == r_count_14_io_out ? io_r_655_b : _GEN_11244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11246 = 10'h290 == r_count_14_io_out ? io_r_656_b : _GEN_11245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11247 = 10'h291 == r_count_14_io_out ? io_r_657_b : _GEN_11246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11248 = 10'h292 == r_count_14_io_out ? io_r_658_b : _GEN_11247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11249 = 10'h293 == r_count_14_io_out ? io_r_659_b : _GEN_11248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11250 = 10'h294 == r_count_14_io_out ? io_r_660_b : _GEN_11249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11251 = 10'h295 == r_count_14_io_out ? io_r_661_b : _GEN_11250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11252 = 10'h296 == r_count_14_io_out ? io_r_662_b : _GEN_11251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11253 = 10'h297 == r_count_14_io_out ? io_r_663_b : _GEN_11252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11254 = 10'h298 == r_count_14_io_out ? io_r_664_b : _GEN_11253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11255 = 10'h299 == r_count_14_io_out ? io_r_665_b : _GEN_11254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11256 = 10'h29a == r_count_14_io_out ? io_r_666_b : _GEN_11255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11257 = 10'h29b == r_count_14_io_out ? io_r_667_b : _GEN_11256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11258 = 10'h29c == r_count_14_io_out ? io_r_668_b : _GEN_11257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11259 = 10'h29d == r_count_14_io_out ? io_r_669_b : _GEN_11258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11260 = 10'h29e == r_count_14_io_out ? io_r_670_b : _GEN_11259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11261 = 10'h29f == r_count_14_io_out ? io_r_671_b : _GEN_11260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11262 = 10'h2a0 == r_count_14_io_out ? io_r_672_b : _GEN_11261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11263 = 10'h2a1 == r_count_14_io_out ? io_r_673_b : _GEN_11262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11264 = 10'h2a2 == r_count_14_io_out ? io_r_674_b : _GEN_11263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11265 = 10'h2a3 == r_count_14_io_out ? io_r_675_b : _GEN_11264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11266 = 10'h2a4 == r_count_14_io_out ? io_r_676_b : _GEN_11265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11267 = 10'h2a5 == r_count_14_io_out ? io_r_677_b : _GEN_11266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11268 = 10'h2a6 == r_count_14_io_out ? io_r_678_b : _GEN_11267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11269 = 10'h2a7 == r_count_14_io_out ? io_r_679_b : _GEN_11268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11270 = 10'h2a8 == r_count_14_io_out ? io_r_680_b : _GEN_11269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11271 = 10'h2a9 == r_count_14_io_out ? io_r_681_b : _GEN_11270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11272 = 10'h2aa == r_count_14_io_out ? io_r_682_b : _GEN_11271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11273 = 10'h2ab == r_count_14_io_out ? io_r_683_b : _GEN_11272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11274 = 10'h2ac == r_count_14_io_out ? io_r_684_b : _GEN_11273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11275 = 10'h2ad == r_count_14_io_out ? io_r_685_b : _GEN_11274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11276 = 10'h2ae == r_count_14_io_out ? io_r_686_b : _GEN_11275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11277 = 10'h2af == r_count_14_io_out ? io_r_687_b : _GEN_11276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11278 = 10'h2b0 == r_count_14_io_out ? io_r_688_b : _GEN_11277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11279 = 10'h2b1 == r_count_14_io_out ? io_r_689_b : _GEN_11278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11280 = 10'h2b2 == r_count_14_io_out ? io_r_690_b : _GEN_11279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11281 = 10'h2b3 == r_count_14_io_out ? io_r_691_b : _GEN_11280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11282 = 10'h2b4 == r_count_14_io_out ? io_r_692_b : _GEN_11281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11283 = 10'h2b5 == r_count_14_io_out ? io_r_693_b : _GEN_11282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11284 = 10'h2b6 == r_count_14_io_out ? io_r_694_b : _GEN_11283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11285 = 10'h2b7 == r_count_14_io_out ? io_r_695_b : _GEN_11284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11286 = 10'h2b8 == r_count_14_io_out ? io_r_696_b : _GEN_11285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11287 = 10'h2b9 == r_count_14_io_out ? io_r_697_b : _GEN_11286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11288 = 10'h2ba == r_count_14_io_out ? io_r_698_b : _GEN_11287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11289 = 10'h2bb == r_count_14_io_out ? io_r_699_b : _GEN_11288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11290 = 10'h2bc == r_count_14_io_out ? io_r_700_b : _GEN_11289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11291 = 10'h2bd == r_count_14_io_out ? io_r_701_b : _GEN_11290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11292 = 10'h2be == r_count_14_io_out ? io_r_702_b : _GEN_11291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11293 = 10'h2bf == r_count_14_io_out ? io_r_703_b : _GEN_11292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11294 = 10'h2c0 == r_count_14_io_out ? io_r_704_b : _GEN_11293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11295 = 10'h2c1 == r_count_14_io_out ? io_r_705_b : _GEN_11294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11296 = 10'h2c2 == r_count_14_io_out ? io_r_706_b : _GEN_11295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11297 = 10'h2c3 == r_count_14_io_out ? io_r_707_b : _GEN_11296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11298 = 10'h2c4 == r_count_14_io_out ? io_r_708_b : _GEN_11297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11299 = 10'h2c5 == r_count_14_io_out ? io_r_709_b : _GEN_11298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11300 = 10'h2c6 == r_count_14_io_out ? io_r_710_b : _GEN_11299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11301 = 10'h2c7 == r_count_14_io_out ? io_r_711_b : _GEN_11300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11302 = 10'h2c8 == r_count_14_io_out ? io_r_712_b : _GEN_11301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11303 = 10'h2c9 == r_count_14_io_out ? io_r_713_b : _GEN_11302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11304 = 10'h2ca == r_count_14_io_out ? io_r_714_b : _GEN_11303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11305 = 10'h2cb == r_count_14_io_out ? io_r_715_b : _GEN_11304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11306 = 10'h2cc == r_count_14_io_out ? io_r_716_b : _GEN_11305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11307 = 10'h2cd == r_count_14_io_out ? io_r_717_b : _GEN_11306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11308 = 10'h2ce == r_count_14_io_out ? io_r_718_b : _GEN_11307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11309 = 10'h2cf == r_count_14_io_out ? io_r_719_b : _GEN_11308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11310 = 10'h2d0 == r_count_14_io_out ? io_r_720_b : _GEN_11309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11311 = 10'h2d1 == r_count_14_io_out ? io_r_721_b : _GEN_11310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11312 = 10'h2d2 == r_count_14_io_out ? io_r_722_b : _GEN_11311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11313 = 10'h2d3 == r_count_14_io_out ? io_r_723_b : _GEN_11312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11314 = 10'h2d4 == r_count_14_io_out ? io_r_724_b : _GEN_11313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11315 = 10'h2d5 == r_count_14_io_out ? io_r_725_b : _GEN_11314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11316 = 10'h2d6 == r_count_14_io_out ? io_r_726_b : _GEN_11315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11317 = 10'h2d7 == r_count_14_io_out ? io_r_727_b : _GEN_11316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11318 = 10'h2d8 == r_count_14_io_out ? io_r_728_b : _GEN_11317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11319 = 10'h2d9 == r_count_14_io_out ? io_r_729_b : _GEN_11318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11320 = 10'h2da == r_count_14_io_out ? io_r_730_b : _GEN_11319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11321 = 10'h2db == r_count_14_io_out ? io_r_731_b : _GEN_11320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11322 = 10'h2dc == r_count_14_io_out ? io_r_732_b : _GEN_11321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11323 = 10'h2dd == r_count_14_io_out ? io_r_733_b : _GEN_11322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11324 = 10'h2de == r_count_14_io_out ? io_r_734_b : _GEN_11323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11325 = 10'h2df == r_count_14_io_out ? io_r_735_b : _GEN_11324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11326 = 10'h2e0 == r_count_14_io_out ? io_r_736_b : _GEN_11325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11327 = 10'h2e1 == r_count_14_io_out ? io_r_737_b : _GEN_11326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11328 = 10'h2e2 == r_count_14_io_out ? io_r_738_b : _GEN_11327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11329 = 10'h2e3 == r_count_14_io_out ? io_r_739_b : _GEN_11328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11330 = 10'h2e4 == r_count_14_io_out ? io_r_740_b : _GEN_11329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11331 = 10'h2e5 == r_count_14_io_out ? io_r_741_b : _GEN_11330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11332 = 10'h2e6 == r_count_14_io_out ? io_r_742_b : _GEN_11331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11333 = 10'h2e7 == r_count_14_io_out ? io_r_743_b : _GEN_11332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11334 = 10'h2e8 == r_count_14_io_out ? io_r_744_b : _GEN_11333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11335 = 10'h2e9 == r_count_14_io_out ? io_r_745_b : _GEN_11334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11336 = 10'h2ea == r_count_14_io_out ? io_r_746_b : _GEN_11335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11337 = 10'h2eb == r_count_14_io_out ? io_r_747_b : _GEN_11336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11338 = 10'h2ec == r_count_14_io_out ? io_r_748_b : _GEN_11337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11341 = 10'h1 == r_count_15_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11342 = 10'h2 == r_count_15_io_out ? io_r_2_b : _GEN_11341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11343 = 10'h3 == r_count_15_io_out ? io_r_3_b : _GEN_11342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11344 = 10'h4 == r_count_15_io_out ? io_r_4_b : _GEN_11343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11345 = 10'h5 == r_count_15_io_out ? io_r_5_b : _GEN_11344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11346 = 10'h6 == r_count_15_io_out ? io_r_6_b : _GEN_11345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11347 = 10'h7 == r_count_15_io_out ? io_r_7_b : _GEN_11346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11348 = 10'h8 == r_count_15_io_out ? io_r_8_b : _GEN_11347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11349 = 10'h9 == r_count_15_io_out ? io_r_9_b : _GEN_11348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11350 = 10'ha == r_count_15_io_out ? io_r_10_b : _GEN_11349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11351 = 10'hb == r_count_15_io_out ? io_r_11_b : _GEN_11350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11352 = 10'hc == r_count_15_io_out ? io_r_12_b : _GEN_11351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11353 = 10'hd == r_count_15_io_out ? io_r_13_b : _GEN_11352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11354 = 10'he == r_count_15_io_out ? io_r_14_b : _GEN_11353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11355 = 10'hf == r_count_15_io_out ? io_r_15_b : _GEN_11354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11356 = 10'h10 == r_count_15_io_out ? io_r_16_b : _GEN_11355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11357 = 10'h11 == r_count_15_io_out ? io_r_17_b : _GEN_11356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11358 = 10'h12 == r_count_15_io_out ? io_r_18_b : _GEN_11357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11359 = 10'h13 == r_count_15_io_out ? io_r_19_b : _GEN_11358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11360 = 10'h14 == r_count_15_io_out ? io_r_20_b : _GEN_11359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11361 = 10'h15 == r_count_15_io_out ? io_r_21_b : _GEN_11360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11362 = 10'h16 == r_count_15_io_out ? io_r_22_b : _GEN_11361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11363 = 10'h17 == r_count_15_io_out ? io_r_23_b : _GEN_11362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11364 = 10'h18 == r_count_15_io_out ? io_r_24_b : _GEN_11363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11365 = 10'h19 == r_count_15_io_out ? io_r_25_b : _GEN_11364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11366 = 10'h1a == r_count_15_io_out ? io_r_26_b : _GEN_11365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11367 = 10'h1b == r_count_15_io_out ? io_r_27_b : _GEN_11366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11368 = 10'h1c == r_count_15_io_out ? io_r_28_b : _GEN_11367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11369 = 10'h1d == r_count_15_io_out ? io_r_29_b : _GEN_11368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11370 = 10'h1e == r_count_15_io_out ? io_r_30_b : _GEN_11369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11371 = 10'h1f == r_count_15_io_out ? io_r_31_b : _GEN_11370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11372 = 10'h20 == r_count_15_io_out ? io_r_32_b : _GEN_11371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11373 = 10'h21 == r_count_15_io_out ? io_r_33_b : _GEN_11372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11374 = 10'h22 == r_count_15_io_out ? io_r_34_b : _GEN_11373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11375 = 10'h23 == r_count_15_io_out ? io_r_35_b : _GEN_11374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11376 = 10'h24 == r_count_15_io_out ? io_r_36_b : _GEN_11375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11377 = 10'h25 == r_count_15_io_out ? io_r_37_b : _GEN_11376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11378 = 10'h26 == r_count_15_io_out ? io_r_38_b : _GEN_11377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11379 = 10'h27 == r_count_15_io_out ? io_r_39_b : _GEN_11378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11380 = 10'h28 == r_count_15_io_out ? io_r_40_b : _GEN_11379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11381 = 10'h29 == r_count_15_io_out ? io_r_41_b : _GEN_11380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11382 = 10'h2a == r_count_15_io_out ? io_r_42_b : _GEN_11381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11383 = 10'h2b == r_count_15_io_out ? io_r_43_b : _GEN_11382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11384 = 10'h2c == r_count_15_io_out ? io_r_44_b : _GEN_11383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11385 = 10'h2d == r_count_15_io_out ? io_r_45_b : _GEN_11384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11386 = 10'h2e == r_count_15_io_out ? io_r_46_b : _GEN_11385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11387 = 10'h2f == r_count_15_io_out ? io_r_47_b : _GEN_11386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11388 = 10'h30 == r_count_15_io_out ? io_r_48_b : _GEN_11387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11389 = 10'h31 == r_count_15_io_out ? io_r_49_b : _GEN_11388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11390 = 10'h32 == r_count_15_io_out ? io_r_50_b : _GEN_11389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11391 = 10'h33 == r_count_15_io_out ? io_r_51_b : _GEN_11390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11392 = 10'h34 == r_count_15_io_out ? io_r_52_b : _GEN_11391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11393 = 10'h35 == r_count_15_io_out ? io_r_53_b : _GEN_11392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11394 = 10'h36 == r_count_15_io_out ? io_r_54_b : _GEN_11393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11395 = 10'h37 == r_count_15_io_out ? io_r_55_b : _GEN_11394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11396 = 10'h38 == r_count_15_io_out ? io_r_56_b : _GEN_11395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11397 = 10'h39 == r_count_15_io_out ? io_r_57_b : _GEN_11396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11398 = 10'h3a == r_count_15_io_out ? io_r_58_b : _GEN_11397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11399 = 10'h3b == r_count_15_io_out ? io_r_59_b : _GEN_11398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11400 = 10'h3c == r_count_15_io_out ? io_r_60_b : _GEN_11399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11401 = 10'h3d == r_count_15_io_out ? io_r_61_b : _GEN_11400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11402 = 10'h3e == r_count_15_io_out ? io_r_62_b : _GEN_11401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11403 = 10'h3f == r_count_15_io_out ? io_r_63_b : _GEN_11402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11404 = 10'h40 == r_count_15_io_out ? io_r_64_b : _GEN_11403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11405 = 10'h41 == r_count_15_io_out ? io_r_65_b : _GEN_11404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11406 = 10'h42 == r_count_15_io_out ? io_r_66_b : _GEN_11405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11407 = 10'h43 == r_count_15_io_out ? io_r_67_b : _GEN_11406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11408 = 10'h44 == r_count_15_io_out ? io_r_68_b : _GEN_11407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11409 = 10'h45 == r_count_15_io_out ? io_r_69_b : _GEN_11408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11410 = 10'h46 == r_count_15_io_out ? io_r_70_b : _GEN_11409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11411 = 10'h47 == r_count_15_io_out ? io_r_71_b : _GEN_11410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11412 = 10'h48 == r_count_15_io_out ? io_r_72_b : _GEN_11411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11413 = 10'h49 == r_count_15_io_out ? io_r_73_b : _GEN_11412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11414 = 10'h4a == r_count_15_io_out ? io_r_74_b : _GEN_11413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11415 = 10'h4b == r_count_15_io_out ? io_r_75_b : _GEN_11414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11416 = 10'h4c == r_count_15_io_out ? io_r_76_b : _GEN_11415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11417 = 10'h4d == r_count_15_io_out ? io_r_77_b : _GEN_11416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11418 = 10'h4e == r_count_15_io_out ? io_r_78_b : _GEN_11417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11419 = 10'h4f == r_count_15_io_out ? io_r_79_b : _GEN_11418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11420 = 10'h50 == r_count_15_io_out ? io_r_80_b : _GEN_11419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11421 = 10'h51 == r_count_15_io_out ? io_r_81_b : _GEN_11420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11422 = 10'h52 == r_count_15_io_out ? io_r_82_b : _GEN_11421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11423 = 10'h53 == r_count_15_io_out ? io_r_83_b : _GEN_11422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11424 = 10'h54 == r_count_15_io_out ? io_r_84_b : _GEN_11423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11425 = 10'h55 == r_count_15_io_out ? io_r_85_b : _GEN_11424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11426 = 10'h56 == r_count_15_io_out ? io_r_86_b : _GEN_11425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11427 = 10'h57 == r_count_15_io_out ? io_r_87_b : _GEN_11426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11428 = 10'h58 == r_count_15_io_out ? io_r_88_b : _GEN_11427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11429 = 10'h59 == r_count_15_io_out ? io_r_89_b : _GEN_11428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11430 = 10'h5a == r_count_15_io_out ? io_r_90_b : _GEN_11429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11431 = 10'h5b == r_count_15_io_out ? io_r_91_b : _GEN_11430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11432 = 10'h5c == r_count_15_io_out ? io_r_92_b : _GEN_11431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11433 = 10'h5d == r_count_15_io_out ? io_r_93_b : _GEN_11432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11434 = 10'h5e == r_count_15_io_out ? io_r_94_b : _GEN_11433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11435 = 10'h5f == r_count_15_io_out ? io_r_95_b : _GEN_11434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11436 = 10'h60 == r_count_15_io_out ? io_r_96_b : _GEN_11435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11437 = 10'h61 == r_count_15_io_out ? io_r_97_b : _GEN_11436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11438 = 10'h62 == r_count_15_io_out ? io_r_98_b : _GEN_11437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11439 = 10'h63 == r_count_15_io_out ? io_r_99_b : _GEN_11438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11440 = 10'h64 == r_count_15_io_out ? io_r_100_b : _GEN_11439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11441 = 10'h65 == r_count_15_io_out ? io_r_101_b : _GEN_11440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11442 = 10'h66 == r_count_15_io_out ? io_r_102_b : _GEN_11441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11443 = 10'h67 == r_count_15_io_out ? io_r_103_b : _GEN_11442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11444 = 10'h68 == r_count_15_io_out ? io_r_104_b : _GEN_11443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11445 = 10'h69 == r_count_15_io_out ? io_r_105_b : _GEN_11444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11446 = 10'h6a == r_count_15_io_out ? io_r_106_b : _GEN_11445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11447 = 10'h6b == r_count_15_io_out ? io_r_107_b : _GEN_11446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11448 = 10'h6c == r_count_15_io_out ? io_r_108_b : _GEN_11447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11449 = 10'h6d == r_count_15_io_out ? io_r_109_b : _GEN_11448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11450 = 10'h6e == r_count_15_io_out ? io_r_110_b : _GEN_11449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11451 = 10'h6f == r_count_15_io_out ? io_r_111_b : _GEN_11450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11452 = 10'h70 == r_count_15_io_out ? io_r_112_b : _GEN_11451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11453 = 10'h71 == r_count_15_io_out ? io_r_113_b : _GEN_11452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11454 = 10'h72 == r_count_15_io_out ? io_r_114_b : _GEN_11453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11455 = 10'h73 == r_count_15_io_out ? io_r_115_b : _GEN_11454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11456 = 10'h74 == r_count_15_io_out ? io_r_116_b : _GEN_11455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11457 = 10'h75 == r_count_15_io_out ? io_r_117_b : _GEN_11456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11458 = 10'h76 == r_count_15_io_out ? io_r_118_b : _GEN_11457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11459 = 10'h77 == r_count_15_io_out ? io_r_119_b : _GEN_11458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11460 = 10'h78 == r_count_15_io_out ? io_r_120_b : _GEN_11459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11461 = 10'h79 == r_count_15_io_out ? io_r_121_b : _GEN_11460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11462 = 10'h7a == r_count_15_io_out ? io_r_122_b : _GEN_11461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11463 = 10'h7b == r_count_15_io_out ? io_r_123_b : _GEN_11462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11464 = 10'h7c == r_count_15_io_out ? io_r_124_b : _GEN_11463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11465 = 10'h7d == r_count_15_io_out ? io_r_125_b : _GEN_11464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11466 = 10'h7e == r_count_15_io_out ? io_r_126_b : _GEN_11465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11467 = 10'h7f == r_count_15_io_out ? io_r_127_b : _GEN_11466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11468 = 10'h80 == r_count_15_io_out ? io_r_128_b : _GEN_11467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11469 = 10'h81 == r_count_15_io_out ? io_r_129_b : _GEN_11468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11470 = 10'h82 == r_count_15_io_out ? io_r_130_b : _GEN_11469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11471 = 10'h83 == r_count_15_io_out ? io_r_131_b : _GEN_11470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11472 = 10'h84 == r_count_15_io_out ? io_r_132_b : _GEN_11471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11473 = 10'h85 == r_count_15_io_out ? io_r_133_b : _GEN_11472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11474 = 10'h86 == r_count_15_io_out ? io_r_134_b : _GEN_11473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11475 = 10'h87 == r_count_15_io_out ? io_r_135_b : _GEN_11474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11476 = 10'h88 == r_count_15_io_out ? io_r_136_b : _GEN_11475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11477 = 10'h89 == r_count_15_io_out ? io_r_137_b : _GEN_11476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11478 = 10'h8a == r_count_15_io_out ? io_r_138_b : _GEN_11477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11479 = 10'h8b == r_count_15_io_out ? io_r_139_b : _GEN_11478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11480 = 10'h8c == r_count_15_io_out ? io_r_140_b : _GEN_11479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11481 = 10'h8d == r_count_15_io_out ? io_r_141_b : _GEN_11480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11482 = 10'h8e == r_count_15_io_out ? io_r_142_b : _GEN_11481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11483 = 10'h8f == r_count_15_io_out ? io_r_143_b : _GEN_11482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11484 = 10'h90 == r_count_15_io_out ? io_r_144_b : _GEN_11483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11485 = 10'h91 == r_count_15_io_out ? io_r_145_b : _GEN_11484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11486 = 10'h92 == r_count_15_io_out ? io_r_146_b : _GEN_11485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11487 = 10'h93 == r_count_15_io_out ? io_r_147_b : _GEN_11486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11488 = 10'h94 == r_count_15_io_out ? io_r_148_b : _GEN_11487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11489 = 10'h95 == r_count_15_io_out ? io_r_149_b : _GEN_11488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11490 = 10'h96 == r_count_15_io_out ? io_r_150_b : _GEN_11489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11491 = 10'h97 == r_count_15_io_out ? io_r_151_b : _GEN_11490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11492 = 10'h98 == r_count_15_io_out ? io_r_152_b : _GEN_11491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11493 = 10'h99 == r_count_15_io_out ? io_r_153_b : _GEN_11492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11494 = 10'h9a == r_count_15_io_out ? io_r_154_b : _GEN_11493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11495 = 10'h9b == r_count_15_io_out ? io_r_155_b : _GEN_11494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11496 = 10'h9c == r_count_15_io_out ? io_r_156_b : _GEN_11495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11497 = 10'h9d == r_count_15_io_out ? io_r_157_b : _GEN_11496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11498 = 10'h9e == r_count_15_io_out ? io_r_158_b : _GEN_11497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11499 = 10'h9f == r_count_15_io_out ? io_r_159_b : _GEN_11498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11500 = 10'ha0 == r_count_15_io_out ? io_r_160_b : _GEN_11499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11501 = 10'ha1 == r_count_15_io_out ? io_r_161_b : _GEN_11500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11502 = 10'ha2 == r_count_15_io_out ? io_r_162_b : _GEN_11501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11503 = 10'ha3 == r_count_15_io_out ? io_r_163_b : _GEN_11502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11504 = 10'ha4 == r_count_15_io_out ? io_r_164_b : _GEN_11503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11505 = 10'ha5 == r_count_15_io_out ? io_r_165_b : _GEN_11504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11506 = 10'ha6 == r_count_15_io_out ? io_r_166_b : _GEN_11505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11507 = 10'ha7 == r_count_15_io_out ? io_r_167_b : _GEN_11506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11508 = 10'ha8 == r_count_15_io_out ? io_r_168_b : _GEN_11507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11509 = 10'ha9 == r_count_15_io_out ? io_r_169_b : _GEN_11508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11510 = 10'haa == r_count_15_io_out ? io_r_170_b : _GEN_11509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11511 = 10'hab == r_count_15_io_out ? io_r_171_b : _GEN_11510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11512 = 10'hac == r_count_15_io_out ? io_r_172_b : _GEN_11511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11513 = 10'had == r_count_15_io_out ? io_r_173_b : _GEN_11512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11514 = 10'hae == r_count_15_io_out ? io_r_174_b : _GEN_11513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11515 = 10'haf == r_count_15_io_out ? io_r_175_b : _GEN_11514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11516 = 10'hb0 == r_count_15_io_out ? io_r_176_b : _GEN_11515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11517 = 10'hb1 == r_count_15_io_out ? io_r_177_b : _GEN_11516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11518 = 10'hb2 == r_count_15_io_out ? io_r_178_b : _GEN_11517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11519 = 10'hb3 == r_count_15_io_out ? io_r_179_b : _GEN_11518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11520 = 10'hb4 == r_count_15_io_out ? io_r_180_b : _GEN_11519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11521 = 10'hb5 == r_count_15_io_out ? io_r_181_b : _GEN_11520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11522 = 10'hb6 == r_count_15_io_out ? io_r_182_b : _GEN_11521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11523 = 10'hb7 == r_count_15_io_out ? io_r_183_b : _GEN_11522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11524 = 10'hb8 == r_count_15_io_out ? io_r_184_b : _GEN_11523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11525 = 10'hb9 == r_count_15_io_out ? io_r_185_b : _GEN_11524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11526 = 10'hba == r_count_15_io_out ? io_r_186_b : _GEN_11525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11527 = 10'hbb == r_count_15_io_out ? io_r_187_b : _GEN_11526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11528 = 10'hbc == r_count_15_io_out ? io_r_188_b : _GEN_11527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11529 = 10'hbd == r_count_15_io_out ? io_r_189_b : _GEN_11528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11530 = 10'hbe == r_count_15_io_out ? io_r_190_b : _GEN_11529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11531 = 10'hbf == r_count_15_io_out ? io_r_191_b : _GEN_11530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11532 = 10'hc0 == r_count_15_io_out ? io_r_192_b : _GEN_11531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11533 = 10'hc1 == r_count_15_io_out ? io_r_193_b : _GEN_11532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11534 = 10'hc2 == r_count_15_io_out ? io_r_194_b : _GEN_11533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11535 = 10'hc3 == r_count_15_io_out ? io_r_195_b : _GEN_11534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11536 = 10'hc4 == r_count_15_io_out ? io_r_196_b : _GEN_11535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11537 = 10'hc5 == r_count_15_io_out ? io_r_197_b : _GEN_11536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11538 = 10'hc6 == r_count_15_io_out ? io_r_198_b : _GEN_11537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11539 = 10'hc7 == r_count_15_io_out ? io_r_199_b : _GEN_11538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11540 = 10'hc8 == r_count_15_io_out ? io_r_200_b : _GEN_11539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11541 = 10'hc9 == r_count_15_io_out ? io_r_201_b : _GEN_11540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11542 = 10'hca == r_count_15_io_out ? io_r_202_b : _GEN_11541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11543 = 10'hcb == r_count_15_io_out ? io_r_203_b : _GEN_11542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11544 = 10'hcc == r_count_15_io_out ? io_r_204_b : _GEN_11543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11545 = 10'hcd == r_count_15_io_out ? io_r_205_b : _GEN_11544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11546 = 10'hce == r_count_15_io_out ? io_r_206_b : _GEN_11545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11547 = 10'hcf == r_count_15_io_out ? io_r_207_b : _GEN_11546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11548 = 10'hd0 == r_count_15_io_out ? io_r_208_b : _GEN_11547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11549 = 10'hd1 == r_count_15_io_out ? io_r_209_b : _GEN_11548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11550 = 10'hd2 == r_count_15_io_out ? io_r_210_b : _GEN_11549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11551 = 10'hd3 == r_count_15_io_out ? io_r_211_b : _GEN_11550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11552 = 10'hd4 == r_count_15_io_out ? io_r_212_b : _GEN_11551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11553 = 10'hd5 == r_count_15_io_out ? io_r_213_b : _GEN_11552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11554 = 10'hd6 == r_count_15_io_out ? io_r_214_b : _GEN_11553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11555 = 10'hd7 == r_count_15_io_out ? io_r_215_b : _GEN_11554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11556 = 10'hd8 == r_count_15_io_out ? io_r_216_b : _GEN_11555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11557 = 10'hd9 == r_count_15_io_out ? io_r_217_b : _GEN_11556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11558 = 10'hda == r_count_15_io_out ? io_r_218_b : _GEN_11557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11559 = 10'hdb == r_count_15_io_out ? io_r_219_b : _GEN_11558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11560 = 10'hdc == r_count_15_io_out ? io_r_220_b : _GEN_11559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11561 = 10'hdd == r_count_15_io_out ? io_r_221_b : _GEN_11560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11562 = 10'hde == r_count_15_io_out ? io_r_222_b : _GEN_11561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11563 = 10'hdf == r_count_15_io_out ? io_r_223_b : _GEN_11562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11564 = 10'he0 == r_count_15_io_out ? io_r_224_b : _GEN_11563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11565 = 10'he1 == r_count_15_io_out ? io_r_225_b : _GEN_11564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11566 = 10'he2 == r_count_15_io_out ? io_r_226_b : _GEN_11565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11567 = 10'he3 == r_count_15_io_out ? io_r_227_b : _GEN_11566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11568 = 10'he4 == r_count_15_io_out ? io_r_228_b : _GEN_11567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11569 = 10'he5 == r_count_15_io_out ? io_r_229_b : _GEN_11568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11570 = 10'he6 == r_count_15_io_out ? io_r_230_b : _GEN_11569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11571 = 10'he7 == r_count_15_io_out ? io_r_231_b : _GEN_11570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11572 = 10'he8 == r_count_15_io_out ? io_r_232_b : _GEN_11571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11573 = 10'he9 == r_count_15_io_out ? io_r_233_b : _GEN_11572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11574 = 10'hea == r_count_15_io_out ? io_r_234_b : _GEN_11573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11575 = 10'heb == r_count_15_io_out ? io_r_235_b : _GEN_11574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11576 = 10'hec == r_count_15_io_out ? io_r_236_b : _GEN_11575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11577 = 10'hed == r_count_15_io_out ? io_r_237_b : _GEN_11576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11578 = 10'hee == r_count_15_io_out ? io_r_238_b : _GEN_11577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11579 = 10'hef == r_count_15_io_out ? io_r_239_b : _GEN_11578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11580 = 10'hf0 == r_count_15_io_out ? io_r_240_b : _GEN_11579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11581 = 10'hf1 == r_count_15_io_out ? io_r_241_b : _GEN_11580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11582 = 10'hf2 == r_count_15_io_out ? io_r_242_b : _GEN_11581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11583 = 10'hf3 == r_count_15_io_out ? io_r_243_b : _GEN_11582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11584 = 10'hf4 == r_count_15_io_out ? io_r_244_b : _GEN_11583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11585 = 10'hf5 == r_count_15_io_out ? io_r_245_b : _GEN_11584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11586 = 10'hf6 == r_count_15_io_out ? io_r_246_b : _GEN_11585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11587 = 10'hf7 == r_count_15_io_out ? io_r_247_b : _GEN_11586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11588 = 10'hf8 == r_count_15_io_out ? io_r_248_b : _GEN_11587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11589 = 10'hf9 == r_count_15_io_out ? io_r_249_b : _GEN_11588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11590 = 10'hfa == r_count_15_io_out ? io_r_250_b : _GEN_11589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11591 = 10'hfb == r_count_15_io_out ? io_r_251_b : _GEN_11590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11592 = 10'hfc == r_count_15_io_out ? io_r_252_b : _GEN_11591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11593 = 10'hfd == r_count_15_io_out ? io_r_253_b : _GEN_11592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11594 = 10'hfe == r_count_15_io_out ? io_r_254_b : _GEN_11593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11595 = 10'hff == r_count_15_io_out ? io_r_255_b : _GEN_11594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11596 = 10'h100 == r_count_15_io_out ? io_r_256_b : _GEN_11595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11597 = 10'h101 == r_count_15_io_out ? io_r_257_b : _GEN_11596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11598 = 10'h102 == r_count_15_io_out ? io_r_258_b : _GEN_11597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11599 = 10'h103 == r_count_15_io_out ? io_r_259_b : _GEN_11598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11600 = 10'h104 == r_count_15_io_out ? io_r_260_b : _GEN_11599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11601 = 10'h105 == r_count_15_io_out ? io_r_261_b : _GEN_11600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11602 = 10'h106 == r_count_15_io_out ? io_r_262_b : _GEN_11601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11603 = 10'h107 == r_count_15_io_out ? io_r_263_b : _GEN_11602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11604 = 10'h108 == r_count_15_io_out ? io_r_264_b : _GEN_11603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11605 = 10'h109 == r_count_15_io_out ? io_r_265_b : _GEN_11604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11606 = 10'h10a == r_count_15_io_out ? io_r_266_b : _GEN_11605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11607 = 10'h10b == r_count_15_io_out ? io_r_267_b : _GEN_11606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11608 = 10'h10c == r_count_15_io_out ? io_r_268_b : _GEN_11607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11609 = 10'h10d == r_count_15_io_out ? io_r_269_b : _GEN_11608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11610 = 10'h10e == r_count_15_io_out ? io_r_270_b : _GEN_11609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11611 = 10'h10f == r_count_15_io_out ? io_r_271_b : _GEN_11610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11612 = 10'h110 == r_count_15_io_out ? io_r_272_b : _GEN_11611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11613 = 10'h111 == r_count_15_io_out ? io_r_273_b : _GEN_11612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11614 = 10'h112 == r_count_15_io_out ? io_r_274_b : _GEN_11613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11615 = 10'h113 == r_count_15_io_out ? io_r_275_b : _GEN_11614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11616 = 10'h114 == r_count_15_io_out ? io_r_276_b : _GEN_11615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11617 = 10'h115 == r_count_15_io_out ? io_r_277_b : _GEN_11616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11618 = 10'h116 == r_count_15_io_out ? io_r_278_b : _GEN_11617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11619 = 10'h117 == r_count_15_io_out ? io_r_279_b : _GEN_11618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11620 = 10'h118 == r_count_15_io_out ? io_r_280_b : _GEN_11619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11621 = 10'h119 == r_count_15_io_out ? io_r_281_b : _GEN_11620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11622 = 10'h11a == r_count_15_io_out ? io_r_282_b : _GEN_11621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11623 = 10'h11b == r_count_15_io_out ? io_r_283_b : _GEN_11622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11624 = 10'h11c == r_count_15_io_out ? io_r_284_b : _GEN_11623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11625 = 10'h11d == r_count_15_io_out ? io_r_285_b : _GEN_11624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11626 = 10'h11e == r_count_15_io_out ? io_r_286_b : _GEN_11625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11627 = 10'h11f == r_count_15_io_out ? io_r_287_b : _GEN_11626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11628 = 10'h120 == r_count_15_io_out ? io_r_288_b : _GEN_11627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11629 = 10'h121 == r_count_15_io_out ? io_r_289_b : _GEN_11628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11630 = 10'h122 == r_count_15_io_out ? io_r_290_b : _GEN_11629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11631 = 10'h123 == r_count_15_io_out ? io_r_291_b : _GEN_11630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11632 = 10'h124 == r_count_15_io_out ? io_r_292_b : _GEN_11631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11633 = 10'h125 == r_count_15_io_out ? io_r_293_b : _GEN_11632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11634 = 10'h126 == r_count_15_io_out ? io_r_294_b : _GEN_11633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11635 = 10'h127 == r_count_15_io_out ? io_r_295_b : _GEN_11634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11636 = 10'h128 == r_count_15_io_out ? io_r_296_b : _GEN_11635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11637 = 10'h129 == r_count_15_io_out ? io_r_297_b : _GEN_11636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11638 = 10'h12a == r_count_15_io_out ? io_r_298_b : _GEN_11637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11639 = 10'h12b == r_count_15_io_out ? io_r_299_b : _GEN_11638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11640 = 10'h12c == r_count_15_io_out ? io_r_300_b : _GEN_11639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11641 = 10'h12d == r_count_15_io_out ? io_r_301_b : _GEN_11640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11642 = 10'h12e == r_count_15_io_out ? io_r_302_b : _GEN_11641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11643 = 10'h12f == r_count_15_io_out ? io_r_303_b : _GEN_11642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11644 = 10'h130 == r_count_15_io_out ? io_r_304_b : _GEN_11643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11645 = 10'h131 == r_count_15_io_out ? io_r_305_b : _GEN_11644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11646 = 10'h132 == r_count_15_io_out ? io_r_306_b : _GEN_11645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11647 = 10'h133 == r_count_15_io_out ? io_r_307_b : _GEN_11646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11648 = 10'h134 == r_count_15_io_out ? io_r_308_b : _GEN_11647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11649 = 10'h135 == r_count_15_io_out ? io_r_309_b : _GEN_11648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11650 = 10'h136 == r_count_15_io_out ? io_r_310_b : _GEN_11649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11651 = 10'h137 == r_count_15_io_out ? io_r_311_b : _GEN_11650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11652 = 10'h138 == r_count_15_io_out ? io_r_312_b : _GEN_11651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11653 = 10'h139 == r_count_15_io_out ? io_r_313_b : _GEN_11652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11654 = 10'h13a == r_count_15_io_out ? io_r_314_b : _GEN_11653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11655 = 10'h13b == r_count_15_io_out ? io_r_315_b : _GEN_11654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11656 = 10'h13c == r_count_15_io_out ? io_r_316_b : _GEN_11655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11657 = 10'h13d == r_count_15_io_out ? io_r_317_b : _GEN_11656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11658 = 10'h13e == r_count_15_io_out ? io_r_318_b : _GEN_11657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11659 = 10'h13f == r_count_15_io_out ? io_r_319_b : _GEN_11658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11660 = 10'h140 == r_count_15_io_out ? io_r_320_b : _GEN_11659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11661 = 10'h141 == r_count_15_io_out ? io_r_321_b : _GEN_11660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11662 = 10'h142 == r_count_15_io_out ? io_r_322_b : _GEN_11661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11663 = 10'h143 == r_count_15_io_out ? io_r_323_b : _GEN_11662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11664 = 10'h144 == r_count_15_io_out ? io_r_324_b : _GEN_11663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11665 = 10'h145 == r_count_15_io_out ? io_r_325_b : _GEN_11664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11666 = 10'h146 == r_count_15_io_out ? io_r_326_b : _GEN_11665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11667 = 10'h147 == r_count_15_io_out ? io_r_327_b : _GEN_11666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11668 = 10'h148 == r_count_15_io_out ? io_r_328_b : _GEN_11667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11669 = 10'h149 == r_count_15_io_out ? io_r_329_b : _GEN_11668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11670 = 10'h14a == r_count_15_io_out ? io_r_330_b : _GEN_11669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11671 = 10'h14b == r_count_15_io_out ? io_r_331_b : _GEN_11670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11672 = 10'h14c == r_count_15_io_out ? io_r_332_b : _GEN_11671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11673 = 10'h14d == r_count_15_io_out ? io_r_333_b : _GEN_11672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11674 = 10'h14e == r_count_15_io_out ? io_r_334_b : _GEN_11673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11675 = 10'h14f == r_count_15_io_out ? io_r_335_b : _GEN_11674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11676 = 10'h150 == r_count_15_io_out ? io_r_336_b : _GEN_11675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11677 = 10'h151 == r_count_15_io_out ? io_r_337_b : _GEN_11676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11678 = 10'h152 == r_count_15_io_out ? io_r_338_b : _GEN_11677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11679 = 10'h153 == r_count_15_io_out ? io_r_339_b : _GEN_11678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11680 = 10'h154 == r_count_15_io_out ? io_r_340_b : _GEN_11679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11681 = 10'h155 == r_count_15_io_out ? io_r_341_b : _GEN_11680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11682 = 10'h156 == r_count_15_io_out ? io_r_342_b : _GEN_11681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11683 = 10'h157 == r_count_15_io_out ? io_r_343_b : _GEN_11682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11684 = 10'h158 == r_count_15_io_out ? io_r_344_b : _GEN_11683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11685 = 10'h159 == r_count_15_io_out ? io_r_345_b : _GEN_11684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11686 = 10'h15a == r_count_15_io_out ? io_r_346_b : _GEN_11685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11687 = 10'h15b == r_count_15_io_out ? io_r_347_b : _GEN_11686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11688 = 10'h15c == r_count_15_io_out ? io_r_348_b : _GEN_11687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11689 = 10'h15d == r_count_15_io_out ? io_r_349_b : _GEN_11688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11690 = 10'h15e == r_count_15_io_out ? io_r_350_b : _GEN_11689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11691 = 10'h15f == r_count_15_io_out ? io_r_351_b : _GEN_11690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11692 = 10'h160 == r_count_15_io_out ? io_r_352_b : _GEN_11691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11693 = 10'h161 == r_count_15_io_out ? io_r_353_b : _GEN_11692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11694 = 10'h162 == r_count_15_io_out ? io_r_354_b : _GEN_11693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11695 = 10'h163 == r_count_15_io_out ? io_r_355_b : _GEN_11694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11696 = 10'h164 == r_count_15_io_out ? io_r_356_b : _GEN_11695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11697 = 10'h165 == r_count_15_io_out ? io_r_357_b : _GEN_11696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11698 = 10'h166 == r_count_15_io_out ? io_r_358_b : _GEN_11697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11699 = 10'h167 == r_count_15_io_out ? io_r_359_b : _GEN_11698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11700 = 10'h168 == r_count_15_io_out ? io_r_360_b : _GEN_11699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11701 = 10'h169 == r_count_15_io_out ? io_r_361_b : _GEN_11700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11702 = 10'h16a == r_count_15_io_out ? io_r_362_b : _GEN_11701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11703 = 10'h16b == r_count_15_io_out ? io_r_363_b : _GEN_11702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11704 = 10'h16c == r_count_15_io_out ? io_r_364_b : _GEN_11703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11705 = 10'h16d == r_count_15_io_out ? io_r_365_b : _GEN_11704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11706 = 10'h16e == r_count_15_io_out ? io_r_366_b : _GEN_11705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11707 = 10'h16f == r_count_15_io_out ? io_r_367_b : _GEN_11706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11708 = 10'h170 == r_count_15_io_out ? io_r_368_b : _GEN_11707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11709 = 10'h171 == r_count_15_io_out ? io_r_369_b : _GEN_11708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11710 = 10'h172 == r_count_15_io_out ? io_r_370_b : _GEN_11709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11711 = 10'h173 == r_count_15_io_out ? io_r_371_b : _GEN_11710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11712 = 10'h174 == r_count_15_io_out ? io_r_372_b : _GEN_11711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11713 = 10'h175 == r_count_15_io_out ? io_r_373_b : _GEN_11712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11714 = 10'h176 == r_count_15_io_out ? io_r_374_b : _GEN_11713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11715 = 10'h177 == r_count_15_io_out ? io_r_375_b : _GEN_11714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11716 = 10'h178 == r_count_15_io_out ? io_r_376_b : _GEN_11715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11717 = 10'h179 == r_count_15_io_out ? io_r_377_b : _GEN_11716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11718 = 10'h17a == r_count_15_io_out ? io_r_378_b : _GEN_11717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11719 = 10'h17b == r_count_15_io_out ? io_r_379_b : _GEN_11718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11720 = 10'h17c == r_count_15_io_out ? io_r_380_b : _GEN_11719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11721 = 10'h17d == r_count_15_io_out ? io_r_381_b : _GEN_11720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11722 = 10'h17e == r_count_15_io_out ? io_r_382_b : _GEN_11721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11723 = 10'h17f == r_count_15_io_out ? io_r_383_b : _GEN_11722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11724 = 10'h180 == r_count_15_io_out ? io_r_384_b : _GEN_11723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11725 = 10'h181 == r_count_15_io_out ? io_r_385_b : _GEN_11724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11726 = 10'h182 == r_count_15_io_out ? io_r_386_b : _GEN_11725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11727 = 10'h183 == r_count_15_io_out ? io_r_387_b : _GEN_11726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11728 = 10'h184 == r_count_15_io_out ? io_r_388_b : _GEN_11727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11729 = 10'h185 == r_count_15_io_out ? io_r_389_b : _GEN_11728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11730 = 10'h186 == r_count_15_io_out ? io_r_390_b : _GEN_11729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11731 = 10'h187 == r_count_15_io_out ? io_r_391_b : _GEN_11730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11732 = 10'h188 == r_count_15_io_out ? io_r_392_b : _GEN_11731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11733 = 10'h189 == r_count_15_io_out ? io_r_393_b : _GEN_11732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11734 = 10'h18a == r_count_15_io_out ? io_r_394_b : _GEN_11733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11735 = 10'h18b == r_count_15_io_out ? io_r_395_b : _GEN_11734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11736 = 10'h18c == r_count_15_io_out ? io_r_396_b : _GEN_11735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11737 = 10'h18d == r_count_15_io_out ? io_r_397_b : _GEN_11736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11738 = 10'h18e == r_count_15_io_out ? io_r_398_b : _GEN_11737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11739 = 10'h18f == r_count_15_io_out ? io_r_399_b : _GEN_11738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11740 = 10'h190 == r_count_15_io_out ? io_r_400_b : _GEN_11739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11741 = 10'h191 == r_count_15_io_out ? io_r_401_b : _GEN_11740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11742 = 10'h192 == r_count_15_io_out ? io_r_402_b : _GEN_11741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11743 = 10'h193 == r_count_15_io_out ? io_r_403_b : _GEN_11742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11744 = 10'h194 == r_count_15_io_out ? io_r_404_b : _GEN_11743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11745 = 10'h195 == r_count_15_io_out ? io_r_405_b : _GEN_11744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11746 = 10'h196 == r_count_15_io_out ? io_r_406_b : _GEN_11745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11747 = 10'h197 == r_count_15_io_out ? io_r_407_b : _GEN_11746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11748 = 10'h198 == r_count_15_io_out ? io_r_408_b : _GEN_11747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11749 = 10'h199 == r_count_15_io_out ? io_r_409_b : _GEN_11748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11750 = 10'h19a == r_count_15_io_out ? io_r_410_b : _GEN_11749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11751 = 10'h19b == r_count_15_io_out ? io_r_411_b : _GEN_11750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11752 = 10'h19c == r_count_15_io_out ? io_r_412_b : _GEN_11751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11753 = 10'h19d == r_count_15_io_out ? io_r_413_b : _GEN_11752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11754 = 10'h19e == r_count_15_io_out ? io_r_414_b : _GEN_11753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11755 = 10'h19f == r_count_15_io_out ? io_r_415_b : _GEN_11754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11756 = 10'h1a0 == r_count_15_io_out ? io_r_416_b : _GEN_11755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11757 = 10'h1a1 == r_count_15_io_out ? io_r_417_b : _GEN_11756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11758 = 10'h1a2 == r_count_15_io_out ? io_r_418_b : _GEN_11757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11759 = 10'h1a3 == r_count_15_io_out ? io_r_419_b : _GEN_11758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11760 = 10'h1a4 == r_count_15_io_out ? io_r_420_b : _GEN_11759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11761 = 10'h1a5 == r_count_15_io_out ? io_r_421_b : _GEN_11760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11762 = 10'h1a6 == r_count_15_io_out ? io_r_422_b : _GEN_11761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11763 = 10'h1a7 == r_count_15_io_out ? io_r_423_b : _GEN_11762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11764 = 10'h1a8 == r_count_15_io_out ? io_r_424_b : _GEN_11763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11765 = 10'h1a9 == r_count_15_io_out ? io_r_425_b : _GEN_11764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11766 = 10'h1aa == r_count_15_io_out ? io_r_426_b : _GEN_11765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11767 = 10'h1ab == r_count_15_io_out ? io_r_427_b : _GEN_11766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11768 = 10'h1ac == r_count_15_io_out ? io_r_428_b : _GEN_11767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11769 = 10'h1ad == r_count_15_io_out ? io_r_429_b : _GEN_11768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11770 = 10'h1ae == r_count_15_io_out ? io_r_430_b : _GEN_11769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11771 = 10'h1af == r_count_15_io_out ? io_r_431_b : _GEN_11770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11772 = 10'h1b0 == r_count_15_io_out ? io_r_432_b : _GEN_11771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11773 = 10'h1b1 == r_count_15_io_out ? io_r_433_b : _GEN_11772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11774 = 10'h1b2 == r_count_15_io_out ? io_r_434_b : _GEN_11773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11775 = 10'h1b3 == r_count_15_io_out ? io_r_435_b : _GEN_11774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11776 = 10'h1b4 == r_count_15_io_out ? io_r_436_b : _GEN_11775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11777 = 10'h1b5 == r_count_15_io_out ? io_r_437_b : _GEN_11776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11778 = 10'h1b6 == r_count_15_io_out ? io_r_438_b : _GEN_11777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11779 = 10'h1b7 == r_count_15_io_out ? io_r_439_b : _GEN_11778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11780 = 10'h1b8 == r_count_15_io_out ? io_r_440_b : _GEN_11779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11781 = 10'h1b9 == r_count_15_io_out ? io_r_441_b : _GEN_11780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11782 = 10'h1ba == r_count_15_io_out ? io_r_442_b : _GEN_11781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11783 = 10'h1bb == r_count_15_io_out ? io_r_443_b : _GEN_11782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11784 = 10'h1bc == r_count_15_io_out ? io_r_444_b : _GEN_11783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11785 = 10'h1bd == r_count_15_io_out ? io_r_445_b : _GEN_11784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11786 = 10'h1be == r_count_15_io_out ? io_r_446_b : _GEN_11785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11787 = 10'h1bf == r_count_15_io_out ? io_r_447_b : _GEN_11786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11788 = 10'h1c0 == r_count_15_io_out ? io_r_448_b : _GEN_11787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11789 = 10'h1c1 == r_count_15_io_out ? io_r_449_b : _GEN_11788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11790 = 10'h1c2 == r_count_15_io_out ? io_r_450_b : _GEN_11789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11791 = 10'h1c3 == r_count_15_io_out ? io_r_451_b : _GEN_11790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11792 = 10'h1c4 == r_count_15_io_out ? io_r_452_b : _GEN_11791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11793 = 10'h1c5 == r_count_15_io_out ? io_r_453_b : _GEN_11792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11794 = 10'h1c6 == r_count_15_io_out ? io_r_454_b : _GEN_11793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11795 = 10'h1c7 == r_count_15_io_out ? io_r_455_b : _GEN_11794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11796 = 10'h1c8 == r_count_15_io_out ? io_r_456_b : _GEN_11795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11797 = 10'h1c9 == r_count_15_io_out ? io_r_457_b : _GEN_11796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11798 = 10'h1ca == r_count_15_io_out ? io_r_458_b : _GEN_11797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11799 = 10'h1cb == r_count_15_io_out ? io_r_459_b : _GEN_11798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11800 = 10'h1cc == r_count_15_io_out ? io_r_460_b : _GEN_11799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11801 = 10'h1cd == r_count_15_io_out ? io_r_461_b : _GEN_11800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11802 = 10'h1ce == r_count_15_io_out ? io_r_462_b : _GEN_11801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11803 = 10'h1cf == r_count_15_io_out ? io_r_463_b : _GEN_11802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11804 = 10'h1d0 == r_count_15_io_out ? io_r_464_b : _GEN_11803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11805 = 10'h1d1 == r_count_15_io_out ? io_r_465_b : _GEN_11804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11806 = 10'h1d2 == r_count_15_io_out ? io_r_466_b : _GEN_11805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11807 = 10'h1d3 == r_count_15_io_out ? io_r_467_b : _GEN_11806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11808 = 10'h1d4 == r_count_15_io_out ? io_r_468_b : _GEN_11807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11809 = 10'h1d5 == r_count_15_io_out ? io_r_469_b : _GEN_11808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11810 = 10'h1d6 == r_count_15_io_out ? io_r_470_b : _GEN_11809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11811 = 10'h1d7 == r_count_15_io_out ? io_r_471_b : _GEN_11810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11812 = 10'h1d8 == r_count_15_io_out ? io_r_472_b : _GEN_11811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11813 = 10'h1d9 == r_count_15_io_out ? io_r_473_b : _GEN_11812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11814 = 10'h1da == r_count_15_io_out ? io_r_474_b : _GEN_11813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11815 = 10'h1db == r_count_15_io_out ? io_r_475_b : _GEN_11814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11816 = 10'h1dc == r_count_15_io_out ? io_r_476_b : _GEN_11815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11817 = 10'h1dd == r_count_15_io_out ? io_r_477_b : _GEN_11816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11818 = 10'h1de == r_count_15_io_out ? io_r_478_b : _GEN_11817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11819 = 10'h1df == r_count_15_io_out ? io_r_479_b : _GEN_11818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11820 = 10'h1e0 == r_count_15_io_out ? io_r_480_b : _GEN_11819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11821 = 10'h1e1 == r_count_15_io_out ? io_r_481_b : _GEN_11820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11822 = 10'h1e2 == r_count_15_io_out ? io_r_482_b : _GEN_11821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11823 = 10'h1e3 == r_count_15_io_out ? io_r_483_b : _GEN_11822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11824 = 10'h1e4 == r_count_15_io_out ? io_r_484_b : _GEN_11823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11825 = 10'h1e5 == r_count_15_io_out ? io_r_485_b : _GEN_11824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11826 = 10'h1e6 == r_count_15_io_out ? io_r_486_b : _GEN_11825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11827 = 10'h1e7 == r_count_15_io_out ? io_r_487_b : _GEN_11826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11828 = 10'h1e8 == r_count_15_io_out ? io_r_488_b : _GEN_11827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11829 = 10'h1e9 == r_count_15_io_out ? io_r_489_b : _GEN_11828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11830 = 10'h1ea == r_count_15_io_out ? io_r_490_b : _GEN_11829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11831 = 10'h1eb == r_count_15_io_out ? io_r_491_b : _GEN_11830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11832 = 10'h1ec == r_count_15_io_out ? io_r_492_b : _GEN_11831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11833 = 10'h1ed == r_count_15_io_out ? io_r_493_b : _GEN_11832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11834 = 10'h1ee == r_count_15_io_out ? io_r_494_b : _GEN_11833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11835 = 10'h1ef == r_count_15_io_out ? io_r_495_b : _GEN_11834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11836 = 10'h1f0 == r_count_15_io_out ? io_r_496_b : _GEN_11835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11837 = 10'h1f1 == r_count_15_io_out ? io_r_497_b : _GEN_11836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11838 = 10'h1f2 == r_count_15_io_out ? io_r_498_b : _GEN_11837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11839 = 10'h1f3 == r_count_15_io_out ? io_r_499_b : _GEN_11838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11840 = 10'h1f4 == r_count_15_io_out ? io_r_500_b : _GEN_11839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11841 = 10'h1f5 == r_count_15_io_out ? io_r_501_b : _GEN_11840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11842 = 10'h1f6 == r_count_15_io_out ? io_r_502_b : _GEN_11841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11843 = 10'h1f7 == r_count_15_io_out ? io_r_503_b : _GEN_11842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11844 = 10'h1f8 == r_count_15_io_out ? io_r_504_b : _GEN_11843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11845 = 10'h1f9 == r_count_15_io_out ? io_r_505_b : _GEN_11844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11846 = 10'h1fa == r_count_15_io_out ? io_r_506_b : _GEN_11845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11847 = 10'h1fb == r_count_15_io_out ? io_r_507_b : _GEN_11846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11848 = 10'h1fc == r_count_15_io_out ? io_r_508_b : _GEN_11847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11849 = 10'h1fd == r_count_15_io_out ? io_r_509_b : _GEN_11848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11850 = 10'h1fe == r_count_15_io_out ? io_r_510_b : _GEN_11849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11851 = 10'h1ff == r_count_15_io_out ? io_r_511_b : _GEN_11850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11852 = 10'h200 == r_count_15_io_out ? io_r_512_b : _GEN_11851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11853 = 10'h201 == r_count_15_io_out ? io_r_513_b : _GEN_11852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11854 = 10'h202 == r_count_15_io_out ? io_r_514_b : _GEN_11853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11855 = 10'h203 == r_count_15_io_out ? io_r_515_b : _GEN_11854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11856 = 10'h204 == r_count_15_io_out ? io_r_516_b : _GEN_11855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11857 = 10'h205 == r_count_15_io_out ? io_r_517_b : _GEN_11856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11858 = 10'h206 == r_count_15_io_out ? io_r_518_b : _GEN_11857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11859 = 10'h207 == r_count_15_io_out ? io_r_519_b : _GEN_11858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11860 = 10'h208 == r_count_15_io_out ? io_r_520_b : _GEN_11859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11861 = 10'h209 == r_count_15_io_out ? io_r_521_b : _GEN_11860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11862 = 10'h20a == r_count_15_io_out ? io_r_522_b : _GEN_11861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11863 = 10'h20b == r_count_15_io_out ? io_r_523_b : _GEN_11862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11864 = 10'h20c == r_count_15_io_out ? io_r_524_b : _GEN_11863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11865 = 10'h20d == r_count_15_io_out ? io_r_525_b : _GEN_11864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11866 = 10'h20e == r_count_15_io_out ? io_r_526_b : _GEN_11865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11867 = 10'h20f == r_count_15_io_out ? io_r_527_b : _GEN_11866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11868 = 10'h210 == r_count_15_io_out ? io_r_528_b : _GEN_11867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11869 = 10'h211 == r_count_15_io_out ? io_r_529_b : _GEN_11868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11870 = 10'h212 == r_count_15_io_out ? io_r_530_b : _GEN_11869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11871 = 10'h213 == r_count_15_io_out ? io_r_531_b : _GEN_11870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11872 = 10'h214 == r_count_15_io_out ? io_r_532_b : _GEN_11871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11873 = 10'h215 == r_count_15_io_out ? io_r_533_b : _GEN_11872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11874 = 10'h216 == r_count_15_io_out ? io_r_534_b : _GEN_11873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11875 = 10'h217 == r_count_15_io_out ? io_r_535_b : _GEN_11874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11876 = 10'h218 == r_count_15_io_out ? io_r_536_b : _GEN_11875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11877 = 10'h219 == r_count_15_io_out ? io_r_537_b : _GEN_11876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11878 = 10'h21a == r_count_15_io_out ? io_r_538_b : _GEN_11877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11879 = 10'h21b == r_count_15_io_out ? io_r_539_b : _GEN_11878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11880 = 10'h21c == r_count_15_io_out ? io_r_540_b : _GEN_11879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11881 = 10'h21d == r_count_15_io_out ? io_r_541_b : _GEN_11880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11882 = 10'h21e == r_count_15_io_out ? io_r_542_b : _GEN_11881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11883 = 10'h21f == r_count_15_io_out ? io_r_543_b : _GEN_11882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11884 = 10'h220 == r_count_15_io_out ? io_r_544_b : _GEN_11883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11885 = 10'h221 == r_count_15_io_out ? io_r_545_b : _GEN_11884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11886 = 10'h222 == r_count_15_io_out ? io_r_546_b : _GEN_11885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11887 = 10'h223 == r_count_15_io_out ? io_r_547_b : _GEN_11886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11888 = 10'h224 == r_count_15_io_out ? io_r_548_b : _GEN_11887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11889 = 10'h225 == r_count_15_io_out ? io_r_549_b : _GEN_11888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11890 = 10'h226 == r_count_15_io_out ? io_r_550_b : _GEN_11889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11891 = 10'h227 == r_count_15_io_out ? io_r_551_b : _GEN_11890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11892 = 10'h228 == r_count_15_io_out ? io_r_552_b : _GEN_11891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11893 = 10'h229 == r_count_15_io_out ? io_r_553_b : _GEN_11892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11894 = 10'h22a == r_count_15_io_out ? io_r_554_b : _GEN_11893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11895 = 10'h22b == r_count_15_io_out ? io_r_555_b : _GEN_11894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11896 = 10'h22c == r_count_15_io_out ? io_r_556_b : _GEN_11895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11897 = 10'h22d == r_count_15_io_out ? io_r_557_b : _GEN_11896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11898 = 10'h22e == r_count_15_io_out ? io_r_558_b : _GEN_11897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11899 = 10'h22f == r_count_15_io_out ? io_r_559_b : _GEN_11898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11900 = 10'h230 == r_count_15_io_out ? io_r_560_b : _GEN_11899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11901 = 10'h231 == r_count_15_io_out ? io_r_561_b : _GEN_11900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11902 = 10'h232 == r_count_15_io_out ? io_r_562_b : _GEN_11901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11903 = 10'h233 == r_count_15_io_out ? io_r_563_b : _GEN_11902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11904 = 10'h234 == r_count_15_io_out ? io_r_564_b : _GEN_11903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11905 = 10'h235 == r_count_15_io_out ? io_r_565_b : _GEN_11904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11906 = 10'h236 == r_count_15_io_out ? io_r_566_b : _GEN_11905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11907 = 10'h237 == r_count_15_io_out ? io_r_567_b : _GEN_11906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11908 = 10'h238 == r_count_15_io_out ? io_r_568_b : _GEN_11907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11909 = 10'h239 == r_count_15_io_out ? io_r_569_b : _GEN_11908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11910 = 10'h23a == r_count_15_io_out ? io_r_570_b : _GEN_11909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11911 = 10'h23b == r_count_15_io_out ? io_r_571_b : _GEN_11910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11912 = 10'h23c == r_count_15_io_out ? io_r_572_b : _GEN_11911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11913 = 10'h23d == r_count_15_io_out ? io_r_573_b : _GEN_11912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11914 = 10'h23e == r_count_15_io_out ? io_r_574_b : _GEN_11913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11915 = 10'h23f == r_count_15_io_out ? io_r_575_b : _GEN_11914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11916 = 10'h240 == r_count_15_io_out ? io_r_576_b : _GEN_11915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11917 = 10'h241 == r_count_15_io_out ? io_r_577_b : _GEN_11916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11918 = 10'h242 == r_count_15_io_out ? io_r_578_b : _GEN_11917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11919 = 10'h243 == r_count_15_io_out ? io_r_579_b : _GEN_11918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11920 = 10'h244 == r_count_15_io_out ? io_r_580_b : _GEN_11919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11921 = 10'h245 == r_count_15_io_out ? io_r_581_b : _GEN_11920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11922 = 10'h246 == r_count_15_io_out ? io_r_582_b : _GEN_11921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11923 = 10'h247 == r_count_15_io_out ? io_r_583_b : _GEN_11922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11924 = 10'h248 == r_count_15_io_out ? io_r_584_b : _GEN_11923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11925 = 10'h249 == r_count_15_io_out ? io_r_585_b : _GEN_11924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11926 = 10'h24a == r_count_15_io_out ? io_r_586_b : _GEN_11925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11927 = 10'h24b == r_count_15_io_out ? io_r_587_b : _GEN_11926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11928 = 10'h24c == r_count_15_io_out ? io_r_588_b : _GEN_11927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11929 = 10'h24d == r_count_15_io_out ? io_r_589_b : _GEN_11928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11930 = 10'h24e == r_count_15_io_out ? io_r_590_b : _GEN_11929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11931 = 10'h24f == r_count_15_io_out ? io_r_591_b : _GEN_11930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11932 = 10'h250 == r_count_15_io_out ? io_r_592_b : _GEN_11931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11933 = 10'h251 == r_count_15_io_out ? io_r_593_b : _GEN_11932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11934 = 10'h252 == r_count_15_io_out ? io_r_594_b : _GEN_11933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11935 = 10'h253 == r_count_15_io_out ? io_r_595_b : _GEN_11934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11936 = 10'h254 == r_count_15_io_out ? io_r_596_b : _GEN_11935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11937 = 10'h255 == r_count_15_io_out ? io_r_597_b : _GEN_11936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11938 = 10'h256 == r_count_15_io_out ? io_r_598_b : _GEN_11937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11939 = 10'h257 == r_count_15_io_out ? io_r_599_b : _GEN_11938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11940 = 10'h258 == r_count_15_io_out ? io_r_600_b : _GEN_11939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11941 = 10'h259 == r_count_15_io_out ? io_r_601_b : _GEN_11940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11942 = 10'h25a == r_count_15_io_out ? io_r_602_b : _GEN_11941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11943 = 10'h25b == r_count_15_io_out ? io_r_603_b : _GEN_11942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11944 = 10'h25c == r_count_15_io_out ? io_r_604_b : _GEN_11943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11945 = 10'h25d == r_count_15_io_out ? io_r_605_b : _GEN_11944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11946 = 10'h25e == r_count_15_io_out ? io_r_606_b : _GEN_11945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11947 = 10'h25f == r_count_15_io_out ? io_r_607_b : _GEN_11946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11948 = 10'h260 == r_count_15_io_out ? io_r_608_b : _GEN_11947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11949 = 10'h261 == r_count_15_io_out ? io_r_609_b : _GEN_11948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11950 = 10'h262 == r_count_15_io_out ? io_r_610_b : _GEN_11949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11951 = 10'h263 == r_count_15_io_out ? io_r_611_b : _GEN_11950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11952 = 10'h264 == r_count_15_io_out ? io_r_612_b : _GEN_11951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11953 = 10'h265 == r_count_15_io_out ? io_r_613_b : _GEN_11952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11954 = 10'h266 == r_count_15_io_out ? io_r_614_b : _GEN_11953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11955 = 10'h267 == r_count_15_io_out ? io_r_615_b : _GEN_11954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11956 = 10'h268 == r_count_15_io_out ? io_r_616_b : _GEN_11955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11957 = 10'h269 == r_count_15_io_out ? io_r_617_b : _GEN_11956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11958 = 10'h26a == r_count_15_io_out ? io_r_618_b : _GEN_11957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11959 = 10'h26b == r_count_15_io_out ? io_r_619_b : _GEN_11958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11960 = 10'h26c == r_count_15_io_out ? io_r_620_b : _GEN_11959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11961 = 10'h26d == r_count_15_io_out ? io_r_621_b : _GEN_11960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11962 = 10'h26e == r_count_15_io_out ? io_r_622_b : _GEN_11961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11963 = 10'h26f == r_count_15_io_out ? io_r_623_b : _GEN_11962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11964 = 10'h270 == r_count_15_io_out ? io_r_624_b : _GEN_11963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11965 = 10'h271 == r_count_15_io_out ? io_r_625_b : _GEN_11964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11966 = 10'h272 == r_count_15_io_out ? io_r_626_b : _GEN_11965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11967 = 10'h273 == r_count_15_io_out ? io_r_627_b : _GEN_11966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11968 = 10'h274 == r_count_15_io_out ? io_r_628_b : _GEN_11967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11969 = 10'h275 == r_count_15_io_out ? io_r_629_b : _GEN_11968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11970 = 10'h276 == r_count_15_io_out ? io_r_630_b : _GEN_11969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11971 = 10'h277 == r_count_15_io_out ? io_r_631_b : _GEN_11970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11972 = 10'h278 == r_count_15_io_out ? io_r_632_b : _GEN_11971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11973 = 10'h279 == r_count_15_io_out ? io_r_633_b : _GEN_11972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11974 = 10'h27a == r_count_15_io_out ? io_r_634_b : _GEN_11973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11975 = 10'h27b == r_count_15_io_out ? io_r_635_b : _GEN_11974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11976 = 10'h27c == r_count_15_io_out ? io_r_636_b : _GEN_11975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11977 = 10'h27d == r_count_15_io_out ? io_r_637_b : _GEN_11976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11978 = 10'h27e == r_count_15_io_out ? io_r_638_b : _GEN_11977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11979 = 10'h27f == r_count_15_io_out ? io_r_639_b : _GEN_11978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11980 = 10'h280 == r_count_15_io_out ? io_r_640_b : _GEN_11979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11981 = 10'h281 == r_count_15_io_out ? io_r_641_b : _GEN_11980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11982 = 10'h282 == r_count_15_io_out ? io_r_642_b : _GEN_11981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11983 = 10'h283 == r_count_15_io_out ? io_r_643_b : _GEN_11982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11984 = 10'h284 == r_count_15_io_out ? io_r_644_b : _GEN_11983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11985 = 10'h285 == r_count_15_io_out ? io_r_645_b : _GEN_11984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11986 = 10'h286 == r_count_15_io_out ? io_r_646_b : _GEN_11985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11987 = 10'h287 == r_count_15_io_out ? io_r_647_b : _GEN_11986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11988 = 10'h288 == r_count_15_io_out ? io_r_648_b : _GEN_11987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11989 = 10'h289 == r_count_15_io_out ? io_r_649_b : _GEN_11988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11990 = 10'h28a == r_count_15_io_out ? io_r_650_b : _GEN_11989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11991 = 10'h28b == r_count_15_io_out ? io_r_651_b : _GEN_11990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11992 = 10'h28c == r_count_15_io_out ? io_r_652_b : _GEN_11991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11993 = 10'h28d == r_count_15_io_out ? io_r_653_b : _GEN_11992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11994 = 10'h28e == r_count_15_io_out ? io_r_654_b : _GEN_11993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11995 = 10'h28f == r_count_15_io_out ? io_r_655_b : _GEN_11994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11996 = 10'h290 == r_count_15_io_out ? io_r_656_b : _GEN_11995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11997 = 10'h291 == r_count_15_io_out ? io_r_657_b : _GEN_11996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11998 = 10'h292 == r_count_15_io_out ? io_r_658_b : _GEN_11997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11999 = 10'h293 == r_count_15_io_out ? io_r_659_b : _GEN_11998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12000 = 10'h294 == r_count_15_io_out ? io_r_660_b : _GEN_11999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12001 = 10'h295 == r_count_15_io_out ? io_r_661_b : _GEN_12000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12002 = 10'h296 == r_count_15_io_out ? io_r_662_b : _GEN_12001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12003 = 10'h297 == r_count_15_io_out ? io_r_663_b : _GEN_12002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12004 = 10'h298 == r_count_15_io_out ? io_r_664_b : _GEN_12003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12005 = 10'h299 == r_count_15_io_out ? io_r_665_b : _GEN_12004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12006 = 10'h29a == r_count_15_io_out ? io_r_666_b : _GEN_12005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12007 = 10'h29b == r_count_15_io_out ? io_r_667_b : _GEN_12006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12008 = 10'h29c == r_count_15_io_out ? io_r_668_b : _GEN_12007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12009 = 10'h29d == r_count_15_io_out ? io_r_669_b : _GEN_12008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12010 = 10'h29e == r_count_15_io_out ? io_r_670_b : _GEN_12009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12011 = 10'h29f == r_count_15_io_out ? io_r_671_b : _GEN_12010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12012 = 10'h2a0 == r_count_15_io_out ? io_r_672_b : _GEN_12011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12013 = 10'h2a1 == r_count_15_io_out ? io_r_673_b : _GEN_12012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12014 = 10'h2a2 == r_count_15_io_out ? io_r_674_b : _GEN_12013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12015 = 10'h2a3 == r_count_15_io_out ? io_r_675_b : _GEN_12014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12016 = 10'h2a4 == r_count_15_io_out ? io_r_676_b : _GEN_12015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12017 = 10'h2a5 == r_count_15_io_out ? io_r_677_b : _GEN_12016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12018 = 10'h2a6 == r_count_15_io_out ? io_r_678_b : _GEN_12017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12019 = 10'h2a7 == r_count_15_io_out ? io_r_679_b : _GEN_12018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12020 = 10'h2a8 == r_count_15_io_out ? io_r_680_b : _GEN_12019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12021 = 10'h2a9 == r_count_15_io_out ? io_r_681_b : _GEN_12020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12022 = 10'h2aa == r_count_15_io_out ? io_r_682_b : _GEN_12021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12023 = 10'h2ab == r_count_15_io_out ? io_r_683_b : _GEN_12022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12024 = 10'h2ac == r_count_15_io_out ? io_r_684_b : _GEN_12023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12025 = 10'h2ad == r_count_15_io_out ? io_r_685_b : _GEN_12024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12026 = 10'h2ae == r_count_15_io_out ? io_r_686_b : _GEN_12025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12027 = 10'h2af == r_count_15_io_out ? io_r_687_b : _GEN_12026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12028 = 10'h2b0 == r_count_15_io_out ? io_r_688_b : _GEN_12027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12029 = 10'h2b1 == r_count_15_io_out ? io_r_689_b : _GEN_12028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12030 = 10'h2b2 == r_count_15_io_out ? io_r_690_b : _GEN_12029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12031 = 10'h2b3 == r_count_15_io_out ? io_r_691_b : _GEN_12030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12032 = 10'h2b4 == r_count_15_io_out ? io_r_692_b : _GEN_12031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12033 = 10'h2b5 == r_count_15_io_out ? io_r_693_b : _GEN_12032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12034 = 10'h2b6 == r_count_15_io_out ? io_r_694_b : _GEN_12033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12035 = 10'h2b7 == r_count_15_io_out ? io_r_695_b : _GEN_12034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12036 = 10'h2b8 == r_count_15_io_out ? io_r_696_b : _GEN_12035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12037 = 10'h2b9 == r_count_15_io_out ? io_r_697_b : _GEN_12036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12038 = 10'h2ba == r_count_15_io_out ? io_r_698_b : _GEN_12037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12039 = 10'h2bb == r_count_15_io_out ? io_r_699_b : _GEN_12038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12040 = 10'h2bc == r_count_15_io_out ? io_r_700_b : _GEN_12039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12041 = 10'h2bd == r_count_15_io_out ? io_r_701_b : _GEN_12040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12042 = 10'h2be == r_count_15_io_out ? io_r_702_b : _GEN_12041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12043 = 10'h2bf == r_count_15_io_out ? io_r_703_b : _GEN_12042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12044 = 10'h2c0 == r_count_15_io_out ? io_r_704_b : _GEN_12043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12045 = 10'h2c1 == r_count_15_io_out ? io_r_705_b : _GEN_12044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12046 = 10'h2c2 == r_count_15_io_out ? io_r_706_b : _GEN_12045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12047 = 10'h2c3 == r_count_15_io_out ? io_r_707_b : _GEN_12046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12048 = 10'h2c4 == r_count_15_io_out ? io_r_708_b : _GEN_12047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12049 = 10'h2c5 == r_count_15_io_out ? io_r_709_b : _GEN_12048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12050 = 10'h2c6 == r_count_15_io_out ? io_r_710_b : _GEN_12049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12051 = 10'h2c7 == r_count_15_io_out ? io_r_711_b : _GEN_12050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12052 = 10'h2c8 == r_count_15_io_out ? io_r_712_b : _GEN_12051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12053 = 10'h2c9 == r_count_15_io_out ? io_r_713_b : _GEN_12052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12054 = 10'h2ca == r_count_15_io_out ? io_r_714_b : _GEN_12053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12055 = 10'h2cb == r_count_15_io_out ? io_r_715_b : _GEN_12054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12056 = 10'h2cc == r_count_15_io_out ? io_r_716_b : _GEN_12055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12057 = 10'h2cd == r_count_15_io_out ? io_r_717_b : _GEN_12056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12058 = 10'h2ce == r_count_15_io_out ? io_r_718_b : _GEN_12057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12059 = 10'h2cf == r_count_15_io_out ? io_r_719_b : _GEN_12058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12060 = 10'h2d0 == r_count_15_io_out ? io_r_720_b : _GEN_12059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12061 = 10'h2d1 == r_count_15_io_out ? io_r_721_b : _GEN_12060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12062 = 10'h2d2 == r_count_15_io_out ? io_r_722_b : _GEN_12061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12063 = 10'h2d3 == r_count_15_io_out ? io_r_723_b : _GEN_12062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12064 = 10'h2d4 == r_count_15_io_out ? io_r_724_b : _GEN_12063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12065 = 10'h2d5 == r_count_15_io_out ? io_r_725_b : _GEN_12064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12066 = 10'h2d6 == r_count_15_io_out ? io_r_726_b : _GEN_12065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12067 = 10'h2d7 == r_count_15_io_out ? io_r_727_b : _GEN_12066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12068 = 10'h2d8 == r_count_15_io_out ? io_r_728_b : _GEN_12067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12069 = 10'h2d9 == r_count_15_io_out ? io_r_729_b : _GEN_12068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12070 = 10'h2da == r_count_15_io_out ? io_r_730_b : _GEN_12069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12071 = 10'h2db == r_count_15_io_out ? io_r_731_b : _GEN_12070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12072 = 10'h2dc == r_count_15_io_out ? io_r_732_b : _GEN_12071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12073 = 10'h2dd == r_count_15_io_out ? io_r_733_b : _GEN_12072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12074 = 10'h2de == r_count_15_io_out ? io_r_734_b : _GEN_12073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12075 = 10'h2df == r_count_15_io_out ? io_r_735_b : _GEN_12074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12076 = 10'h2e0 == r_count_15_io_out ? io_r_736_b : _GEN_12075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12077 = 10'h2e1 == r_count_15_io_out ? io_r_737_b : _GEN_12076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12078 = 10'h2e2 == r_count_15_io_out ? io_r_738_b : _GEN_12077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12079 = 10'h2e3 == r_count_15_io_out ? io_r_739_b : _GEN_12078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12080 = 10'h2e4 == r_count_15_io_out ? io_r_740_b : _GEN_12079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12081 = 10'h2e5 == r_count_15_io_out ? io_r_741_b : _GEN_12080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12082 = 10'h2e6 == r_count_15_io_out ? io_r_742_b : _GEN_12081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12083 = 10'h2e7 == r_count_15_io_out ? io_r_743_b : _GEN_12082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12084 = 10'h2e8 == r_count_15_io_out ? io_r_744_b : _GEN_12083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12085 = 10'h2e9 == r_count_15_io_out ? io_r_745_b : _GEN_12084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12086 = 10'h2ea == r_count_15_io_out ? io_r_746_b : _GEN_12085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12087 = 10'h2eb == r_count_15_io_out ? io_r_747_b : _GEN_12086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12088 = 10'h2ec == r_count_15_io_out ? io_r_748_b : _GEN_12087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12091 = 10'h1 == r_count_16_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12092 = 10'h2 == r_count_16_io_out ? io_r_2_b : _GEN_12091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12093 = 10'h3 == r_count_16_io_out ? io_r_3_b : _GEN_12092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12094 = 10'h4 == r_count_16_io_out ? io_r_4_b : _GEN_12093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12095 = 10'h5 == r_count_16_io_out ? io_r_5_b : _GEN_12094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12096 = 10'h6 == r_count_16_io_out ? io_r_6_b : _GEN_12095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12097 = 10'h7 == r_count_16_io_out ? io_r_7_b : _GEN_12096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12098 = 10'h8 == r_count_16_io_out ? io_r_8_b : _GEN_12097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12099 = 10'h9 == r_count_16_io_out ? io_r_9_b : _GEN_12098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12100 = 10'ha == r_count_16_io_out ? io_r_10_b : _GEN_12099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12101 = 10'hb == r_count_16_io_out ? io_r_11_b : _GEN_12100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12102 = 10'hc == r_count_16_io_out ? io_r_12_b : _GEN_12101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12103 = 10'hd == r_count_16_io_out ? io_r_13_b : _GEN_12102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12104 = 10'he == r_count_16_io_out ? io_r_14_b : _GEN_12103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12105 = 10'hf == r_count_16_io_out ? io_r_15_b : _GEN_12104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12106 = 10'h10 == r_count_16_io_out ? io_r_16_b : _GEN_12105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12107 = 10'h11 == r_count_16_io_out ? io_r_17_b : _GEN_12106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12108 = 10'h12 == r_count_16_io_out ? io_r_18_b : _GEN_12107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12109 = 10'h13 == r_count_16_io_out ? io_r_19_b : _GEN_12108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12110 = 10'h14 == r_count_16_io_out ? io_r_20_b : _GEN_12109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12111 = 10'h15 == r_count_16_io_out ? io_r_21_b : _GEN_12110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12112 = 10'h16 == r_count_16_io_out ? io_r_22_b : _GEN_12111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12113 = 10'h17 == r_count_16_io_out ? io_r_23_b : _GEN_12112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12114 = 10'h18 == r_count_16_io_out ? io_r_24_b : _GEN_12113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12115 = 10'h19 == r_count_16_io_out ? io_r_25_b : _GEN_12114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12116 = 10'h1a == r_count_16_io_out ? io_r_26_b : _GEN_12115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12117 = 10'h1b == r_count_16_io_out ? io_r_27_b : _GEN_12116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12118 = 10'h1c == r_count_16_io_out ? io_r_28_b : _GEN_12117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12119 = 10'h1d == r_count_16_io_out ? io_r_29_b : _GEN_12118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12120 = 10'h1e == r_count_16_io_out ? io_r_30_b : _GEN_12119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12121 = 10'h1f == r_count_16_io_out ? io_r_31_b : _GEN_12120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12122 = 10'h20 == r_count_16_io_out ? io_r_32_b : _GEN_12121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12123 = 10'h21 == r_count_16_io_out ? io_r_33_b : _GEN_12122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12124 = 10'h22 == r_count_16_io_out ? io_r_34_b : _GEN_12123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12125 = 10'h23 == r_count_16_io_out ? io_r_35_b : _GEN_12124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12126 = 10'h24 == r_count_16_io_out ? io_r_36_b : _GEN_12125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12127 = 10'h25 == r_count_16_io_out ? io_r_37_b : _GEN_12126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12128 = 10'h26 == r_count_16_io_out ? io_r_38_b : _GEN_12127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12129 = 10'h27 == r_count_16_io_out ? io_r_39_b : _GEN_12128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12130 = 10'h28 == r_count_16_io_out ? io_r_40_b : _GEN_12129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12131 = 10'h29 == r_count_16_io_out ? io_r_41_b : _GEN_12130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12132 = 10'h2a == r_count_16_io_out ? io_r_42_b : _GEN_12131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12133 = 10'h2b == r_count_16_io_out ? io_r_43_b : _GEN_12132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12134 = 10'h2c == r_count_16_io_out ? io_r_44_b : _GEN_12133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12135 = 10'h2d == r_count_16_io_out ? io_r_45_b : _GEN_12134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12136 = 10'h2e == r_count_16_io_out ? io_r_46_b : _GEN_12135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12137 = 10'h2f == r_count_16_io_out ? io_r_47_b : _GEN_12136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12138 = 10'h30 == r_count_16_io_out ? io_r_48_b : _GEN_12137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12139 = 10'h31 == r_count_16_io_out ? io_r_49_b : _GEN_12138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12140 = 10'h32 == r_count_16_io_out ? io_r_50_b : _GEN_12139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12141 = 10'h33 == r_count_16_io_out ? io_r_51_b : _GEN_12140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12142 = 10'h34 == r_count_16_io_out ? io_r_52_b : _GEN_12141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12143 = 10'h35 == r_count_16_io_out ? io_r_53_b : _GEN_12142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12144 = 10'h36 == r_count_16_io_out ? io_r_54_b : _GEN_12143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12145 = 10'h37 == r_count_16_io_out ? io_r_55_b : _GEN_12144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12146 = 10'h38 == r_count_16_io_out ? io_r_56_b : _GEN_12145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12147 = 10'h39 == r_count_16_io_out ? io_r_57_b : _GEN_12146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12148 = 10'h3a == r_count_16_io_out ? io_r_58_b : _GEN_12147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12149 = 10'h3b == r_count_16_io_out ? io_r_59_b : _GEN_12148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12150 = 10'h3c == r_count_16_io_out ? io_r_60_b : _GEN_12149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12151 = 10'h3d == r_count_16_io_out ? io_r_61_b : _GEN_12150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12152 = 10'h3e == r_count_16_io_out ? io_r_62_b : _GEN_12151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12153 = 10'h3f == r_count_16_io_out ? io_r_63_b : _GEN_12152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12154 = 10'h40 == r_count_16_io_out ? io_r_64_b : _GEN_12153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12155 = 10'h41 == r_count_16_io_out ? io_r_65_b : _GEN_12154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12156 = 10'h42 == r_count_16_io_out ? io_r_66_b : _GEN_12155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12157 = 10'h43 == r_count_16_io_out ? io_r_67_b : _GEN_12156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12158 = 10'h44 == r_count_16_io_out ? io_r_68_b : _GEN_12157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12159 = 10'h45 == r_count_16_io_out ? io_r_69_b : _GEN_12158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12160 = 10'h46 == r_count_16_io_out ? io_r_70_b : _GEN_12159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12161 = 10'h47 == r_count_16_io_out ? io_r_71_b : _GEN_12160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12162 = 10'h48 == r_count_16_io_out ? io_r_72_b : _GEN_12161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12163 = 10'h49 == r_count_16_io_out ? io_r_73_b : _GEN_12162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12164 = 10'h4a == r_count_16_io_out ? io_r_74_b : _GEN_12163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12165 = 10'h4b == r_count_16_io_out ? io_r_75_b : _GEN_12164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12166 = 10'h4c == r_count_16_io_out ? io_r_76_b : _GEN_12165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12167 = 10'h4d == r_count_16_io_out ? io_r_77_b : _GEN_12166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12168 = 10'h4e == r_count_16_io_out ? io_r_78_b : _GEN_12167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12169 = 10'h4f == r_count_16_io_out ? io_r_79_b : _GEN_12168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12170 = 10'h50 == r_count_16_io_out ? io_r_80_b : _GEN_12169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12171 = 10'h51 == r_count_16_io_out ? io_r_81_b : _GEN_12170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12172 = 10'h52 == r_count_16_io_out ? io_r_82_b : _GEN_12171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12173 = 10'h53 == r_count_16_io_out ? io_r_83_b : _GEN_12172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12174 = 10'h54 == r_count_16_io_out ? io_r_84_b : _GEN_12173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12175 = 10'h55 == r_count_16_io_out ? io_r_85_b : _GEN_12174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12176 = 10'h56 == r_count_16_io_out ? io_r_86_b : _GEN_12175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12177 = 10'h57 == r_count_16_io_out ? io_r_87_b : _GEN_12176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12178 = 10'h58 == r_count_16_io_out ? io_r_88_b : _GEN_12177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12179 = 10'h59 == r_count_16_io_out ? io_r_89_b : _GEN_12178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12180 = 10'h5a == r_count_16_io_out ? io_r_90_b : _GEN_12179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12181 = 10'h5b == r_count_16_io_out ? io_r_91_b : _GEN_12180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12182 = 10'h5c == r_count_16_io_out ? io_r_92_b : _GEN_12181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12183 = 10'h5d == r_count_16_io_out ? io_r_93_b : _GEN_12182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12184 = 10'h5e == r_count_16_io_out ? io_r_94_b : _GEN_12183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12185 = 10'h5f == r_count_16_io_out ? io_r_95_b : _GEN_12184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12186 = 10'h60 == r_count_16_io_out ? io_r_96_b : _GEN_12185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12187 = 10'h61 == r_count_16_io_out ? io_r_97_b : _GEN_12186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12188 = 10'h62 == r_count_16_io_out ? io_r_98_b : _GEN_12187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12189 = 10'h63 == r_count_16_io_out ? io_r_99_b : _GEN_12188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12190 = 10'h64 == r_count_16_io_out ? io_r_100_b : _GEN_12189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12191 = 10'h65 == r_count_16_io_out ? io_r_101_b : _GEN_12190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12192 = 10'h66 == r_count_16_io_out ? io_r_102_b : _GEN_12191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12193 = 10'h67 == r_count_16_io_out ? io_r_103_b : _GEN_12192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12194 = 10'h68 == r_count_16_io_out ? io_r_104_b : _GEN_12193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12195 = 10'h69 == r_count_16_io_out ? io_r_105_b : _GEN_12194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12196 = 10'h6a == r_count_16_io_out ? io_r_106_b : _GEN_12195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12197 = 10'h6b == r_count_16_io_out ? io_r_107_b : _GEN_12196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12198 = 10'h6c == r_count_16_io_out ? io_r_108_b : _GEN_12197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12199 = 10'h6d == r_count_16_io_out ? io_r_109_b : _GEN_12198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12200 = 10'h6e == r_count_16_io_out ? io_r_110_b : _GEN_12199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12201 = 10'h6f == r_count_16_io_out ? io_r_111_b : _GEN_12200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12202 = 10'h70 == r_count_16_io_out ? io_r_112_b : _GEN_12201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12203 = 10'h71 == r_count_16_io_out ? io_r_113_b : _GEN_12202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12204 = 10'h72 == r_count_16_io_out ? io_r_114_b : _GEN_12203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12205 = 10'h73 == r_count_16_io_out ? io_r_115_b : _GEN_12204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12206 = 10'h74 == r_count_16_io_out ? io_r_116_b : _GEN_12205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12207 = 10'h75 == r_count_16_io_out ? io_r_117_b : _GEN_12206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12208 = 10'h76 == r_count_16_io_out ? io_r_118_b : _GEN_12207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12209 = 10'h77 == r_count_16_io_out ? io_r_119_b : _GEN_12208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12210 = 10'h78 == r_count_16_io_out ? io_r_120_b : _GEN_12209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12211 = 10'h79 == r_count_16_io_out ? io_r_121_b : _GEN_12210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12212 = 10'h7a == r_count_16_io_out ? io_r_122_b : _GEN_12211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12213 = 10'h7b == r_count_16_io_out ? io_r_123_b : _GEN_12212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12214 = 10'h7c == r_count_16_io_out ? io_r_124_b : _GEN_12213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12215 = 10'h7d == r_count_16_io_out ? io_r_125_b : _GEN_12214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12216 = 10'h7e == r_count_16_io_out ? io_r_126_b : _GEN_12215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12217 = 10'h7f == r_count_16_io_out ? io_r_127_b : _GEN_12216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12218 = 10'h80 == r_count_16_io_out ? io_r_128_b : _GEN_12217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12219 = 10'h81 == r_count_16_io_out ? io_r_129_b : _GEN_12218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12220 = 10'h82 == r_count_16_io_out ? io_r_130_b : _GEN_12219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12221 = 10'h83 == r_count_16_io_out ? io_r_131_b : _GEN_12220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12222 = 10'h84 == r_count_16_io_out ? io_r_132_b : _GEN_12221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12223 = 10'h85 == r_count_16_io_out ? io_r_133_b : _GEN_12222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12224 = 10'h86 == r_count_16_io_out ? io_r_134_b : _GEN_12223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12225 = 10'h87 == r_count_16_io_out ? io_r_135_b : _GEN_12224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12226 = 10'h88 == r_count_16_io_out ? io_r_136_b : _GEN_12225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12227 = 10'h89 == r_count_16_io_out ? io_r_137_b : _GEN_12226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12228 = 10'h8a == r_count_16_io_out ? io_r_138_b : _GEN_12227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12229 = 10'h8b == r_count_16_io_out ? io_r_139_b : _GEN_12228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12230 = 10'h8c == r_count_16_io_out ? io_r_140_b : _GEN_12229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12231 = 10'h8d == r_count_16_io_out ? io_r_141_b : _GEN_12230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12232 = 10'h8e == r_count_16_io_out ? io_r_142_b : _GEN_12231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12233 = 10'h8f == r_count_16_io_out ? io_r_143_b : _GEN_12232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12234 = 10'h90 == r_count_16_io_out ? io_r_144_b : _GEN_12233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12235 = 10'h91 == r_count_16_io_out ? io_r_145_b : _GEN_12234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12236 = 10'h92 == r_count_16_io_out ? io_r_146_b : _GEN_12235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12237 = 10'h93 == r_count_16_io_out ? io_r_147_b : _GEN_12236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12238 = 10'h94 == r_count_16_io_out ? io_r_148_b : _GEN_12237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12239 = 10'h95 == r_count_16_io_out ? io_r_149_b : _GEN_12238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12240 = 10'h96 == r_count_16_io_out ? io_r_150_b : _GEN_12239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12241 = 10'h97 == r_count_16_io_out ? io_r_151_b : _GEN_12240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12242 = 10'h98 == r_count_16_io_out ? io_r_152_b : _GEN_12241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12243 = 10'h99 == r_count_16_io_out ? io_r_153_b : _GEN_12242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12244 = 10'h9a == r_count_16_io_out ? io_r_154_b : _GEN_12243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12245 = 10'h9b == r_count_16_io_out ? io_r_155_b : _GEN_12244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12246 = 10'h9c == r_count_16_io_out ? io_r_156_b : _GEN_12245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12247 = 10'h9d == r_count_16_io_out ? io_r_157_b : _GEN_12246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12248 = 10'h9e == r_count_16_io_out ? io_r_158_b : _GEN_12247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12249 = 10'h9f == r_count_16_io_out ? io_r_159_b : _GEN_12248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12250 = 10'ha0 == r_count_16_io_out ? io_r_160_b : _GEN_12249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12251 = 10'ha1 == r_count_16_io_out ? io_r_161_b : _GEN_12250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12252 = 10'ha2 == r_count_16_io_out ? io_r_162_b : _GEN_12251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12253 = 10'ha3 == r_count_16_io_out ? io_r_163_b : _GEN_12252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12254 = 10'ha4 == r_count_16_io_out ? io_r_164_b : _GEN_12253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12255 = 10'ha5 == r_count_16_io_out ? io_r_165_b : _GEN_12254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12256 = 10'ha6 == r_count_16_io_out ? io_r_166_b : _GEN_12255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12257 = 10'ha7 == r_count_16_io_out ? io_r_167_b : _GEN_12256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12258 = 10'ha8 == r_count_16_io_out ? io_r_168_b : _GEN_12257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12259 = 10'ha9 == r_count_16_io_out ? io_r_169_b : _GEN_12258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12260 = 10'haa == r_count_16_io_out ? io_r_170_b : _GEN_12259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12261 = 10'hab == r_count_16_io_out ? io_r_171_b : _GEN_12260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12262 = 10'hac == r_count_16_io_out ? io_r_172_b : _GEN_12261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12263 = 10'had == r_count_16_io_out ? io_r_173_b : _GEN_12262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12264 = 10'hae == r_count_16_io_out ? io_r_174_b : _GEN_12263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12265 = 10'haf == r_count_16_io_out ? io_r_175_b : _GEN_12264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12266 = 10'hb0 == r_count_16_io_out ? io_r_176_b : _GEN_12265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12267 = 10'hb1 == r_count_16_io_out ? io_r_177_b : _GEN_12266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12268 = 10'hb2 == r_count_16_io_out ? io_r_178_b : _GEN_12267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12269 = 10'hb3 == r_count_16_io_out ? io_r_179_b : _GEN_12268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12270 = 10'hb4 == r_count_16_io_out ? io_r_180_b : _GEN_12269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12271 = 10'hb5 == r_count_16_io_out ? io_r_181_b : _GEN_12270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12272 = 10'hb6 == r_count_16_io_out ? io_r_182_b : _GEN_12271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12273 = 10'hb7 == r_count_16_io_out ? io_r_183_b : _GEN_12272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12274 = 10'hb8 == r_count_16_io_out ? io_r_184_b : _GEN_12273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12275 = 10'hb9 == r_count_16_io_out ? io_r_185_b : _GEN_12274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12276 = 10'hba == r_count_16_io_out ? io_r_186_b : _GEN_12275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12277 = 10'hbb == r_count_16_io_out ? io_r_187_b : _GEN_12276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12278 = 10'hbc == r_count_16_io_out ? io_r_188_b : _GEN_12277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12279 = 10'hbd == r_count_16_io_out ? io_r_189_b : _GEN_12278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12280 = 10'hbe == r_count_16_io_out ? io_r_190_b : _GEN_12279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12281 = 10'hbf == r_count_16_io_out ? io_r_191_b : _GEN_12280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12282 = 10'hc0 == r_count_16_io_out ? io_r_192_b : _GEN_12281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12283 = 10'hc1 == r_count_16_io_out ? io_r_193_b : _GEN_12282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12284 = 10'hc2 == r_count_16_io_out ? io_r_194_b : _GEN_12283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12285 = 10'hc3 == r_count_16_io_out ? io_r_195_b : _GEN_12284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12286 = 10'hc4 == r_count_16_io_out ? io_r_196_b : _GEN_12285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12287 = 10'hc5 == r_count_16_io_out ? io_r_197_b : _GEN_12286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12288 = 10'hc6 == r_count_16_io_out ? io_r_198_b : _GEN_12287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12289 = 10'hc7 == r_count_16_io_out ? io_r_199_b : _GEN_12288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12290 = 10'hc8 == r_count_16_io_out ? io_r_200_b : _GEN_12289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12291 = 10'hc9 == r_count_16_io_out ? io_r_201_b : _GEN_12290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12292 = 10'hca == r_count_16_io_out ? io_r_202_b : _GEN_12291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12293 = 10'hcb == r_count_16_io_out ? io_r_203_b : _GEN_12292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12294 = 10'hcc == r_count_16_io_out ? io_r_204_b : _GEN_12293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12295 = 10'hcd == r_count_16_io_out ? io_r_205_b : _GEN_12294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12296 = 10'hce == r_count_16_io_out ? io_r_206_b : _GEN_12295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12297 = 10'hcf == r_count_16_io_out ? io_r_207_b : _GEN_12296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12298 = 10'hd0 == r_count_16_io_out ? io_r_208_b : _GEN_12297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12299 = 10'hd1 == r_count_16_io_out ? io_r_209_b : _GEN_12298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12300 = 10'hd2 == r_count_16_io_out ? io_r_210_b : _GEN_12299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12301 = 10'hd3 == r_count_16_io_out ? io_r_211_b : _GEN_12300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12302 = 10'hd4 == r_count_16_io_out ? io_r_212_b : _GEN_12301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12303 = 10'hd5 == r_count_16_io_out ? io_r_213_b : _GEN_12302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12304 = 10'hd6 == r_count_16_io_out ? io_r_214_b : _GEN_12303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12305 = 10'hd7 == r_count_16_io_out ? io_r_215_b : _GEN_12304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12306 = 10'hd8 == r_count_16_io_out ? io_r_216_b : _GEN_12305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12307 = 10'hd9 == r_count_16_io_out ? io_r_217_b : _GEN_12306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12308 = 10'hda == r_count_16_io_out ? io_r_218_b : _GEN_12307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12309 = 10'hdb == r_count_16_io_out ? io_r_219_b : _GEN_12308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12310 = 10'hdc == r_count_16_io_out ? io_r_220_b : _GEN_12309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12311 = 10'hdd == r_count_16_io_out ? io_r_221_b : _GEN_12310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12312 = 10'hde == r_count_16_io_out ? io_r_222_b : _GEN_12311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12313 = 10'hdf == r_count_16_io_out ? io_r_223_b : _GEN_12312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12314 = 10'he0 == r_count_16_io_out ? io_r_224_b : _GEN_12313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12315 = 10'he1 == r_count_16_io_out ? io_r_225_b : _GEN_12314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12316 = 10'he2 == r_count_16_io_out ? io_r_226_b : _GEN_12315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12317 = 10'he3 == r_count_16_io_out ? io_r_227_b : _GEN_12316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12318 = 10'he4 == r_count_16_io_out ? io_r_228_b : _GEN_12317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12319 = 10'he5 == r_count_16_io_out ? io_r_229_b : _GEN_12318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12320 = 10'he6 == r_count_16_io_out ? io_r_230_b : _GEN_12319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12321 = 10'he7 == r_count_16_io_out ? io_r_231_b : _GEN_12320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12322 = 10'he8 == r_count_16_io_out ? io_r_232_b : _GEN_12321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12323 = 10'he9 == r_count_16_io_out ? io_r_233_b : _GEN_12322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12324 = 10'hea == r_count_16_io_out ? io_r_234_b : _GEN_12323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12325 = 10'heb == r_count_16_io_out ? io_r_235_b : _GEN_12324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12326 = 10'hec == r_count_16_io_out ? io_r_236_b : _GEN_12325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12327 = 10'hed == r_count_16_io_out ? io_r_237_b : _GEN_12326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12328 = 10'hee == r_count_16_io_out ? io_r_238_b : _GEN_12327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12329 = 10'hef == r_count_16_io_out ? io_r_239_b : _GEN_12328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12330 = 10'hf0 == r_count_16_io_out ? io_r_240_b : _GEN_12329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12331 = 10'hf1 == r_count_16_io_out ? io_r_241_b : _GEN_12330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12332 = 10'hf2 == r_count_16_io_out ? io_r_242_b : _GEN_12331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12333 = 10'hf3 == r_count_16_io_out ? io_r_243_b : _GEN_12332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12334 = 10'hf4 == r_count_16_io_out ? io_r_244_b : _GEN_12333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12335 = 10'hf5 == r_count_16_io_out ? io_r_245_b : _GEN_12334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12336 = 10'hf6 == r_count_16_io_out ? io_r_246_b : _GEN_12335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12337 = 10'hf7 == r_count_16_io_out ? io_r_247_b : _GEN_12336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12338 = 10'hf8 == r_count_16_io_out ? io_r_248_b : _GEN_12337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12339 = 10'hf9 == r_count_16_io_out ? io_r_249_b : _GEN_12338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12340 = 10'hfa == r_count_16_io_out ? io_r_250_b : _GEN_12339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12341 = 10'hfb == r_count_16_io_out ? io_r_251_b : _GEN_12340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12342 = 10'hfc == r_count_16_io_out ? io_r_252_b : _GEN_12341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12343 = 10'hfd == r_count_16_io_out ? io_r_253_b : _GEN_12342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12344 = 10'hfe == r_count_16_io_out ? io_r_254_b : _GEN_12343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12345 = 10'hff == r_count_16_io_out ? io_r_255_b : _GEN_12344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12346 = 10'h100 == r_count_16_io_out ? io_r_256_b : _GEN_12345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12347 = 10'h101 == r_count_16_io_out ? io_r_257_b : _GEN_12346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12348 = 10'h102 == r_count_16_io_out ? io_r_258_b : _GEN_12347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12349 = 10'h103 == r_count_16_io_out ? io_r_259_b : _GEN_12348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12350 = 10'h104 == r_count_16_io_out ? io_r_260_b : _GEN_12349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12351 = 10'h105 == r_count_16_io_out ? io_r_261_b : _GEN_12350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12352 = 10'h106 == r_count_16_io_out ? io_r_262_b : _GEN_12351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12353 = 10'h107 == r_count_16_io_out ? io_r_263_b : _GEN_12352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12354 = 10'h108 == r_count_16_io_out ? io_r_264_b : _GEN_12353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12355 = 10'h109 == r_count_16_io_out ? io_r_265_b : _GEN_12354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12356 = 10'h10a == r_count_16_io_out ? io_r_266_b : _GEN_12355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12357 = 10'h10b == r_count_16_io_out ? io_r_267_b : _GEN_12356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12358 = 10'h10c == r_count_16_io_out ? io_r_268_b : _GEN_12357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12359 = 10'h10d == r_count_16_io_out ? io_r_269_b : _GEN_12358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12360 = 10'h10e == r_count_16_io_out ? io_r_270_b : _GEN_12359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12361 = 10'h10f == r_count_16_io_out ? io_r_271_b : _GEN_12360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12362 = 10'h110 == r_count_16_io_out ? io_r_272_b : _GEN_12361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12363 = 10'h111 == r_count_16_io_out ? io_r_273_b : _GEN_12362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12364 = 10'h112 == r_count_16_io_out ? io_r_274_b : _GEN_12363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12365 = 10'h113 == r_count_16_io_out ? io_r_275_b : _GEN_12364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12366 = 10'h114 == r_count_16_io_out ? io_r_276_b : _GEN_12365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12367 = 10'h115 == r_count_16_io_out ? io_r_277_b : _GEN_12366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12368 = 10'h116 == r_count_16_io_out ? io_r_278_b : _GEN_12367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12369 = 10'h117 == r_count_16_io_out ? io_r_279_b : _GEN_12368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12370 = 10'h118 == r_count_16_io_out ? io_r_280_b : _GEN_12369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12371 = 10'h119 == r_count_16_io_out ? io_r_281_b : _GEN_12370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12372 = 10'h11a == r_count_16_io_out ? io_r_282_b : _GEN_12371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12373 = 10'h11b == r_count_16_io_out ? io_r_283_b : _GEN_12372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12374 = 10'h11c == r_count_16_io_out ? io_r_284_b : _GEN_12373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12375 = 10'h11d == r_count_16_io_out ? io_r_285_b : _GEN_12374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12376 = 10'h11e == r_count_16_io_out ? io_r_286_b : _GEN_12375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12377 = 10'h11f == r_count_16_io_out ? io_r_287_b : _GEN_12376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12378 = 10'h120 == r_count_16_io_out ? io_r_288_b : _GEN_12377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12379 = 10'h121 == r_count_16_io_out ? io_r_289_b : _GEN_12378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12380 = 10'h122 == r_count_16_io_out ? io_r_290_b : _GEN_12379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12381 = 10'h123 == r_count_16_io_out ? io_r_291_b : _GEN_12380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12382 = 10'h124 == r_count_16_io_out ? io_r_292_b : _GEN_12381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12383 = 10'h125 == r_count_16_io_out ? io_r_293_b : _GEN_12382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12384 = 10'h126 == r_count_16_io_out ? io_r_294_b : _GEN_12383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12385 = 10'h127 == r_count_16_io_out ? io_r_295_b : _GEN_12384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12386 = 10'h128 == r_count_16_io_out ? io_r_296_b : _GEN_12385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12387 = 10'h129 == r_count_16_io_out ? io_r_297_b : _GEN_12386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12388 = 10'h12a == r_count_16_io_out ? io_r_298_b : _GEN_12387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12389 = 10'h12b == r_count_16_io_out ? io_r_299_b : _GEN_12388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12390 = 10'h12c == r_count_16_io_out ? io_r_300_b : _GEN_12389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12391 = 10'h12d == r_count_16_io_out ? io_r_301_b : _GEN_12390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12392 = 10'h12e == r_count_16_io_out ? io_r_302_b : _GEN_12391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12393 = 10'h12f == r_count_16_io_out ? io_r_303_b : _GEN_12392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12394 = 10'h130 == r_count_16_io_out ? io_r_304_b : _GEN_12393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12395 = 10'h131 == r_count_16_io_out ? io_r_305_b : _GEN_12394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12396 = 10'h132 == r_count_16_io_out ? io_r_306_b : _GEN_12395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12397 = 10'h133 == r_count_16_io_out ? io_r_307_b : _GEN_12396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12398 = 10'h134 == r_count_16_io_out ? io_r_308_b : _GEN_12397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12399 = 10'h135 == r_count_16_io_out ? io_r_309_b : _GEN_12398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12400 = 10'h136 == r_count_16_io_out ? io_r_310_b : _GEN_12399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12401 = 10'h137 == r_count_16_io_out ? io_r_311_b : _GEN_12400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12402 = 10'h138 == r_count_16_io_out ? io_r_312_b : _GEN_12401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12403 = 10'h139 == r_count_16_io_out ? io_r_313_b : _GEN_12402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12404 = 10'h13a == r_count_16_io_out ? io_r_314_b : _GEN_12403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12405 = 10'h13b == r_count_16_io_out ? io_r_315_b : _GEN_12404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12406 = 10'h13c == r_count_16_io_out ? io_r_316_b : _GEN_12405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12407 = 10'h13d == r_count_16_io_out ? io_r_317_b : _GEN_12406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12408 = 10'h13e == r_count_16_io_out ? io_r_318_b : _GEN_12407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12409 = 10'h13f == r_count_16_io_out ? io_r_319_b : _GEN_12408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12410 = 10'h140 == r_count_16_io_out ? io_r_320_b : _GEN_12409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12411 = 10'h141 == r_count_16_io_out ? io_r_321_b : _GEN_12410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12412 = 10'h142 == r_count_16_io_out ? io_r_322_b : _GEN_12411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12413 = 10'h143 == r_count_16_io_out ? io_r_323_b : _GEN_12412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12414 = 10'h144 == r_count_16_io_out ? io_r_324_b : _GEN_12413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12415 = 10'h145 == r_count_16_io_out ? io_r_325_b : _GEN_12414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12416 = 10'h146 == r_count_16_io_out ? io_r_326_b : _GEN_12415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12417 = 10'h147 == r_count_16_io_out ? io_r_327_b : _GEN_12416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12418 = 10'h148 == r_count_16_io_out ? io_r_328_b : _GEN_12417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12419 = 10'h149 == r_count_16_io_out ? io_r_329_b : _GEN_12418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12420 = 10'h14a == r_count_16_io_out ? io_r_330_b : _GEN_12419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12421 = 10'h14b == r_count_16_io_out ? io_r_331_b : _GEN_12420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12422 = 10'h14c == r_count_16_io_out ? io_r_332_b : _GEN_12421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12423 = 10'h14d == r_count_16_io_out ? io_r_333_b : _GEN_12422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12424 = 10'h14e == r_count_16_io_out ? io_r_334_b : _GEN_12423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12425 = 10'h14f == r_count_16_io_out ? io_r_335_b : _GEN_12424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12426 = 10'h150 == r_count_16_io_out ? io_r_336_b : _GEN_12425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12427 = 10'h151 == r_count_16_io_out ? io_r_337_b : _GEN_12426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12428 = 10'h152 == r_count_16_io_out ? io_r_338_b : _GEN_12427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12429 = 10'h153 == r_count_16_io_out ? io_r_339_b : _GEN_12428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12430 = 10'h154 == r_count_16_io_out ? io_r_340_b : _GEN_12429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12431 = 10'h155 == r_count_16_io_out ? io_r_341_b : _GEN_12430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12432 = 10'h156 == r_count_16_io_out ? io_r_342_b : _GEN_12431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12433 = 10'h157 == r_count_16_io_out ? io_r_343_b : _GEN_12432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12434 = 10'h158 == r_count_16_io_out ? io_r_344_b : _GEN_12433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12435 = 10'h159 == r_count_16_io_out ? io_r_345_b : _GEN_12434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12436 = 10'h15a == r_count_16_io_out ? io_r_346_b : _GEN_12435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12437 = 10'h15b == r_count_16_io_out ? io_r_347_b : _GEN_12436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12438 = 10'h15c == r_count_16_io_out ? io_r_348_b : _GEN_12437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12439 = 10'h15d == r_count_16_io_out ? io_r_349_b : _GEN_12438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12440 = 10'h15e == r_count_16_io_out ? io_r_350_b : _GEN_12439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12441 = 10'h15f == r_count_16_io_out ? io_r_351_b : _GEN_12440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12442 = 10'h160 == r_count_16_io_out ? io_r_352_b : _GEN_12441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12443 = 10'h161 == r_count_16_io_out ? io_r_353_b : _GEN_12442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12444 = 10'h162 == r_count_16_io_out ? io_r_354_b : _GEN_12443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12445 = 10'h163 == r_count_16_io_out ? io_r_355_b : _GEN_12444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12446 = 10'h164 == r_count_16_io_out ? io_r_356_b : _GEN_12445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12447 = 10'h165 == r_count_16_io_out ? io_r_357_b : _GEN_12446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12448 = 10'h166 == r_count_16_io_out ? io_r_358_b : _GEN_12447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12449 = 10'h167 == r_count_16_io_out ? io_r_359_b : _GEN_12448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12450 = 10'h168 == r_count_16_io_out ? io_r_360_b : _GEN_12449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12451 = 10'h169 == r_count_16_io_out ? io_r_361_b : _GEN_12450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12452 = 10'h16a == r_count_16_io_out ? io_r_362_b : _GEN_12451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12453 = 10'h16b == r_count_16_io_out ? io_r_363_b : _GEN_12452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12454 = 10'h16c == r_count_16_io_out ? io_r_364_b : _GEN_12453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12455 = 10'h16d == r_count_16_io_out ? io_r_365_b : _GEN_12454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12456 = 10'h16e == r_count_16_io_out ? io_r_366_b : _GEN_12455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12457 = 10'h16f == r_count_16_io_out ? io_r_367_b : _GEN_12456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12458 = 10'h170 == r_count_16_io_out ? io_r_368_b : _GEN_12457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12459 = 10'h171 == r_count_16_io_out ? io_r_369_b : _GEN_12458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12460 = 10'h172 == r_count_16_io_out ? io_r_370_b : _GEN_12459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12461 = 10'h173 == r_count_16_io_out ? io_r_371_b : _GEN_12460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12462 = 10'h174 == r_count_16_io_out ? io_r_372_b : _GEN_12461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12463 = 10'h175 == r_count_16_io_out ? io_r_373_b : _GEN_12462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12464 = 10'h176 == r_count_16_io_out ? io_r_374_b : _GEN_12463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12465 = 10'h177 == r_count_16_io_out ? io_r_375_b : _GEN_12464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12466 = 10'h178 == r_count_16_io_out ? io_r_376_b : _GEN_12465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12467 = 10'h179 == r_count_16_io_out ? io_r_377_b : _GEN_12466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12468 = 10'h17a == r_count_16_io_out ? io_r_378_b : _GEN_12467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12469 = 10'h17b == r_count_16_io_out ? io_r_379_b : _GEN_12468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12470 = 10'h17c == r_count_16_io_out ? io_r_380_b : _GEN_12469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12471 = 10'h17d == r_count_16_io_out ? io_r_381_b : _GEN_12470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12472 = 10'h17e == r_count_16_io_out ? io_r_382_b : _GEN_12471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12473 = 10'h17f == r_count_16_io_out ? io_r_383_b : _GEN_12472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12474 = 10'h180 == r_count_16_io_out ? io_r_384_b : _GEN_12473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12475 = 10'h181 == r_count_16_io_out ? io_r_385_b : _GEN_12474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12476 = 10'h182 == r_count_16_io_out ? io_r_386_b : _GEN_12475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12477 = 10'h183 == r_count_16_io_out ? io_r_387_b : _GEN_12476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12478 = 10'h184 == r_count_16_io_out ? io_r_388_b : _GEN_12477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12479 = 10'h185 == r_count_16_io_out ? io_r_389_b : _GEN_12478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12480 = 10'h186 == r_count_16_io_out ? io_r_390_b : _GEN_12479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12481 = 10'h187 == r_count_16_io_out ? io_r_391_b : _GEN_12480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12482 = 10'h188 == r_count_16_io_out ? io_r_392_b : _GEN_12481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12483 = 10'h189 == r_count_16_io_out ? io_r_393_b : _GEN_12482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12484 = 10'h18a == r_count_16_io_out ? io_r_394_b : _GEN_12483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12485 = 10'h18b == r_count_16_io_out ? io_r_395_b : _GEN_12484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12486 = 10'h18c == r_count_16_io_out ? io_r_396_b : _GEN_12485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12487 = 10'h18d == r_count_16_io_out ? io_r_397_b : _GEN_12486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12488 = 10'h18e == r_count_16_io_out ? io_r_398_b : _GEN_12487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12489 = 10'h18f == r_count_16_io_out ? io_r_399_b : _GEN_12488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12490 = 10'h190 == r_count_16_io_out ? io_r_400_b : _GEN_12489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12491 = 10'h191 == r_count_16_io_out ? io_r_401_b : _GEN_12490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12492 = 10'h192 == r_count_16_io_out ? io_r_402_b : _GEN_12491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12493 = 10'h193 == r_count_16_io_out ? io_r_403_b : _GEN_12492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12494 = 10'h194 == r_count_16_io_out ? io_r_404_b : _GEN_12493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12495 = 10'h195 == r_count_16_io_out ? io_r_405_b : _GEN_12494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12496 = 10'h196 == r_count_16_io_out ? io_r_406_b : _GEN_12495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12497 = 10'h197 == r_count_16_io_out ? io_r_407_b : _GEN_12496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12498 = 10'h198 == r_count_16_io_out ? io_r_408_b : _GEN_12497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12499 = 10'h199 == r_count_16_io_out ? io_r_409_b : _GEN_12498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12500 = 10'h19a == r_count_16_io_out ? io_r_410_b : _GEN_12499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12501 = 10'h19b == r_count_16_io_out ? io_r_411_b : _GEN_12500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12502 = 10'h19c == r_count_16_io_out ? io_r_412_b : _GEN_12501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12503 = 10'h19d == r_count_16_io_out ? io_r_413_b : _GEN_12502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12504 = 10'h19e == r_count_16_io_out ? io_r_414_b : _GEN_12503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12505 = 10'h19f == r_count_16_io_out ? io_r_415_b : _GEN_12504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12506 = 10'h1a0 == r_count_16_io_out ? io_r_416_b : _GEN_12505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12507 = 10'h1a1 == r_count_16_io_out ? io_r_417_b : _GEN_12506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12508 = 10'h1a2 == r_count_16_io_out ? io_r_418_b : _GEN_12507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12509 = 10'h1a3 == r_count_16_io_out ? io_r_419_b : _GEN_12508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12510 = 10'h1a4 == r_count_16_io_out ? io_r_420_b : _GEN_12509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12511 = 10'h1a5 == r_count_16_io_out ? io_r_421_b : _GEN_12510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12512 = 10'h1a6 == r_count_16_io_out ? io_r_422_b : _GEN_12511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12513 = 10'h1a7 == r_count_16_io_out ? io_r_423_b : _GEN_12512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12514 = 10'h1a8 == r_count_16_io_out ? io_r_424_b : _GEN_12513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12515 = 10'h1a9 == r_count_16_io_out ? io_r_425_b : _GEN_12514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12516 = 10'h1aa == r_count_16_io_out ? io_r_426_b : _GEN_12515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12517 = 10'h1ab == r_count_16_io_out ? io_r_427_b : _GEN_12516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12518 = 10'h1ac == r_count_16_io_out ? io_r_428_b : _GEN_12517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12519 = 10'h1ad == r_count_16_io_out ? io_r_429_b : _GEN_12518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12520 = 10'h1ae == r_count_16_io_out ? io_r_430_b : _GEN_12519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12521 = 10'h1af == r_count_16_io_out ? io_r_431_b : _GEN_12520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12522 = 10'h1b0 == r_count_16_io_out ? io_r_432_b : _GEN_12521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12523 = 10'h1b1 == r_count_16_io_out ? io_r_433_b : _GEN_12522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12524 = 10'h1b2 == r_count_16_io_out ? io_r_434_b : _GEN_12523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12525 = 10'h1b3 == r_count_16_io_out ? io_r_435_b : _GEN_12524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12526 = 10'h1b4 == r_count_16_io_out ? io_r_436_b : _GEN_12525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12527 = 10'h1b5 == r_count_16_io_out ? io_r_437_b : _GEN_12526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12528 = 10'h1b6 == r_count_16_io_out ? io_r_438_b : _GEN_12527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12529 = 10'h1b7 == r_count_16_io_out ? io_r_439_b : _GEN_12528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12530 = 10'h1b8 == r_count_16_io_out ? io_r_440_b : _GEN_12529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12531 = 10'h1b9 == r_count_16_io_out ? io_r_441_b : _GEN_12530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12532 = 10'h1ba == r_count_16_io_out ? io_r_442_b : _GEN_12531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12533 = 10'h1bb == r_count_16_io_out ? io_r_443_b : _GEN_12532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12534 = 10'h1bc == r_count_16_io_out ? io_r_444_b : _GEN_12533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12535 = 10'h1bd == r_count_16_io_out ? io_r_445_b : _GEN_12534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12536 = 10'h1be == r_count_16_io_out ? io_r_446_b : _GEN_12535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12537 = 10'h1bf == r_count_16_io_out ? io_r_447_b : _GEN_12536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12538 = 10'h1c0 == r_count_16_io_out ? io_r_448_b : _GEN_12537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12539 = 10'h1c1 == r_count_16_io_out ? io_r_449_b : _GEN_12538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12540 = 10'h1c2 == r_count_16_io_out ? io_r_450_b : _GEN_12539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12541 = 10'h1c3 == r_count_16_io_out ? io_r_451_b : _GEN_12540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12542 = 10'h1c4 == r_count_16_io_out ? io_r_452_b : _GEN_12541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12543 = 10'h1c5 == r_count_16_io_out ? io_r_453_b : _GEN_12542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12544 = 10'h1c6 == r_count_16_io_out ? io_r_454_b : _GEN_12543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12545 = 10'h1c7 == r_count_16_io_out ? io_r_455_b : _GEN_12544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12546 = 10'h1c8 == r_count_16_io_out ? io_r_456_b : _GEN_12545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12547 = 10'h1c9 == r_count_16_io_out ? io_r_457_b : _GEN_12546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12548 = 10'h1ca == r_count_16_io_out ? io_r_458_b : _GEN_12547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12549 = 10'h1cb == r_count_16_io_out ? io_r_459_b : _GEN_12548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12550 = 10'h1cc == r_count_16_io_out ? io_r_460_b : _GEN_12549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12551 = 10'h1cd == r_count_16_io_out ? io_r_461_b : _GEN_12550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12552 = 10'h1ce == r_count_16_io_out ? io_r_462_b : _GEN_12551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12553 = 10'h1cf == r_count_16_io_out ? io_r_463_b : _GEN_12552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12554 = 10'h1d0 == r_count_16_io_out ? io_r_464_b : _GEN_12553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12555 = 10'h1d1 == r_count_16_io_out ? io_r_465_b : _GEN_12554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12556 = 10'h1d2 == r_count_16_io_out ? io_r_466_b : _GEN_12555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12557 = 10'h1d3 == r_count_16_io_out ? io_r_467_b : _GEN_12556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12558 = 10'h1d4 == r_count_16_io_out ? io_r_468_b : _GEN_12557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12559 = 10'h1d5 == r_count_16_io_out ? io_r_469_b : _GEN_12558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12560 = 10'h1d6 == r_count_16_io_out ? io_r_470_b : _GEN_12559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12561 = 10'h1d7 == r_count_16_io_out ? io_r_471_b : _GEN_12560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12562 = 10'h1d8 == r_count_16_io_out ? io_r_472_b : _GEN_12561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12563 = 10'h1d9 == r_count_16_io_out ? io_r_473_b : _GEN_12562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12564 = 10'h1da == r_count_16_io_out ? io_r_474_b : _GEN_12563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12565 = 10'h1db == r_count_16_io_out ? io_r_475_b : _GEN_12564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12566 = 10'h1dc == r_count_16_io_out ? io_r_476_b : _GEN_12565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12567 = 10'h1dd == r_count_16_io_out ? io_r_477_b : _GEN_12566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12568 = 10'h1de == r_count_16_io_out ? io_r_478_b : _GEN_12567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12569 = 10'h1df == r_count_16_io_out ? io_r_479_b : _GEN_12568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12570 = 10'h1e0 == r_count_16_io_out ? io_r_480_b : _GEN_12569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12571 = 10'h1e1 == r_count_16_io_out ? io_r_481_b : _GEN_12570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12572 = 10'h1e2 == r_count_16_io_out ? io_r_482_b : _GEN_12571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12573 = 10'h1e3 == r_count_16_io_out ? io_r_483_b : _GEN_12572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12574 = 10'h1e4 == r_count_16_io_out ? io_r_484_b : _GEN_12573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12575 = 10'h1e5 == r_count_16_io_out ? io_r_485_b : _GEN_12574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12576 = 10'h1e6 == r_count_16_io_out ? io_r_486_b : _GEN_12575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12577 = 10'h1e7 == r_count_16_io_out ? io_r_487_b : _GEN_12576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12578 = 10'h1e8 == r_count_16_io_out ? io_r_488_b : _GEN_12577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12579 = 10'h1e9 == r_count_16_io_out ? io_r_489_b : _GEN_12578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12580 = 10'h1ea == r_count_16_io_out ? io_r_490_b : _GEN_12579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12581 = 10'h1eb == r_count_16_io_out ? io_r_491_b : _GEN_12580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12582 = 10'h1ec == r_count_16_io_out ? io_r_492_b : _GEN_12581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12583 = 10'h1ed == r_count_16_io_out ? io_r_493_b : _GEN_12582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12584 = 10'h1ee == r_count_16_io_out ? io_r_494_b : _GEN_12583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12585 = 10'h1ef == r_count_16_io_out ? io_r_495_b : _GEN_12584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12586 = 10'h1f0 == r_count_16_io_out ? io_r_496_b : _GEN_12585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12587 = 10'h1f1 == r_count_16_io_out ? io_r_497_b : _GEN_12586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12588 = 10'h1f2 == r_count_16_io_out ? io_r_498_b : _GEN_12587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12589 = 10'h1f3 == r_count_16_io_out ? io_r_499_b : _GEN_12588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12590 = 10'h1f4 == r_count_16_io_out ? io_r_500_b : _GEN_12589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12591 = 10'h1f5 == r_count_16_io_out ? io_r_501_b : _GEN_12590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12592 = 10'h1f6 == r_count_16_io_out ? io_r_502_b : _GEN_12591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12593 = 10'h1f7 == r_count_16_io_out ? io_r_503_b : _GEN_12592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12594 = 10'h1f8 == r_count_16_io_out ? io_r_504_b : _GEN_12593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12595 = 10'h1f9 == r_count_16_io_out ? io_r_505_b : _GEN_12594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12596 = 10'h1fa == r_count_16_io_out ? io_r_506_b : _GEN_12595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12597 = 10'h1fb == r_count_16_io_out ? io_r_507_b : _GEN_12596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12598 = 10'h1fc == r_count_16_io_out ? io_r_508_b : _GEN_12597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12599 = 10'h1fd == r_count_16_io_out ? io_r_509_b : _GEN_12598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12600 = 10'h1fe == r_count_16_io_out ? io_r_510_b : _GEN_12599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12601 = 10'h1ff == r_count_16_io_out ? io_r_511_b : _GEN_12600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12602 = 10'h200 == r_count_16_io_out ? io_r_512_b : _GEN_12601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12603 = 10'h201 == r_count_16_io_out ? io_r_513_b : _GEN_12602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12604 = 10'h202 == r_count_16_io_out ? io_r_514_b : _GEN_12603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12605 = 10'h203 == r_count_16_io_out ? io_r_515_b : _GEN_12604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12606 = 10'h204 == r_count_16_io_out ? io_r_516_b : _GEN_12605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12607 = 10'h205 == r_count_16_io_out ? io_r_517_b : _GEN_12606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12608 = 10'h206 == r_count_16_io_out ? io_r_518_b : _GEN_12607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12609 = 10'h207 == r_count_16_io_out ? io_r_519_b : _GEN_12608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12610 = 10'h208 == r_count_16_io_out ? io_r_520_b : _GEN_12609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12611 = 10'h209 == r_count_16_io_out ? io_r_521_b : _GEN_12610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12612 = 10'h20a == r_count_16_io_out ? io_r_522_b : _GEN_12611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12613 = 10'h20b == r_count_16_io_out ? io_r_523_b : _GEN_12612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12614 = 10'h20c == r_count_16_io_out ? io_r_524_b : _GEN_12613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12615 = 10'h20d == r_count_16_io_out ? io_r_525_b : _GEN_12614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12616 = 10'h20e == r_count_16_io_out ? io_r_526_b : _GEN_12615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12617 = 10'h20f == r_count_16_io_out ? io_r_527_b : _GEN_12616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12618 = 10'h210 == r_count_16_io_out ? io_r_528_b : _GEN_12617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12619 = 10'h211 == r_count_16_io_out ? io_r_529_b : _GEN_12618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12620 = 10'h212 == r_count_16_io_out ? io_r_530_b : _GEN_12619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12621 = 10'h213 == r_count_16_io_out ? io_r_531_b : _GEN_12620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12622 = 10'h214 == r_count_16_io_out ? io_r_532_b : _GEN_12621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12623 = 10'h215 == r_count_16_io_out ? io_r_533_b : _GEN_12622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12624 = 10'h216 == r_count_16_io_out ? io_r_534_b : _GEN_12623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12625 = 10'h217 == r_count_16_io_out ? io_r_535_b : _GEN_12624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12626 = 10'h218 == r_count_16_io_out ? io_r_536_b : _GEN_12625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12627 = 10'h219 == r_count_16_io_out ? io_r_537_b : _GEN_12626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12628 = 10'h21a == r_count_16_io_out ? io_r_538_b : _GEN_12627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12629 = 10'h21b == r_count_16_io_out ? io_r_539_b : _GEN_12628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12630 = 10'h21c == r_count_16_io_out ? io_r_540_b : _GEN_12629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12631 = 10'h21d == r_count_16_io_out ? io_r_541_b : _GEN_12630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12632 = 10'h21e == r_count_16_io_out ? io_r_542_b : _GEN_12631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12633 = 10'h21f == r_count_16_io_out ? io_r_543_b : _GEN_12632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12634 = 10'h220 == r_count_16_io_out ? io_r_544_b : _GEN_12633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12635 = 10'h221 == r_count_16_io_out ? io_r_545_b : _GEN_12634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12636 = 10'h222 == r_count_16_io_out ? io_r_546_b : _GEN_12635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12637 = 10'h223 == r_count_16_io_out ? io_r_547_b : _GEN_12636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12638 = 10'h224 == r_count_16_io_out ? io_r_548_b : _GEN_12637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12639 = 10'h225 == r_count_16_io_out ? io_r_549_b : _GEN_12638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12640 = 10'h226 == r_count_16_io_out ? io_r_550_b : _GEN_12639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12641 = 10'h227 == r_count_16_io_out ? io_r_551_b : _GEN_12640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12642 = 10'h228 == r_count_16_io_out ? io_r_552_b : _GEN_12641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12643 = 10'h229 == r_count_16_io_out ? io_r_553_b : _GEN_12642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12644 = 10'h22a == r_count_16_io_out ? io_r_554_b : _GEN_12643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12645 = 10'h22b == r_count_16_io_out ? io_r_555_b : _GEN_12644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12646 = 10'h22c == r_count_16_io_out ? io_r_556_b : _GEN_12645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12647 = 10'h22d == r_count_16_io_out ? io_r_557_b : _GEN_12646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12648 = 10'h22e == r_count_16_io_out ? io_r_558_b : _GEN_12647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12649 = 10'h22f == r_count_16_io_out ? io_r_559_b : _GEN_12648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12650 = 10'h230 == r_count_16_io_out ? io_r_560_b : _GEN_12649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12651 = 10'h231 == r_count_16_io_out ? io_r_561_b : _GEN_12650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12652 = 10'h232 == r_count_16_io_out ? io_r_562_b : _GEN_12651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12653 = 10'h233 == r_count_16_io_out ? io_r_563_b : _GEN_12652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12654 = 10'h234 == r_count_16_io_out ? io_r_564_b : _GEN_12653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12655 = 10'h235 == r_count_16_io_out ? io_r_565_b : _GEN_12654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12656 = 10'h236 == r_count_16_io_out ? io_r_566_b : _GEN_12655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12657 = 10'h237 == r_count_16_io_out ? io_r_567_b : _GEN_12656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12658 = 10'h238 == r_count_16_io_out ? io_r_568_b : _GEN_12657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12659 = 10'h239 == r_count_16_io_out ? io_r_569_b : _GEN_12658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12660 = 10'h23a == r_count_16_io_out ? io_r_570_b : _GEN_12659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12661 = 10'h23b == r_count_16_io_out ? io_r_571_b : _GEN_12660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12662 = 10'h23c == r_count_16_io_out ? io_r_572_b : _GEN_12661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12663 = 10'h23d == r_count_16_io_out ? io_r_573_b : _GEN_12662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12664 = 10'h23e == r_count_16_io_out ? io_r_574_b : _GEN_12663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12665 = 10'h23f == r_count_16_io_out ? io_r_575_b : _GEN_12664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12666 = 10'h240 == r_count_16_io_out ? io_r_576_b : _GEN_12665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12667 = 10'h241 == r_count_16_io_out ? io_r_577_b : _GEN_12666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12668 = 10'h242 == r_count_16_io_out ? io_r_578_b : _GEN_12667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12669 = 10'h243 == r_count_16_io_out ? io_r_579_b : _GEN_12668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12670 = 10'h244 == r_count_16_io_out ? io_r_580_b : _GEN_12669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12671 = 10'h245 == r_count_16_io_out ? io_r_581_b : _GEN_12670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12672 = 10'h246 == r_count_16_io_out ? io_r_582_b : _GEN_12671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12673 = 10'h247 == r_count_16_io_out ? io_r_583_b : _GEN_12672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12674 = 10'h248 == r_count_16_io_out ? io_r_584_b : _GEN_12673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12675 = 10'h249 == r_count_16_io_out ? io_r_585_b : _GEN_12674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12676 = 10'h24a == r_count_16_io_out ? io_r_586_b : _GEN_12675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12677 = 10'h24b == r_count_16_io_out ? io_r_587_b : _GEN_12676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12678 = 10'h24c == r_count_16_io_out ? io_r_588_b : _GEN_12677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12679 = 10'h24d == r_count_16_io_out ? io_r_589_b : _GEN_12678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12680 = 10'h24e == r_count_16_io_out ? io_r_590_b : _GEN_12679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12681 = 10'h24f == r_count_16_io_out ? io_r_591_b : _GEN_12680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12682 = 10'h250 == r_count_16_io_out ? io_r_592_b : _GEN_12681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12683 = 10'h251 == r_count_16_io_out ? io_r_593_b : _GEN_12682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12684 = 10'h252 == r_count_16_io_out ? io_r_594_b : _GEN_12683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12685 = 10'h253 == r_count_16_io_out ? io_r_595_b : _GEN_12684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12686 = 10'h254 == r_count_16_io_out ? io_r_596_b : _GEN_12685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12687 = 10'h255 == r_count_16_io_out ? io_r_597_b : _GEN_12686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12688 = 10'h256 == r_count_16_io_out ? io_r_598_b : _GEN_12687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12689 = 10'h257 == r_count_16_io_out ? io_r_599_b : _GEN_12688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12690 = 10'h258 == r_count_16_io_out ? io_r_600_b : _GEN_12689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12691 = 10'h259 == r_count_16_io_out ? io_r_601_b : _GEN_12690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12692 = 10'h25a == r_count_16_io_out ? io_r_602_b : _GEN_12691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12693 = 10'h25b == r_count_16_io_out ? io_r_603_b : _GEN_12692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12694 = 10'h25c == r_count_16_io_out ? io_r_604_b : _GEN_12693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12695 = 10'h25d == r_count_16_io_out ? io_r_605_b : _GEN_12694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12696 = 10'h25e == r_count_16_io_out ? io_r_606_b : _GEN_12695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12697 = 10'h25f == r_count_16_io_out ? io_r_607_b : _GEN_12696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12698 = 10'h260 == r_count_16_io_out ? io_r_608_b : _GEN_12697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12699 = 10'h261 == r_count_16_io_out ? io_r_609_b : _GEN_12698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12700 = 10'h262 == r_count_16_io_out ? io_r_610_b : _GEN_12699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12701 = 10'h263 == r_count_16_io_out ? io_r_611_b : _GEN_12700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12702 = 10'h264 == r_count_16_io_out ? io_r_612_b : _GEN_12701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12703 = 10'h265 == r_count_16_io_out ? io_r_613_b : _GEN_12702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12704 = 10'h266 == r_count_16_io_out ? io_r_614_b : _GEN_12703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12705 = 10'h267 == r_count_16_io_out ? io_r_615_b : _GEN_12704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12706 = 10'h268 == r_count_16_io_out ? io_r_616_b : _GEN_12705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12707 = 10'h269 == r_count_16_io_out ? io_r_617_b : _GEN_12706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12708 = 10'h26a == r_count_16_io_out ? io_r_618_b : _GEN_12707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12709 = 10'h26b == r_count_16_io_out ? io_r_619_b : _GEN_12708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12710 = 10'h26c == r_count_16_io_out ? io_r_620_b : _GEN_12709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12711 = 10'h26d == r_count_16_io_out ? io_r_621_b : _GEN_12710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12712 = 10'h26e == r_count_16_io_out ? io_r_622_b : _GEN_12711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12713 = 10'h26f == r_count_16_io_out ? io_r_623_b : _GEN_12712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12714 = 10'h270 == r_count_16_io_out ? io_r_624_b : _GEN_12713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12715 = 10'h271 == r_count_16_io_out ? io_r_625_b : _GEN_12714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12716 = 10'h272 == r_count_16_io_out ? io_r_626_b : _GEN_12715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12717 = 10'h273 == r_count_16_io_out ? io_r_627_b : _GEN_12716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12718 = 10'h274 == r_count_16_io_out ? io_r_628_b : _GEN_12717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12719 = 10'h275 == r_count_16_io_out ? io_r_629_b : _GEN_12718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12720 = 10'h276 == r_count_16_io_out ? io_r_630_b : _GEN_12719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12721 = 10'h277 == r_count_16_io_out ? io_r_631_b : _GEN_12720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12722 = 10'h278 == r_count_16_io_out ? io_r_632_b : _GEN_12721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12723 = 10'h279 == r_count_16_io_out ? io_r_633_b : _GEN_12722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12724 = 10'h27a == r_count_16_io_out ? io_r_634_b : _GEN_12723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12725 = 10'h27b == r_count_16_io_out ? io_r_635_b : _GEN_12724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12726 = 10'h27c == r_count_16_io_out ? io_r_636_b : _GEN_12725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12727 = 10'h27d == r_count_16_io_out ? io_r_637_b : _GEN_12726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12728 = 10'h27e == r_count_16_io_out ? io_r_638_b : _GEN_12727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12729 = 10'h27f == r_count_16_io_out ? io_r_639_b : _GEN_12728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12730 = 10'h280 == r_count_16_io_out ? io_r_640_b : _GEN_12729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12731 = 10'h281 == r_count_16_io_out ? io_r_641_b : _GEN_12730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12732 = 10'h282 == r_count_16_io_out ? io_r_642_b : _GEN_12731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12733 = 10'h283 == r_count_16_io_out ? io_r_643_b : _GEN_12732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12734 = 10'h284 == r_count_16_io_out ? io_r_644_b : _GEN_12733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12735 = 10'h285 == r_count_16_io_out ? io_r_645_b : _GEN_12734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12736 = 10'h286 == r_count_16_io_out ? io_r_646_b : _GEN_12735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12737 = 10'h287 == r_count_16_io_out ? io_r_647_b : _GEN_12736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12738 = 10'h288 == r_count_16_io_out ? io_r_648_b : _GEN_12737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12739 = 10'h289 == r_count_16_io_out ? io_r_649_b : _GEN_12738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12740 = 10'h28a == r_count_16_io_out ? io_r_650_b : _GEN_12739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12741 = 10'h28b == r_count_16_io_out ? io_r_651_b : _GEN_12740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12742 = 10'h28c == r_count_16_io_out ? io_r_652_b : _GEN_12741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12743 = 10'h28d == r_count_16_io_out ? io_r_653_b : _GEN_12742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12744 = 10'h28e == r_count_16_io_out ? io_r_654_b : _GEN_12743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12745 = 10'h28f == r_count_16_io_out ? io_r_655_b : _GEN_12744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12746 = 10'h290 == r_count_16_io_out ? io_r_656_b : _GEN_12745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12747 = 10'h291 == r_count_16_io_out ? io_r_657_b : _GEN_12746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12748 = 10'h292 == r_count_16_io_out ? io_r_658_b : _GEN_12747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12749 = 10'h293 == r_count_16_io_out ? io_r_659_b : _GEN_12748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12750 = 10'h294 == r_count_16_io_out ? io_r_660_b : _GEN_12749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12751 = 10'h295 == r_count_16_io_out ? io_r_661_b : _GEN_12750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12752 = 10'h296 == r_count_16_io_out ? io_r_662_b : _GEN_12751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12753 = 10'h297 == r_count_16_io_out ? io_r_663_b : _GEN_12752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12754 = 10'h298 == r_count_16_io_out ? io_r_664_b : _GEN_12753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12755 = 10'h299 == r_count_16_io_out ? io_r_665_b : _GEN_12754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12756 = 10'h29a == r_count_16_io_out ? io_r_666_b : _GEN_12755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12757 = 10'h29b == r_count_16_io_out ? io_r_667_b : _GEN_12756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12758 = 10'h29c == r_count_16_io_out ? io_r_668_b : _GEN_12757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12759 = 10'h29d == r_count_16_io_out ? io_r_669_b : _GEN_12758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12760 = 10'h29e == r_count_16_io_out ? io_r_670_b : _GEN_12759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12761 = 10'h29f == r_count_16_io_out ? io_r_671_b : _GEN_12760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12762 = 10'h2a0 == r_count_16_io_out ? io_r_672_b : _GEN_12761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12763 = 10'h2a1 == r_count_16_io_out ? io_r_673_b : _GEN_12762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12764 = 10'h2a2 == r_count_16_io_out ? io_r_674_b : _GEN_12763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12765 = 10'h2a3 == r_count_16_io_out ? io_r_675_b : _GEN_12764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12766 = 10'h2a4 == r_count_16_io_out ? io_r_676_b : _GEN_12765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12767 = 10'h2a5 == r_count_16_io_out ? io_r_677_b : _GEN_12766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12768 = 10'h2a6 == r_count_16_io_out ? io_r_678_b : _GEN_12767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12769 = 10'h2a7 == r_count_16_io_out ? io_r_679_b : _GEN_12768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12770 = 10'h2a8 == r_count_16_io_out ? io_r_680_b : _GEN_12769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12771 = 10'h2a9 == r_count_16_io_out ? io_r_681_b : _GEN_12770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12772 = 10'h2aa == r_count_16_io_out ? io_r_682_b : _GEN_12771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12773 = 10'h2ab == r_count_16_io_out ? io_r_683_b : _GEN_12772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12774 = 10'h2ac == r_count_16_io_out ? io_r_684_b : _GEN_12773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12775 = 10'h2ad == r_count_16_io_out ? io_r_685_b : _GEN_12774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12776 = 10'h2ae == r_count_16_io_out ? io_r_686_b : _GEN_12775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12777 = 10'h2af == r_count_16_io_out ? io_r_687_b : _GEN_12776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12778 = 10'h2b0 == r_count_16_io_out ? io_r_688_b : _GEN_12777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12779 = 10'h2b1 == r_count_16_io_out ? io_r_689_b : _GEN_12778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12780 = 10'h2b2 == r_count_16_io_out ? io_r_690_b : _GEN_12779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12781 = 10'h2b3 == r_count_16_io_out ? io_r_691_b : _GEN_12780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12782 = 10'h2b4 == r_count_16_io_out ? io_r_692_b : _GEN_12781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12783 = 10'h2b5 == r_count_16_io_out ? io_r_693_b : _GEN_12782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12784 = 10'h2b6 == r_count_16_io_out ? io_r_694_b : _GEN_12783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12785 = 10'h2b7 == r_count_16_io_out ? io_r_695_b : _GEN_12784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12786 = 10'h2b8 == r_count_16_io_out ? io_r_696_b : _GEN_12785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12787 = 10'h2b9 == r_count_16_io_out ? io_r_697_b : _GEN_12786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12788 = 10'h2ba == r_count_16_io_out ? io_r_698_b : _GEN_12787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12789 = 10'h2bb == r_count_16_io_out ? io_r_699_b : _GEN_12788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12790 = 10'h2bc == r_count_16_io_out ? io_r_700_b : _GEN_12789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12791 = 10'h2bd == r_count_16_io_out ? io_r_701_b : _GEN_12790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12792 = 10'h2be == r_count_16_io_out ? io_r_702_b : _GEN_12791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12793 = 10'h2bf == r_count_16_io_out ? io_r_703_b : _GEN_12792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12794 = 10'h2c0 == r_count_16_io_out ? io_r_704_b : _GEN_12793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12795 = 10'h2c1 == r_count_16_io_out ? io_r_705_b : _GEN_12794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12796 = 10'h2c2 == r_count_16_io_out ? io_r_706_b : _GEN_12795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12797 = 10'h2c3 == r_count_16_io_out ? io_r_707_b : _GEN_12796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12798 = 10'h2c4 == r_count_16_io_out ? io_r_708_b : _GEN_12797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12799 = 10'h2c5 == r_count_16_io_out ? io_r_709_b : _GEN_12798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12800 = 10'h2c6 == r_count_16_io_out ? io_r_710_b : _GEN_12799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12801 = 10'h2c7 == r_count_16_io_out ? io_r_711_b : _GEN_12800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12802 = 10'h2c8 == r_count_16_io_out ? io_r_712_b : _GEN_12801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12803 = 10'h2c9 == r_count_16_io_out ? io_r_713_b : _GEN_12802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12804 = 10'h2ca == r_count_16_io_out ? io_r_714_b : _GEN_12803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12805 = 10'h2cb == r_count_16_io_out ? io_r_715_b : _GEN_12804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12806 = 10'h2cc == r_count_16_io_out ? io_r_716_b : _GEN_12805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12807 = 10'h2cd == r_count_16_io_out ? io_r_717_b : _GEN_12806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12808 = 10'h2ce == r_count_16_io_out ? io_r_718_b : _GEN_12807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12809 = 10'h2cf == r_count_16_io_out ? io_r_719_b : _GEN_12808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12810 = 10'h2d0 == r_count_16_io_out ? io_r_720_b : _GEN_12809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12811 = 10'h2d1 == r_count_16_io_out ? io_r_721_b : _GEN_12810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12812 = 10'h2d2 == r_count_16_io_out ? io_r_722_b : _GEN_12811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12813 = 10'h2d3 == r_count_16_io_out ? io_r_723_b : _GEN_12812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12814 = 10'h2d4 == r_count_16_io_out ? io_r_724_b : _GEN_12813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12815 = 10'h2d5 == r_count_16_io_out ? io_r_725_b : _GEN_12814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12816 = 10'h2d6 == r_count_16_io_out ? io_r_726_b : _GEN_12815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12817 = 10'h2d7 == r_count_16_io_out ? io_r_727_b : _GEN_12816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12818 = 10'h2d8 == r_count_16_io_out ? io_r_728_b : _GEN_12817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12819 = 10'h2d9 == r_count_16_io_out ? io_r_729_b : _GEN_12818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12820 = 10'h2da == r_count_16_io_out ? io_r_730_b : _GEN_12819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12821 = 10'h2db == r_count_16_io_out ? io_r_731_b : _GEN_12820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12822 = 10'h2dc == r_count_16_io_out ? io_r_732_b : _GEN_12821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12823 = 10'h2dd == r_count_16_io_out ? io_r_733_b : _GEN_12822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12824 = 10'h2de == r_count_16_io_out ? io_r_734_b : _GEN_12823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12825 = 10'h2df == r_count_16_io_out ? io_r_735_b : _GEN_12824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12826 = 10'h2e0 == r_count_16_io_out ? io_r_736_b : _GEN_12825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12827 = 10'h2e1 == r_count_16_io_out ? io_r_737_b : _GEN_12826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12828 = 10'h2e2 == r_count_16_io_out ? io_r_738_b : _GEN_12827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12829 = 10'h2e3 == r_count_16_io_out ? io_r_739_b : _GEN_12828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12830 = 10'h2e4 == r_count_16_io_out ? io_r_740_b : _GEN_12829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12831 = 10'h2e5 == r_count_16_io_out ? io_r_741_b : _GEN_12830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12832 = 10'h2e6 == r_count_16_io_out ? io_r_742_b : _GEN_12831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12833 = 10'h2e7 == r_count_16_io_out ? io_r_743_b : _GEN_12832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12834 = 10'h2e8 == r_count_16_io_out ? io_r_744_b : _GEN_12833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12835 = 10'h2e9 == r_count_16_io_out ? io_r_745_b : _GEN_12834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12836 = 10'h2ea == r_count_16_io_out ? io_r_746_b : _GEN_12835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12837 = 10'h2eb == r_count_16_io_out ? io_r_747_b : _GEN_12836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12838 = 10'h2ec == r_count_16_io_out ? io_r_748_b : _GEN_12837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12841 = 10'h1 == r_count_17_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12842 = 10'h2 == r_count_17_io_out ? io_r_2_b : _GEN_12841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12843 = 10'h3 == r_count_17_io_out ? io_r_3_b : _GEN_12842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12844 = 10'h4 == r_count_17_io_out ? io_r_4_b : _GEN_12843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12845 = 10'h5 == r_count_17_io_out ? io_r_5_b : _GEN_12844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12846 = 10'h6 == r_count_17_io_out ? io_r_6_b : _GEN_12845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12847 = 10'h7 == r_count_17_io_out ? io_r_7_b : _GEN_12846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12848 = 10'h8 == r_count_17_io_out ? io_r_8_b : _GEN_12847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12849 = 10'h9 == r_count_17_io_out ? io_r_9_b : _GEN_12848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12850 = 10'ha == r_count_17_io_out ? io_r_10_b : _GEN_12849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12851 = 10'hb == r_count_17_io_out ? io_r_11_b : _GEN_12850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12852 = 10'hc == r_count_17_io_out ? io_r_12_b : _GEN_12851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12853 = 10'hd == r_count_17_io_out ? io_r_13_b : _GEN_12852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12854 = 10'he == r_count_17_io_out ? io_r_14_b : _GEN_12853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12855 = 10'hf == r_count_17_io_out ? io_r_15_b : _GEN_12854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12856 = 10'h10 == r_count_17_io_out ? io_r_16_b : _GEN_12855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12857 = 10'h11 == r_count_17_io_out ? io_r_17_b : _GEN_12856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12858 = 10'h12 == r_count_17_io_out ? io_r_18_b : _GEN_12857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12859 = 10'h13 == r_count_17_io_out ? io_r_19_b : _GEN_12858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12860 = 10'h14 == r_count_17_io_out ? io_r_20_b : _GEN_12859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12861 = 10'h15 == r_count_17_io_out ? io_r_21_b : _GEN_12860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12862 = 10'h16 == r_count_17_io_out ? io_r_22_b : _GEN_12861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12863 = 10'h17 == r_count_17_io_out ? io_r_23_b : _GEN_12862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12864 = 10'h18 == r_count_17_io_out ? io_r_24_b : _GEN_12863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12865 = 10'h19 == r_count_17_io_out ? io_r_25_b : _GEN_12864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12866 = 10'h1a == r_count_17_io_out ? io_r_26_b : _GEN_12865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12867 = 10'h1b == r_count_17_io_out ? io_r_27_b : _GEN_12866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12868 = 10'h1c == r_count_17_io_out ? io_r_28_b : _GEN_12867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12869 = 10'h1d == r_count_17_io_out ? io_r_29_b : _GEN_12868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12870 = 10'h1e == r_count_17_io_out ? io_r_30_b : _GEN_12869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12871 = 10'h1f == r_count_17_io_out ? io_r_31_b : _GEN_12870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12872 = 10'h20 == r_count_17_io_out ? io_r_32_b : _GEN_12871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12873 = 10'h21 == r_count_17_io_out ? io_r_33_b : _GEN_12872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12874 = 10'h22 == r_count_17_io_out ? io_r_34_b : _GEN_12873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12875 = 10'h23 == r_count_17_io_out ? io_r_35_b : _GEN_12874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12876 = 10'h24 == r_count_17_io_out ? io_r_36_b : _GEN_12875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12877 = 10'h25 == r_count_17_io_out ? io_r_37_b : _GEN_12876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12878 = 10'h26 == r_count_17_io_out ? io_r_38_b : _GEN_12877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12879 = 10'h27 == r_count_17_io_out ? io_r_39_b : _GEN_12878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12880 = 10'h28 == r_count_17_io_out ? io_r_40_b : _GEN_12879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12881 = 10'h29 == r_count_17_io_out ? io_r_41_b : _GEN_12880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12882 = 10'h2a == r_count_17_io_out ? io_r_42_b : _GEN_12881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12883 = 10'h2b == r_count_17_io_out ? io_r_43_b : _GEN_12882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12884 = 10'h2c == r_count_17_io_out ? io_r_44_b : _GEN_12883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12885 = 10'h2d == r_count_17_io_out ? io_r_45_b : _GEN_12884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12886 = 10'h2e == r_count_17_io_out ? io_r_46_b : _GEN_12885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12887 = 10'h2f == r_count_17_io_out ? io_r_47_b : _GEN_12886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12888 = 10'h30 == r_count_17_io_out ? io_r_48_b : _GEN_12887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12889 = 10'h31 == r_count_17_io_out ? io_r_49_b : _GEN_12888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12890 = 10'h32 == r_count_17_io_out ? io_r_50_b : _GEN_12889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12891 = 10'h33 == r_count_17_io_out ? io_r_51_b : _GEN_12890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12892 = 10'h34 == r_count_17_io_out ? io_r_52_b : _GEN_12891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12893 = 10'h35 == r_count_17_io_out ? io_r_53_b : _GEN_12892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12894 = 10'h36 == r_count_17_io_out ? io_r_54_b : _GEN_12893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12895 = 10'h37 == r_count_17_io_out ? io_r_55_b : _GEN_12894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12896 = 10'h38 == r_count_17_io_out ? io_r_56_b : _GEN_12895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12897 = 10'h39 == r_count_17_io_out ? io_r_57_b : _GEN_12896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12898 = 10'h3a == r_count_17_io_out ? io_r_58_b : _GEN_12897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12899 = 10'h3b == r_count_17_io_out ? io_r_59_b : _GEN_12898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12900 = 10'h3c == r_count_17_io_out ? io_r_60_b : _GEN_12899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12901 = 10'h3d == r_count_17_io_out ? io_r_61_b : _GEN_12900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12902 = 10'h3e == r_count_17_io_out ? io_r_62_b : _GEN_12901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12903 = 10'h3f == r_count_17_io_out ? io_r_63_b : _GEN_12902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12904 = 10'h40 == r_count_17_io_out ? io_r_64_b : _GEN_12903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12905 = 10'h41 == r_count_17_io_out ? io_r_65_b : _GEN_12904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12906 = 10'h42 == r_count_17_io_out ? io_r_66_b : _GEN_12905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12907 = 10'h43 == r_count_17_io_out ? io_r_67_b : _GEN_12906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12908 = 10'h44 == r_count_17_io_out ? io_r_68_b : _GEN_12907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12909 = 10'h45 == r_count_17_io_out ? io_r_69_b : _GEN_12908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12910 = 10'h46 == r_count_17_io_out ? io_r_70_b : _GEN_12909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12911 = 10'h47 == r_count_17_io_out ? io_r_71_b : _GEN_12910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12912 = 10'h48 == r_count_17_io_out ? io_r_72_b : _GEN_12911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12913 = 10'h49 == r_count_17_io_out ? io_r_73_b : _GEN_12912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12914 = 10'h4a == r_count_17_io_out ? io_r_74_b : _GEN_12913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12915 = 10'h4b == r_count_17_io_out ? io_r_75_b : _GEN_12914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12916 = 10'h4c == r_count_17_io_out ? io_r_76_b : _GEN_12915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12917 = 10'h4d == r_count_17_io_out ? io_r_77_b : _GEN_12916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12918 = 10'h4e == r_count_17_io_out ? io_r_78_b : _GEN_12917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12919 = 10'h4f == r_count_17_io_out ? io_r_79_b : _GEN_12918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12920 = 10'h50 == r_count_17_io_out ? io_r_80_b : _GEN_12919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12921 = 10'h51 == r_count_17_io_out ? io_r_81_b : _GEN_12920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12922 = 10'h52 == r_count_17_io_out ? io_r_82_b : _GEN_12921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12923 = 10'h53 == r_count_17_io_out ? io_r_83_b : _GEN_12922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12924 = 10'h54 == r_count_17_io_out ? io_r_84_b : _GEN_12923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12925 = 10'h55 == r_count_17_io_out ? io_r_85_b : _GEN_12924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12926 = 10'h56 == r_count_17_io_out ? io_r_86_b : _GEN_12925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12927 = 10'h57 == r_count_17_io_out ? io_r_87_b : _GEN_12926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12928 = 10'h58 == r_count_17_io_out ? io_r_88_b : _GEN_12927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12929 = 10'h59 == r_count_17_io_out ? io_r_89_b : _GEN_12928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12930 = 10'h5a == r_count_17_io_out ? io_r_90_b : _GEN_12929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12931 = 10'h5b == r_count_17_io_out ? io_r_91_b : _GEN_12930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12932 = 10'h5c == r_count_17_io_out ? io_r_92_b : _GEN_12931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12933 = 10'h5d == r_count_17_io_out ? io_r_93_b : _GEN_12932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12934 = 10'h5e == r_count_17_io_out ? io_r_94_b : _GEN_12933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12935 = 10'h5f == r_count_17_io_out ? io_r_95_b : _GEN_12934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12936 = 10'h60 == r_count_17_io_out ? io_r_96_b : _GEN_12935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12937 = 10'h61 == r_count_17_io_out ? io_r_97_b : _GEN_12936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12938 = 10'h62 == r_count_17_io_out ? io_r_98_b : _GEN_12937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12939 = 10'h63 == r_count_17_io_out ? io_r_99_b : _GEN_12938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12940 = 10'h64 == r_count_17_io_out ? io_r_100_b : _GEN_12939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12941 = 10'h65 == r_count_17_io_out ? io_r_101_b : _GEN_12940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12942 = 10'h66 == r_count_17_io_out ? io_r_102_b : _GEN_12941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12943 = 10'h67 == r_count_17_io_out ? io_r_103_b : _GEN_12942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12944 = 10'h68 == r_count_17_io_out ? io_r_104_b : _GEN_12943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12945 = 10'h69 == r_count_17_io_out ? io_r_105_b : _GEN_12944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12946 = 10'h6a == r_count_17_io_out ? io_r_106_b : _GEN_12945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12947 = 10'h6b == r_count_17_io_out ? io_r_107_b : _GEN_12946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12948 = 10'h6c == r_count_17_io_out ? io_r_108_b : _GEN_12947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12949 = 10'h6d == r_count_17_io_out ? io_r_109_b : _GEN_12948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12950 = 10'h6e == r_count_17_io_out ? io_r_110_b : _GEN_12949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12951 = 10'h6f == r_count_17_io_out ? io_r_111_b : _GEN_12950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12952 = 10'h70 == r_count_17_io_out ? io_r_112_b : _GEN_12951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12953 = 10'h71 == r_count_17_io_out ? io_r_113_b : _GEN_12952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12954 = 10'h72 == r_count_17_io_out ? io_r_114_b : _GEN_12953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12955 = 10'h73 == r_count_17_io_out ? io_r_115_b : _GEN_12954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12956 = 10'h74 == r_count_17_io_out ? io_r_116_b : _GEN_12955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12957 = 10'h75 == r_count_17_io_out ? io_r_117_b : _GEN_12956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12958 = 10'h76 == r_count_17_io_out ? io_r_118_b : _GEN_12957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12959 = 10'h77 == r_count_17_io_out ? io_r_119_b : _GEN_12958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12960 = 10'h78 == r_count_17_io_out ? io_r_120_b : _GEN_12959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12961 = 10'h79 == r_count_17_io_out ? io_r_121_b : _GEN_12960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12962 = 10'h7a == r_count_17_io_out ? io_r_122_b : _GEN_12961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12963 = 10'h7b == r_count_17_io_out ? io_r_123_b : _GEN_12962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12964 = 10'h7c == r_count_17_io_out ? io_r_124_b : _GEN_12963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12965 = 10'h7d == r_count_17_io_out ? io_r_125_b : _GEN_12964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12966 = 10'h7e == r_count_17_io_out ? io_r_126_b : _GEN_12965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12967 = 10'h7f == r_count_17_io_out ? io_r_127_b : _GEN_12966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12968 = 10'h80 == r_count_17_io_out ? io_r_128_b : _GEN_12967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12969 = 10'h81 == r_count_17_io_out ? io_r_129_b : _GEN_12968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12970 = 10'h82 == r_count_17_io_out ? io_r_130_b : _GEN_12969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12971 = 10'h83 == r_count_17_io_out ? io_r_131_b : _GEN_12970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12972 = 10'h84 == r_count_17_io_out ? io_r_132_b : _GEN_12971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12973 = 10'h85 == r_count_17_io_out ? io_r_133_b : _GEN_12972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12974 = 10'h86 == r_count_17_io_out ? io_r_134_b : _GEN_12973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12975 = 10'h87 == r_count_17_io_out ? io_r_135_b : _GEN_12974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12976 = 10'h88 == r_count_17_io_out ? io_r_136_b : _GEN_12975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12977 = 10'h89 == r_count_17_io_out ? io_r_137_b : _GEN_12976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12978 = 10'h8a == r_count_17_io_out ? io_r_138_b : _GEN_12977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12979 = 10'h8b == r_count_17_io_out ? io_r_139_b : _GEN_12978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12980 = 10'h8c == r_count_17_io_out ? io_r_140_b : _GEN_12979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12981 = 10'h8d == r_count_17_io_out ? io_r_141_b : _GEN_12980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12982 = 10'h8e == r_count_17_io_out ? io_r_142_b : _GEN_12981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12983 = 10'h8f == r_count_17_io_out ? io_r_143_b : _GEN_12982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12984 = 10'h90 == r_count_17_io_out ? io_r_144_b : _GEN_12983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12985 = 10'h91 == r_count_17_io_out ? io_r_145_b : _GEN_12984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12986 = 10'h92 == r_count_17_io_out ? io_r_146_b : _GEN_12985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12987 = 10'h93 == r_count_17_io_out ? io_r_147_b : _GEN_12986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12988 = 10'h94 == r_count_17_io_out ? io_r_148_b : _GEN_12987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12989 = 10'h95 == r_count_17_io_out ? io_r_149_b : _GEN_12988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12990 = 10'h96 == r_count_17_io_out ? io_r_150_b : _GEN_12989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12991 = 10'h97 == r_count_17_io_out ? io_r_151_b : _GEN_12990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12992 = 10'h98 == r_count_17_io_out ? io_r_152_b : _GEN_12991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12993 = 10'h99 == r_count_17_io_out ? io_r_153_b : _GEN_12992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12994 = 10'h9a == r_count_17_io_out ? io_r_154_b : _GEN_12993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12995 = 10'h9b == r_count_17_io_out ? io_r_155_b : _GEN_12994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12996 = 10'h9c == r_count_17_io_out ? io_r_156_b : _GEN_12995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12997 = 10'h9d == r_count_17_io_out ? io_r_157_b : _GEN_12996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12998 = 10'h9e == r_count_17_io_out ? io_r_158_b : _GEN_12997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12999 = 10'h9f == r_count_17_io_out ? io_r_159_b : _GEN_12998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13000 = 10'ha0 == r_count_17_io_out ? io_r_160_b : _GEN_12999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13001 = 10'ha1 == r_count_17_io_out ? io_r_161_b : _GEN_13000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13002 = 10'ha2 == r_count_17_io_out ? io_r_162_b : _GEN_13001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13003 = 10'ha3 == r_count_17_io_out ? io_r_163_b : _GEN_13002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13004 = 10'ha4 == r_count_17_io_out ? io_r_164_b : _GEN_13003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13005 = 10'ha5 == r_count_17_io_out ? io_r_165_b : _GEN_13004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13006 = 10'ha6 == r_count_17_io_out ? io_r_166_b : _GEN_13005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13007 = 10'ha7 == r_count_17_io_out ? io_r_167_b : _GEN_13006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13008 = 10'ha8 == r_count_17_io_out ? io_r_168_b : _GEN_13007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13009 = 10'ha9 == r_count_17_io_out ? io_r_169_b : _GEN_13008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13010 = 10'haa == r_count_17_io_out ? io_r_170_b : _GEN_13009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13011 = 10'hab == r_count_17_io_out ? io_r_171_b : _GEN_13010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13012 = 10'hac == r_count_17_io_out ? io_r_172_b : _GEN_13011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13013 = 10'had == r_count_17_io_out ? io_r_173_b : _GEN_13012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13014 = 10'hae == r_count_17_io_out ? io_r_174_b : _GEN_13013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13015 = 10'haf == r_count_17_io_out ? io_r_175_b : _GEN_13014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13016 = 10'hb0 == r_count_17_io_out ? io_r_176_b : _GEN_13015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13017 = 10'hb1 == r_count_17_io_out ? io_r_177_b : _GEN_13016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13018 = 10'hb2 == r_count_17_io_out ? io_r_178_b : _GEN_13017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13019 = 10'hb3 == r_count_17_io_out ? io_r_179_b : _GEN_13018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13020 = 10'hb4 == r_count_17_io_out ? io_r_180_b : _GEN_13019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13021 = 10'hb5 == r_count_17_io_out ? io_r_181_b : _GEN_13020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13022 = 10'hb6 == r_count_17_io_out ? io_r_182_b : _GEN_13021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13023 = 10'hb7 == r_count_17_io_out ? io_r_183_b : _GEN_13022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13024 = 10'hb8 == r_count_17_io_out ? io_r_184_b : _GEN_13023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13025 = 10'hb9 == r_count_17_io_out ? io_r_185_b : _GEN_13024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13026 = 10'hba == r_count_17_io_out ? io_r_186_b : _GEN_13025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13027 = 10'hbb == r_count_17_io_out ? io_r_187_b : _GEN_13026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13028 = 10'hbc == r_count_17_io_out ? io_r_188_b : _GEN_13027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13029 = 10'hbd == r_count_17_io_out ? io_r_189_b : _GEN_13028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13030 = 10'hbe == r_count_17_io_out ? io_r_190_b : _GEN_13029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13031 = 10'hbf == r_count_17_io_out ? io_r_191_b : _GEN_13030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13032 = 10'hc0 == r_count_17_io_out ? io_r_192_b : _GEN_13031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13033 = 10'hc1 == r_count_17_io_out ? io_r_193_b : _GEN_13032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13034 = 10'hc2 == r_count_17_io_out ? io_r_194_b : _GEN_13033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13035 = 10'hc3 == r_count_17_io_out ? io_r_195_b : _GEN_13034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13036 = 10'hc4 == r_count_17_io_out ? io_r_196_b : _GEN_13035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13037 = 10'hc5 == r_count_17_io_out ? io_r_197_b : _GEN_13036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13038 = 10'hc6 == r_count_17_io_out ? io_r_198_b : _GEN_13037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13039 = 10'hc7 == r_count_17_io_out ? io_r_199_b : _GEN_13038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13040 = 10'hc8 == r_count_17_io_out ? io_r_200_b : _GEN_13039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13041 = 10'hc9 == r_count_17_io_out ? io_r_201_b : _GEN_13040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13042 = 10'hca == r_count_17_io_out ? io_r_202_b : _GEN_13041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13043 = 10'hcb == r_count_17_io_out ? io_r_203_b : _GEN_13042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13044 = 10'hcc == r_count_17_io_out ? io_r_204_b : _GEN_13043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13045 = 10'hcd == r_count_17_io_out ? io_r_205_b : _GEN_13044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13046 = 10'hce == r_count_17_io_out ? io_r_206_b : _GEN_13045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13047 = 10'hcf == r_count_17_io_out ? io_r_207_b : _GEN_13046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13048 = 10'hd0 == r_count_17_io_out ? io_r_208_b : _GEN_13047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13049 = 10'hd1 == r_count_17_io_out ? io_r_209_b : _GEN_13048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13050 = 10'hd2 == r_count_17_io_out ? io_r_210_b : _GEN_13049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13051 = 10'hd3 == r_count_17_io_out ? io_r_211_b : _GEN_13050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13052 = 10'hd4 == r_count_17_io_out ? io_r_212_b : _GEN_13051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13053 = 10'hd5 == r_count_17_io_out ? io_r_213_b : _GEN_13052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13054 = 10'hd6 == r_count_17_io_out ? io_r_214_b : _GEN_13053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13055 = 10'hd7 == r_count_17_io_out ? io_r_215_b : _GEN_13054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13056 = 10'hd8 == r_count_17_io_out ? io_r_216_b : _GEN_13055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13057 = 10'hd9 == r_count_17_io_out ? io_r_217_b : _GEN_13056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13058 = 10'hda == r_count_17_io_out ? io_r_218_b : _GEN_13057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13059 = 10'hdb == r_count_17_io_out ? io_r_219_b : _GEN_13058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13060 = 10'hdc == r_count_17_io_out ? io_r_220_b : _GEN_13059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13061 = 10'hdd == r_count_17_io_out ? io_r_221_b : _GEN_13060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13062 = 10'hde == r_count_17_io_out ? io_r_222_b : _GEN_13061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13063 = 10'hdf == r_count_17_io_out ? io_r_223_b : _GEN_13062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13064 = 10'he0 == r_count_17_io_out ? io_r_224_b : _GEN_13063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13065 = 10'he1 == r_count_17_io_out ? io_r_225_b : _GEN_13064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13066 = 10'he2 == r_count_17_io_out ? io_r_226_b : _GEN_13065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13067 = 10'he3 == r_count_17_io_out ? io_r_227_b : _GEN_13066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13068 = 10'he4 == r_count_17_io_out ? io_r_228_b : _GEN_13067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13069 = 10'he5 == r_count_17_io_out ? io_r_229_b : _GEN_13068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13070 = 10'he6 == r_count_17_io_out ? io_r_230_b : _GEN_13069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13071 = 10'he7 == r_count_17_io_out ? io_r_231_b : _GEN_13070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13072 = 10'he8 == r_count_17_io_out ? io_r_232_b : _GEN_13071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13073 = 10'he9 == r_count_17_io_out ? io_r_233_b : _GEN_13072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13074 = 10'hea == r_count_17_io_out ? io_r_234_b : _GEN_13073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13075 = 10'heb == r_count_17_io_out ? io_r_235_b : _GEN_13074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13076 = 10'hec == r_count_17_io_out ? io_r_236_b : _GEN_13075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13077 = 10'hed == r_count_17_io_out ? io_r_237_b : _GEN_13076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13078 = 10'hee == r_count_17_io_out ? io_r_238_b : _GEN_13077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13079 = 10'hef == r_count_17_io_out ? io_r_239_b : _GEN_13078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13080 = 10'hf0 == r_count_17_io_out ? io_r_240_b : _GEN_13079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13081 = 10'hf1 == r_count_17_io_out ? io_r_241_b : _GEN_13080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13082 = 10'hf2 == r_count_17_io_out ? io_r_242_b : _GEN_13081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13083 = 10'hf3 == r_count_17_io_out ? io_r_243_b : _GEN_13082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13084 = 10'hf4 == r_count_17_io_out ? io_r_244_b : _GEN_13083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13085 = 10'hf5 == r_count_17_io_out ? io_r_245_b : _GEN_13084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13086 = 10'hf6 == r_count_17_io_out ? io_r_246_b : _GEN_13085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13087 = 10'hf7 == r_count_17_io_out ? io_r_247_b : _GEN_13086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13088 = 10'hf8 == r_count_17_io_out ? io_r_248_b : _GEN_13087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13089 = 10'hf9 == r_count_17_io_out ? io_r_249_b : _GEN_13088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13090 = 10'hfa == r_count_17_io_out ? io_r_250_b : _GEN_13089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13091 = 10'hfb == r_count_17_io_out ? io_r_251_b : _GEN_13090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13092 = 10'hfc == r_count_17_io_out ? io_r_252_b : _GEN_13091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13093 = 10'hfd == r_count_17_io_out ? io_r_253_b : _GEN_13092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13094 = 10'hfe == r_count_17_io_out ? io_r_254_b : _GEN_13093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13095 = 10'hff == r_count_17_io_out ? io_r_255_b : _GEN_13094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13096 = 10'h100 == r_count_17_io_out ? io_r_256_b : _GEN_13095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13097 = 10'h101 == r_count_17_io_out ? io_r_257_b : _GEN_13096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13098 = 10'h102 == r_count_17_io_out ? io_r_258_b : _GEN_13097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13099 = 10'h103 == r_count_17_io_out ? io_r_259_b : _GEN_13098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13100 = 10'h104 == r_count_17_io_out ? io_r_260_b : _GEN_13099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13101 = 10'h105 == r_count_17_io_out ? io_r_261_b : _GEN_13100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13102 = 10'h106 == r_count_17_io_out ? io_r_262_b : _GEN_13101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13103 = 10'h107 == r_count_17_io_out ? io_r_263_b : _GEN_13102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13104 = 10'h108 == r_count_17_io_out ? io_r_264_b : _GEN_13103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13105 = 10'h109 == r_count_17_io_out ? io_r_265_b : _GEN_13104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13106 = 10'h10a == r_count_17_io_out ? io_r_266_b : _GEN_13105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13107 = 10'h10b == r_count_17_io_out ? io_r_267_b : _GEN_13106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13108 = 10'h10c == r_count_17_io_out ? io_r_268_b : _GEN_13107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13109 = 10'h10d == r_count_17_io_out ? io_r_269_b : _GEN_13108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13110 = 10'h10e == r_count_17_io_out ? io_r_270_b : _GEN_13109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13111 = 10'h10f == r_count_17_io_out ? io_r_271_b : _GEN_13110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13112 = 10'h110 == r_count_17_io_out ? io_r_272_b : _GEN_13111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13113 = 10'h111 == r_count_17_io_out ? io_r_273_b : _GEN_13112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13114 = 10'h112 == r_count_17_io_out ? io_r_274_b : _GEN_13113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13115 = 10'h113 == r_count_17_io_out ? io_r_275_b : _GEN_13114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13116 = 10'h114 == r_count_17_io_out ? io_r_276_b : _GEN_13115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13117 = 10'h115 == r_count_17_io_out ? io_r_277_b : _GEN_13116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13118 = 10'h116 == r_count_17_io_out ? io_r_278_b : _GEN_13117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13119 = 10'h117 == r_count_17_io_out ? io_r_279_b : _GEN_13118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13120 = 10'h118 == r_count_17_io_out ? io_r_280_b : _GEN_13119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13121 = 10'h119 == r_count_17_io_out ? io_r_281_b : _GEN_13120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13122 = 10'h11a == r_count_17_io_out ? io_r_282_b : _GEN_13121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13123 = 10'h11b == r_count_17_io_out ? io_r_283_b : _GEN_13122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13124 = 10'h11c == r_count_17_io_out ? io_r_284_b : _GEN_13123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13125 = 10'h11d == r_count_17_io_out ? io_r_285_b : _GEN_13124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13126 = 10'h11e == r_count_17_io_out ? io_r_286_b : _GEN_13125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13127 = 10'h11f == r_count_17_io_out ? io_r_287_b : _GEN_13126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13128 = 10'h120 == r_count_17_io_out ? io_r_288_b : _GEN_13127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13129 = 10'h121 == r_count_17_io_out ? io_r_289_b : _GEN_13128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13130 = 10'h122 == r_count_17_io_out ? io_r_290_b : _GEN_13129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13131 = 10'h123 == r_count_17_io_out ? io_r_291_b : _GEN_13130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13132 = 10'h124 == r_count_17_io_out ? io_r_292_b : _GEN_13131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13133 = 10'h125 == r_count_17_io_out ? io_r_293_b : _GEN_13132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13134 = 10'h126 == r_count_17_io_out ? io_r_294_b : _GEN_13133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13135 = 10'h127 == r_count_17_io_out ? io_r_295_b : _GEN_13134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13136 = 10'h128 == r_count_17_io_out ? io_r_296_b : _GEN_13135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13137 = 10'h129 == r_count_17_io_out ? io_r_297_b : _GEN_13136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13138 = 10'h12a == r_count_17_io_out ? io_r_298_b : _GEN_13137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13139 = 10'h12b == r_count_17_io_out ? io_r_299_b : _GEN_13138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13140 = 10'h12c == r_count_17_io_out ? io_r_300_b : _GEN_13139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13141 = 10'h12d == r_count_17_io_out ? io_r_301_b : _GEN_13140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13142 = 10'h12e == r_count_17_io_out ? io_r_302_b : _GEN_13141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13143 = 10'h12f == r_count_17_io_out ? io_r_303_b : _GEN_13142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13144 = 10'h130 == r_count_17_io_out ? io_r_304_b : _GEN_13143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13145 = 10'h131 == r_count_17_io_out ? io_r_305_b : _GEN_13144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13146 = 10'h132 == r_count_17_io_out ? io_r_306_b : _GEN_13145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13147 = 10'h133 == r_count_17_io_out ? io_r_307_b : _GEN_13146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13148 = 10'h134 == r_count_17_io_out ? io_r_308_b : _GEN_13147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13149 = 10'h135 == r_count_17_io_out ? io_r_309_b : _GEN_13148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13150 = 10'h136 == r_count_17_io_out ? io_r_310_b : _GEN_13149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13151 = 10'h137 == r_count_17_io_out ? io_r_311_b : _GEN_13150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13152 = 10'h138 == r_count_17_io_out ? io_r_312_b : _GEN_13151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13153 = 10'h139 == r_count_17_io_out ? io_r_313_b : _GEN_13152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13154 = 10'h13a == r_count_17_io_out ? io_r_314_b : _GEN_13153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13155 = 10'h13b == r_count_17_io_out ? io_r_315_b : _GEN_13154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13156 = 10'h13c == r_count_17_io_out ? io_r_316_b : _GEN_13155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13157 = 10'h13d == r_count_17_io_out ? io_r_317_b : _GEN_13156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13158 = 10'h13e == r_count_17_io_out ? io_r_318_b : _GEN_13157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13159 = 10'h13f == r_count_17_io_out ? io_r_319_b : _GEN_13158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13160 = 10'h140 == r_count_17_io_out ? io_r_320_b : _GEN_13159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13161 = 10'h141 == r_count_17_io_out ? io_r_321_b : _GEN_13160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13162 = 10'h142 == r_count_17_io_out ? io_r_322_b : _GEN_13161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13163 = 10'h143 == r_count_17_io_out ? io_r_323_b : _GEN_13162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13164 = 10'h144 == r_count_17_io_out ? io_r_324_b : _GEN_13163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13165 = 10'h145 == r_count_17_io_out ? io_r_325_b : _GEN_13164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13166 = 10'h146 == r_count_17_io_out ? io_r_326_b : _GEN_13165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13167 = 10'h147 == r_count_17_io_out ? io_r_327_b : _GEN_13166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13168 = 10'h148 == r_count_17_io_out ? io_r_328_b : _GEN_13167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13169 = 10'h149 == r_count_17_io_out ? io_r_329_b : _GEN_13168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13170 = 10'h14a == r_count_17_io_out ? io_r_330_b : _GEN_13169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13171 = 10'h14b == r_count_17_io_out ? io_r_331_b : _GEN_13170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13172 = 10'h14c == r_count_17_io_out ? io_r_332_b : _GEN_13171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13173 = 10'h14d == r_count_17_io_out ? io_r_333_b : _GEN_13172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13174 = 10'h14e == r_count_17_io_out ? io_r_334_b : _GEN_13173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13175 = 10'h14f == r_count_17_io_out ? io_r_335_b : _GEN_13174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13176 = 10'h150 == r_count_17_io_out ? io_r_336_b : _GEN_13175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13177 = 10'h151 == r_count_17_io_out ? io_r_337_b : _GEN_13176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13178 = 10'h152 == r_count_17_io_out ? io_r_338_b : _GEN_13177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13179 = 10'h153 == r_count_17_io_out ? io_r_339_b : _GEN_13178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13180 = 10'h154 == r_count_17_io_out ? io_r_340_b : _GEN_13179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13181 = 10'h155 == r_count_17_io_out ? io_r_341_b : _GEN_13180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13182 = 10'h156 == r_count_17_io_out ? io_r_342_b : _GEN_13181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13183 = 10'h157 == r_count_17_io_out ? io_r_343_b : _GEN_13182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13184 = 10'h158 == r_count_17_io_out ? io_r_344_b : _GEN_13183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13185 = 10'h159 == r_count_17_io_out ? io_r_345_b : _GEN_13184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13186 = 10'h15a == r_count_17_io_out ? io_r_346_b : _GEN_13185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13187 = 10'h15b == r_count_17_io_out ? io_r_347_b : _GEN_13186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13188 = 10'h15c == r_count_17_io_out ? io_r_348_b : _GEN_13187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13189 = 10'h15d == r_count_17_io_out ? io_r_349_b : _GEN_13188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13190 = 10'h15e == r_count_17_io_out ? io_r_350_b : _GEN_13189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13191 = 10'h15f == r_count_17_io_out ? io_r_351_b : _GEN_13190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13192 = 10'h160 == r_count_17_io_out ? io_r_352_b : _GEN_13191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13193 = 10'h161 == r_count_17_io_out ? io_r_353_b : _GEN_13192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13194 = 10'h162 == r_count_17_io_out ? io_r_354_b : _GEN_13193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13195 = 10'h163 == r_count_17_io_out ? io_r_355_b : _GEN_13194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13196 = 10'h164 == r_count_17_io_out ? io_r_356_b : _GEN_13195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13197 = 10'h165 == r_count_17_io_out ? io_r_357_b : _GEN_13196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13198 = 10'h166 == r_count_17_io_out ? io_r_358_b : _GEN_13197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13199 = 10'h167 == r_count_17_io_out ? io_r_359_b : _GEN_13198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13200 = 10'h168 == r_count_17_io_out ? io_r_360_b : _GEN_13199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13201 = 10'h169 == r_count_17_io_out ? io_r_361_b : _GEN_13200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13202 = 10'h16a == r_count_17_io_out ? io_r_362_b : _GEN_13201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13203 = 10'h16b == r_count_17_io_out ? io_r_363_b : _GEN_13202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13204 = 10'h16c == r_count_17_io_out ? io_r_364_b : _GEN_13203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13205 = 10'h16d == r_count_17_io_out ? io_r_365_b : _GEN_13204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13206 = 10'h16e == r_count_17_io_out ? io_r_366_b : _GEN_13205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13207 = 10'h16f == r_count_17_io_out ? io_r_367_b : _GEN_13206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13208 = 10'h170 == r_count_17_io_out ? io_r_368_b : _GEN_13207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13209 = 10'h171 == r_count_17_io_out ? io_r_369_b : _GEN_13208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13210 = 10'h172 == r_count_17_io_out ? io_r_370_b : _GEN_13209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13211 = 10'h173 == r_count_17_io_out ? io_r_371_b : _GEN_13210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13212 = 10'h174 == r_count_17_io_out ? io_r_372_b : _GEN_13211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13213 = 10'h175 == r_count_17_io_out ? io_r_373_b : _GEN_13212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13214 = 10'h176 == r_count_17_io_out ? io_r_374_b : _GEN_13213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13215 = 10'h177 == r_count_17_io_out ? io_r_375_b : _GEN_13214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13216 = 10'h178 == r_count_17_io_out ? io_r_376_b : _GEN_13215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13217 = 10'h179 == r_count_17_io_out ? io_r_377_b : _GEN_13216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13218 = 10'h17a == r_count_17_io_out ? io_r_378_b : _GEN_13217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13219 = 10'h17b == r_count_17_io_out ? io_r_379_b : _GEN_13218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13220 = 10'h17c == r_count_17_io_out ? io_r_380_b : _GEN_13219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13221 = 10'h17d == r_count_17_io_out ? io_r_381_b : _GEN_13220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13222 = 10'h17e == r_count_17_io_out ? io_r_382_b : _GEN_13221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13223 = 10'h17f == r_count_17_io_out ? io_r_383_b : _GEN_13222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13224 = 10'h180 == r_count_17_io_out ? io_r_384_b : _GEN_13223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13225 = 10'h181 == r_count_17_io_out ? io_r_385_b : _GEN_13224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13226 = 10'h182 == r_count_17_io_out ? io_r_386_b : _GEN_13225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13227 = 10'h183 == r_count_17_io_out ? io_r_387_b : _GEN_13226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13228 = 10'h184 == r_count_17_io_out ? io_r_388_b : _GEN_13227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13229 = 10'h185 == r_count_17_io_out ? io_r_389_b : _GEN_13228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13230 = 10'h186 == r_count_17_io_out ? io_r_390_b : _GEN_13229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13231 = 10'h187 == r_count_17_io_out ? io_r_391_b : _GEN_13230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13232 = 10'h188 == r_count_17_io_out ? io_r_392_b : _GEN_13231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13233 = 10'h189 == r_count_17_io_out ? io_r_393_b : _GEN_13232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13234 = 10'h18a == r_count_17_io_out ? io_r_394_b : _GEN_13233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13235 = 10'h18b == r_count_17_io_out ? io_r_395_b : _GEN_13234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13236 = 10'h18c == r_count_17_io_out ? io_r_396_b : _GEN_13235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13237 = 10'h18d == r_count_17_io_out ? io_r_397_b : _GEN_13236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13238 = 10'h18e == r_count_17_io_out ? io_r_398_b : _GEN_13237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13239 = 10'h18f == r_count_17_io_out ? io_r_399_b : _GEN_13238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13240 = 10'h190 == r_count_17_io_out ? io_r_400_b : _GEN_13239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13241 = 10'h191 == r_count_17_io_out ? io_r_401_b : _GEN_13240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13242 = 10'h192 == r_count_17_io_out ? io_r_402_b : _GEN_13241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13243 = 10'h193 == r_count_17_io_out ? io_r_403_b : _GEN_13242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13244 = 10'h194 == r_count_17_io_out ? io_r_404_b : _GEN_13243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13245 = 10'h195 == r_count_17_io_out ? io_r_405_b : _GEN_13244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13246 = 10'h196 == r_count_17_io_out ? io_r_406_b : _GEN_13245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13247 = 10'h197 == r_count_17_io_out ? io_r_407_b : _GEN_13246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13248 = 10'h198 == r_count_17_io_out ? io_r_408_b : _GEN_13247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13249 = 10'h199 == r_count_17_io_out ? io_r_409_b : _GEN_13248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13250 = 10'h19a == r_count_17_io_out ? io_r_410_b : _GEN_13249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13251 = 10'h19b == r_count_17_io_out ? io_r_411_b : _GEN_13250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13252 = 10'h19c == r_count_17_io_out ? io_r_412_b : _GEN_13251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13253 = 10'h19d == r_count_17_io_out ? io_r_413_b : _GEN_13252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13254 = 10'h19e == r_count_17_io_out ? io_r_414_b : _GEN_13253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13255 = 10'h19f == r_count_17_io_out ? io_r_415_b : _GEN_13254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13256 = 10'h1a0 == r_count_17_io_out ? io_r_416_b : _GEN_13255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13257 = 10'h1a1 == r_count_17_io_out ? io_r_417_b : _GEN_13256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13258 = 10'h1a2 == r_count_17_io_out ? io_r_418_b : _GEN_13257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13259 = 10'h1a3 == r_count_17_io_out ? io_r_419_b : _GEN_13258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13260 = 10'h1a4 == r_count_17_io_out ? io_r_420_b : _GEN_13259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13261 = 10'h1a5 == r_count_17_io_out ? io_r_421_b : _GEN_13260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13262 = 10'h1a6 == r_count_17_io_out ? io_r_422_b : _GEN_13261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13263 = 10'h1a7 == r_count_17_io_out ? io_r_423_b : _GEN_13262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13264 = 10'h1a8 == r_count_17_io_out ? io_r_424_b : _GEN_13263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13265 = 10'h1a9 == r_count_17_io_out ? io_r_425_b : _GEN_13264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13266 = 10'h1aa == r_count_17_io_out ? io_r_426_b : _GEN_13265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13267 = 10'h1ab == r_count_17_io_out ? io_r_427_b : _GEN_13266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13268 = 10'h1ac == r_count_17_io_out ? io_r_428_b : _GEN_13267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13269 = 10'h1ad == r_count_17_io_out ? io_r_429_b : _GEN_13268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13270 = 10'h1ae == r_count_17_io_out ? io_r_430_b : _GEN_13269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13271 = 10'h1af == r_count_17_io_out ? io_r_431_b : _GEN_13270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13272 = 10'h1b0 == r_count_17_io_out ? io_r_432_b : _GEN_13271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13273 = 10'h1b1 == r_count_17_io_out ? io_r_433_b : _GEN_13272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13274 = 10'h1b2 == r_count_17_io_out ? io_r_434_b : _GEN_13273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13275 = 10'h1b3 == r_count_17_io_out ? io_r_435_b : _GEN_13274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13276 = 10'h1b4 == r_count_17_io_out ? io_r_436_b : _GEN_13275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13277 = 10'h1b5 == r_count_17_io_out ? io_r_437_b : _GEN_13276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13278 = 10'h1b6 == r_count_17_io_out ? io_r_438_b : _GEN_13277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13279 = 10'h1b7 == r_count_17_io_out ? io_r_439_b : _GEN_13278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13280 = 10'h1b8 == r_count_17_io_out ? io_r_440_b : _GEN_13279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13281 = 10'h1b9 == r_count_17_io_out ? io_r_441_b : _GEN_13280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13282 = 10'h1ba == r_count_17_io_out ? io_r_442_b : _GEN_13281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13283 = 10'h1bb == r_count_17_io_out ? io_r_443_b : _GEN_13282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13284 = 10'h1bc == r_count_17_io_out ? io_r_444_b : _GEN_13283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13285 = 10'h1bd == r_count_17_io_out ? io_r_445_b : _GEN_13284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13286 = 10'h1be == r_count_17_io_out ? io_r_446_b : _GEN_13285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13287 = 10'h1bf == r_count_17_io_out ? io_r_447_b : _GEN_13286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13288 = 10'h1c0 == r_count_17_io_out ? io_r_448_b : _GEN_13287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13289 = 10'h1c1 == r_count_17_io_out ? io_r_449_b : _GEN_13288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13290 = 10'h1c2 == r_count_17_io_out ? io_r_450_b : _GEN_13289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13291 = 10'h1c3 == r_count_17_io_out ? io_r_451_b : _GEN_13290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13292 = 10'h1c4 == r_count_17_io_out ? io_r_452_b : _GEN_13291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13293 = 10'h1c5 == r_count_17_io_out ? io_r_453_b : _GEN_13292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13294 = 10'h1c6 == r_count_17_io_out ? io_r_454_b : _GEN_13293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13295 = 10'h1c7 == r_count_17_io_out ? io_r_455_b : _GEN_13294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13296 = 10'h1c8 == r_count_17_io_out ? io_r_456_b : _GEN_13295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13297 = 10'h1c9 == r_count_17_io_out ? io_r_457_b : _GEN_13296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13298 = 10'h1ca == r_count_17_io_out ? io_r_458_b : _GEN_13297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13299 = 10'h1cb == r_count_17_io_out ? io_r_459_b : _GEN_13298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13300 = 10'h1cc == r_count_17_io_out ? io_r_460_b : _GEN_13299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13301 = 10'h1cd == r_count_17_io_out ? io_r_461_b : _GEN_13300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13302 = 10'h1ce == r_count_17_io_out ? io_r_462_b : _GEN_13301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13303 = 10'h1cf == r_count_17_io_out ? io_r_463_b : _GEN_13302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13304 = 10'h1d0 == r_count_17_io_out ? io_r_464_b : _GEN_13303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13305 = 10'h1d1 == r_count_17_io_out ? io_r_465_b : _GEN_13304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13306 = 10'h1d2 == r_count_17_io_out ? io_r_466_b : _GEN_13305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13307 = 10'h1d3 == r_count_17_io_out ? io_r_467_b : _GEN_13306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13308 = 10'h1d4 == r_count_17_io_out ? io_r_468_b : _GEN_13307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13309 = 10'h1d5 == r_count_17_io_out ? io_r_469_b : _GEN_13308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13310 = 10'h1d6 == r_count_17_io_out ? io_r_470_b : _GEN_13309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13311 = 10'h1d7 == r_count_17_io_out ? io_r_471_b : _GEN_13310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13312 = 10'h1d8 == r_count_17_io_out ? io_r_472_b : _GEN_13311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13313 = 10'h1d9 == r_count_17_io_out ? io_r_473_b : _GEN_13312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13314 = 10'h1da == r_count_17_io_out ? io_r_474_b : _GEN_13313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13315 = 10'h1db == r_count_17_io_out ? io_r_475_b : _GEN_13314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13316 = 10'h1dc == r_count_17_io_out ? io_r_476_b : _GEN_13315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13317 = 10'h1dd == r_count_17_io_out ? io_r_477_b : _GEN_13316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13318 = 10'h1de == r_count_17_io_out ? io_r_478_b : _GEN_13317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13319 = 10'h1df == r_count_17_io_out ? io_r_479_b : _GEN_13318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13320 = 10'h1e0 == r_count_17_io_out ? io_r_480_b : _GEN_13319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13321 = 10'h1e1 == r_count_17_io_out ? io_r_481_b : _GEN_13320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13322 = 10'h1e2 == r_count_17_io_out ? io_r_482_b : _GEN_13321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13323 = 10'h1e3 == r_count_17_io_out ? io_r_483_b : _GEN_13322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13324 = 10'h1e4 == r_count_17_io_out ? io_r_484_b : _GEN_13323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13325 = 10'h1e5 == r_count_17_io_out ? io_r_485_b : _GEN_13324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13326 = 10'h1e6 == r_count_17_io_out ? io_r_486_b : _GEN_13325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13327 = 10'h1e7 == r_count_17_io_out ? io_r_487_b : _GEN_13326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13328 = 10'h1e8 == r_count_17_io_out ? io_r_488_b : _GEN_13327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13329 = 10'h1e9 == r_count_17_io_out ? io_r_489_b : _GEN_13328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13330 = 10'h1ea == r_count_17_io_out ? io_r_490_b : _GEN_13329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13331 = 10'h1eb == r_count_17_io_out ? io_r_491_b : _GEN_13330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13332 = 10'h1ec == r_count_17_io_out ? io_r_492_b : _GEN_13331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13333 = 10'h1ed == r_count_17_io_out ? io_r_493_b : _GEN_13332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13334 = 10'h1ee == r_count_17_io_out ? io_r_494_b : _GEN_13333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13335 = 10'h1ef == r_count_17_io_out ? io_r_495_b : _GEN_13334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13336 = 10'h1f0 == r_count_17_io_out ? io_r_496_b : _GEN_13335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13337 = 10'h1f1 == r_count_17_io_out ? io_r_497_b : _GEN_13336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13338 = 10'h1f2 == r_count_17_io_out ? io_r_498_b : _GEN_13337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13339 = 10'h1f3 == r_count_17_io_out ? io_r_499_b : _GEN_13338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13340 = 10'h1f4 == r_count_17_io_out ? io_r_500_b : _GEN_13339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13341 = 10'h1f5 == r_count_17_io_out ? io_r_501_b : _GEN_13340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13342 = 10'h1f6 == r_count_17_io_out ? io_r_502_b : _GEN_13341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13343 = 10'h1f7 == r_count_17_io_out ? io_r_503_b : _GEN_13342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13344 = 10'h1f8 == r_count_17_io_out ? io_r_504_b : _GEN_13343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13345 = 10'h1f9 == r_count_17_io_out ? io_r_505_b : _GEN_13344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13346 = 10'h1fa == r_count_17_io_out ? io_r_506_b : _GEN_13345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13347 = 10'h1fb == r_count_17_io_out ? io_r_507_b : _GEN_13346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13348 = 10'h1fc == r_count_17_io_out ? io_r_508_b : _GEN_13347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13349 = 10'h1fd == r_count_17_io_out ? io_r_509_b : _GEN_13348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13350 = 10'h1fe == r_count_17_io_out ? io_r_510_b : _GEN_13349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13351 = 10'h1ff == r_count_17_io_out ? io_r_511_b : _GEN_13350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13352 = 10'h200 == r_count_17_io_out ? io_r_512_b : _GEN_13351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13353 = 10'h201 == r_count_17_io_out ? io_r_513_b : _GEN_13352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13354 = 10'h202 == r_count_17_io_out ? io_r_514_b : _GEN_13353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13355 = 10'h203 == r_count_17_io_out ? io_r_515_b : _GEN_13354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13356 = 10'h204 == r_count_17_io_out ? io_r_516_b : _GEN_13355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13357 = 10'h205 == r_count_17_io_out ? io_r_517_b : _GEN_13356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13358 = 10'h206 == r_count_17_io_out ? io_r_518_b : _GEN_13357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13359 = 10'h207 == r_count_17_io_out ? io_r_519_b : _GEN_13358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13360 = 10'h208 == r_count_17_io_out ? io_r_520_b : _GEN_13359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13361 = 10'h209 == r_count_17_io_out ? io_r_521_b : _GEN_13360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13362 = 10'h20a == r_count_17_io_out ? io_r_522_b : _GEN_13361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13363 = 10'h20b == r_count_17_io_out ? io_r_523_b : _GEN_13362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13364 = 10'h20c == r_count_17_io_out ? io_r_524_b : _GEN_13363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13365 = 10'h20d == r_count_17_io_out ? io_r_525_b : _GEN_13364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13366 = 10'h20e == r_count_17_io_out ? io_r_526_b : _GEN_13365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13367 = 10'h20f == r_count_17_io_out ? io_r_527_b : _GEN_13366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13368 = 10'h210 == r_count_17_io_out ? io_r_528_b : _GEN_13367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13369 = 10'h211 == r_count_17_io_out ? io_r_529_b : _GEN_13368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13370 = 10'h212 == r_count_17_io_out ? io_r_530_b : _GEN_13369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13371 = 10'h213 == r_count_17_io_out ? io_r_531_b : _GEN_13370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13372 = 10'h214 == r_count_17_io_out ? io_r_532_b : _GEN_13371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13373 = 10'h215 == r_count_17_io_out ? io_r_533_b : _GEN_13372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13374 = 10'h216 == r_count_17_io_out ? io_r_534_b : _GEN_13373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13375 = 10'h217 == r_count_17_io_out ? io_r_535_b : _GEN_13374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13376 = 10'h218 == r_count_17_io_out ? io_r_536_b : _GEN_13375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13377 = 10'h219 == r_count_17_io_out ? io_r_537_b : _GEN_13376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13378 = 10'h21a == r_count_17_io_out ? io_r_538_b : _GEN_13377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13379 = 10'h21b == r_count_17_io_out ? io_r_539_b : _GEN_13378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13380 = 10'h21c == r_count_17_io_out ? io_r_540_b : _GEN_13379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13381 = 10'h21d == r_count_17_io_out ? io_r_541_b : _GEN_13380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13382 = 10'h21e == r_count_17_io_out ? io_r_542_b : _GEN_13381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13383 = 10'h21f == r_count_17_io_out ? io_r_543_b : _GEN_13382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13384 = 10'h220 == r_count_17_io_out ? io_r_544_b : _GEN_13383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13385 = 10'h221 == r_count_17_io_out ? io_r_545_b : _GEN_13384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13386 = 10'h222 == r_count_17_io_out ? io_r_546_b : _GEN_13385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13387 = 10'h223 == r_count_17_io_out ? io_r_547_b : _GEN_13386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13388 = 10'h224 == r_count_17_io_out ? io_r_548_b : _GEN_13387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13389 = 10'h225 == r_count_17_io_out ? io_r_549_b : _GEN_13388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13390 = 10'h226 == r_count_17_io_out ? io_r_550_b : _GEN_13389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13391 = 10'h227 == r_count_17_io_out ? io_r_551_b : _GEN_13390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13392 = 10'h228 == r_count_17_io_out ? io_r_552_b : _GEN_13391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13393 = 10'h229 == r_count_17_io_out ? io_r_553_b : _GEN_13392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13394 = 10'h22a == r_count_17_io_out ? io_r_554_b : _GEN_13393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13395 = 10'h22b == r_count_17_io_out ? io_r_555_b : _GEN_13394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13396 = 10'h22c == r_count_17_io_out ? io_r_556_b : _GEN_13395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13397 = 10'h22d == r_count_17_io_out ? io_r_557_b : _GEN_13396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13398 = 10'h22e == r_count_17_io_out ? io_r_558_b : _GEN_13397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13399 = 10'h22f == r_count_17_io_out ? io_r_559_b : _GEN_13398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13400 = 10'h230 == r_count_17_io_out ? io_r_560_b : _GEN_13399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13401 = 10'h231 == r_count_17_io_out ? io_r_561_b : _GEN_13400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13402 = 10'h232 == r_count_17_io_out ? io_r_562_b : _GEN_13401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13403 = 10'h233 == r_count_17_io_out ? io_r_563_b : _GEN_13402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13404 = 10'h234 == r_count_17_io_out ? io_r_564_b : _GEN_13403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13405 = 10'h235 == r_count_17_io_out ? io_r_565_b : _GEN_13404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13406 = 10'h236 == r_count_17_io_out ? io_r_566_b : _GEN_13405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13407 = 10'h237 == r_count_17_io_out ? io_r_567_b : _GEN_13406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13408 = 10'h238 == r_count_17_io_out ? io_r_568_b : _GEN_13407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13409 = 10'h239 == r_count_17_io_out ? io_r_569_b : _GEN_13408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13410 = 10'h23a == r_count_17_io_out ? io_r_570_b : _GEN_13409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13411 = 10'h23b == r_count_17_io_out ? io_r_571_b : _GEN_13410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13412 = 10'h23c == r_count_17_io_out ? io_r_572_b : _GEN_13411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13413 = 10'h23d == r_count_17_io_out ? io_r_573_b : _GEN_13412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13414 = 10'h23e == r_count_17_io_out ? io_r_574_b : _GEN_13413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13415 = 10'h23f == r_count_17_io_out ? io_r_575_b : _GEN_13414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13416 = 10'h240 == r_count_17_io_out ? io_r_576_b : _GEN_13415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13417 = 10'h241 == r_count_17_io_out ? io_r_577_b : _GEN_13416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13418 = 10'h242 == r_count_17_io_out ? io_r_578_b : _GEN_13417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13419 = 10'h243 == r_count_17_io_out ? io_r_579_b : _GEN_13418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13420 = 10'h244 == r_count_17_io_out ? io_r_580_b : _GEN_13419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13421 = 10'h245 == r_count_17_io_out ? io_r_581_b : _GEN_13420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13422 = 10'h246 == r_count_17_io_out ? io_r_582_b : _GEN_13421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13423 = 10'h247 == r_count_17_io_out ? io_r_583_b : _GEN_13422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13424 = 10'h248 == r_count_17_io_out ? io_r_584_b : _GEN_13423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13425 = 10'h249 == r_count_17_io_out ? io_r_585_b : _GEN_13424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13426 = 10'h24a == r_count_17_io_out ? io_r_586_b : _GEN_13425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13427 = 10'h24b == r_count_17_io_out ? io_r_587_b : _GEN_13426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13428 = 10'h24c == r_count_17_io_out ? io_r_588_b : _GEN_13427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13429 = 10'h24d == r_count_17_io_out ? io_r_589_b : _GEN_13428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13430 = 10'h24e == r_count_17_io_out ? io_r_590_b : _GEN_13429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13431 = 10'h24f == r_count_17_io_out ? io_r_591_b : _GEN_13430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13432 = 10'h250 == r_count_17_io_out ? io_r_592_b : _GEN_13431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13433 = 10'h251 == r_count_17_io_out ? io_r_593_b : _GEN_13432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13434 = 10'h252 == r_count_17_io_out ? io_r_594_b : _GEN_13433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13435 = 10'h253 == r_count_17_io_out ? io_r_595_b : _GEN_13434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13436 = 10'h254 == r_count_17_io_out ? io_r_596_b : _GEN_13435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13437 = 10'h255 == r_count_17_io_out ? io_r_597_b : _GEN_13436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13438 = 10'h256 == r_count_17_io_out ? io_r_598_b : _GEN_13437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13439 = 10'h257 == r_count_17_io_out ? io_r_599_b : _GEN_13438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13440 = 10'h258 == r_count_17_io_out ? io_r_600_b : _GEN_13439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13441 = 10'h259 == r_count_17_io_out ? io_r_601_b : _GEN_13440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13442 = 10'h25a == r_count_17_io_out ? io_r_602_b : _GEN_13441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13443 = 10'h25b == r_count_17_io_out ? io_r_603_b : _GEN_13442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13444 = 10'h25c == r_count_17_io_out ? io_r_604_b : _GEN_13443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13445 = 10'h25d == r_count_17_io_out ? io_r_605_b : _GEN_13444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13446 = 10'h25e == r_count_17_io_out ? io_r_606_b : _GEN_13445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13447 = 10'h25f == r_count_17_io_out ? io_r_607_b : _GEN_13446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13448 = 10'h260 == r_count_17_io_out ? io_r_608_b : _GEN_13447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13449 = 10'h261 == r_count_17_io_out ? io_r_609_b : _GEN_13448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13450 = 10'h262 == r_count_17_io_out ? io_r_610_b : _GEN_13449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13451 = 10'h263 == r_count_17_io_out ? io_r_611_b : _GEN_13450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13452 = 10'h264 == r_count_17_io_out ? io_r_612_b : _GEN_13451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13453 = 10'h265 == r_count_17_io_out ? io_r_613_b : _GEN_13452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13454 = 10'h266 == r_count_17_io_out ? io_r_614_b : _GEN_13453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13455 = 10'h267 == r_count_17_io_out ? io_r_615_b : _GEN_13454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13456 = 10'h268 == r_count_17_io_out ? io_r_616_b : _GEN_13455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13457 = 10'h269 == r_count_17_io_out ? io_r_617_b : _GEN_13456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13458 = 10'h26a == r_count_17_io_out ? io_r_618_b : _GEN_13457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13459 = 10'h26b == r_count_17_io_out ? io_r_619_b : _GEN_13458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13460 = 10'h26c == r_count_17_io_out ? io_r_620_b : _GEN_13459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13461 = 10'h26d == r_count_17_io_out ? io_r_621_b : _GEN_13460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13462 = 10'h26e == r_count_17_io_out ? io_r_622_b : _GEN_13461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13463 = 10'h26f == r_count_17_io_out ? io_r_623_b : _GEN_13462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13464 = 10'h270 == r_count_17_io_out ? io_r_624_b : _GEN_13463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13465 = 10'h271 == r_count_17_io_out ? io_r_625_b : _GEN_13464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13466 = 10'h272 == r_count_17_io_out ? io_r_626_b : _GEN_13465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13467 = 10'h273 == r_count_17_io_out ? io_r_627_b : _GEN_13466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13468 = 10'h274 == r_count_17_io_out ? io_r_628_b : _GEN_13467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13469 = 10'h275 == r_count_17_io_out ? io_r_629_b : _GEN_13468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13470 = 10'h276 == r_count_17_io_out ? io_r_630_b : _GEN_13469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13471 = 10'h277 == r_count_17_io_out ? io_r_631_b : _GEN_13470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13472 = 10'h278 == r_count_17_io_out ? io_r_632_b : _GEN_13471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13473 = 10'h279 == r_count_17_io_out ? io_r_633_b : _GEN_13472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13474 = 10'h27a == r_count_17_io_out ? io_r_634_b : _GEN_13473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13475 = 10'h27b == r_count_17_io_out ? io_r_635_b : _GEN_13474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13476 = 10'h27c == r_count_17_io_out ? io_r_636_b : _GEN_13475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13477 = 10'h27d == r_count_17_io_out ? io_r_637_b : _GEN_13476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13478 = 10'h27e == r_count_17_io_out ? io_r_638_b : _GEN_13477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13479 = 10'h27f == r_count_17_io_out ? io_r_639_b : _GEN_13478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13480 = 10'h280 == r_count_17_io_out ? io_r_640_b : _GEN_13479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13481 = 10'h281 == r_count_17_io_out ? io_r_641_b : _GEN_13480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13482 = 10'h282 == r_count_17_io_out ? io_r_642_b : _GEN_13481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13483 = 10'h283 == r_count_17_io_out ? io_r_643_b : _GEN_13482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13484 = 10'h284 == r_count_17_io_out ? io_r_644_b : _GEN_13483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13485 = 10'h285 == r_count_17_io_out ? io_r_645_b : _GEN_13484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13486 = 10'h286 == r_count_17_io_out ? io_r_646_b : _GEN_13485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13487 = 10'h287 == r_count_17_io_out ? io_r_647_b : _GEN_13486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13488 = 10'h288 == r_count_17_io_out ? io_r_648_b : _GEN_13487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13489 = 10'h289 == r_count_17_io_out ? io_r_649_b : _GEN_13488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13490 = 10'h28a == r_count_17_io_out ? io_r_650_b : _GEN_13489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13491 = 10'h28b == r_count_17_io_out ? io_r_651_b : _GEN_13490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13492 = 10'h28c == r_count_17_io_out ? io_r_652_b : _GEN_13491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13493 = 10'h28d == r_count_17_io_out ? io_r_653_b : _GEN_13492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13494 = 10'h28e == r_count_17_io_out ? io_r_654_b : _GEN_13493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13495 = 10'h28f == r_count_17_io_out ? io_r_655_b : _GEN_13494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13496 = 10'h290 == r_count_17_io_out ? io_r_656_b : _GEN_13495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13497 = 10'h291 == r_count_17_io_out ? io_r_657_b : _GEN_13496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13498 = 10'h292 == r_count_17_io_out ? io_r_658_b : _GEN_13497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13499 = 10'h293 == r_count_17_io_out ? io_r_659_b : _GEN_13498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13500 = 10'h294 == r_count_17_io_out ? io_r_660_b : _GEN_13499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13501 = 10'h295 == r_count_17_io_out ? io_r_661_b : _GEN_13500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13502 = 10'h296 == r_count_17_io_out ? io_r_662_b : _GEN_13501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13503 = 10'h297 == r_count_17_io_out ? io_r_663_b : _GEN_13502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13504 = 10'h298 == r_count_17_io_out ? io_r_664_b : _GEN_13503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13505 = 10'h299 == r_count_17_io_out ? io_r_665_b : _GEN_13504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13506 = 10'h29a == r_count_17_io_out ? io_r_666_b : _GEN_13505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13507 = 10'h29b == r_count_17_io_out ? io_r_667_b : _GEN_13506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13508 = 10'h29c == r_count_17_io_out ? io_r_668_b : _GEN_13507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13509 = 10'h29d == r_count_17_io_out ? io_r_669_b : _GEN_13508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13510 = 10'h29e == r_count_17_io_out ? io_r_670_b : _GEN_13509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13511 = 10'h29f == r_count_17_io_out ? io_r_671_b : _GEN_13510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13512 = 10'h2a0 == r_count_17_io_out ? io_r_672_b : _GEN_13511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13513 = 10'h2a1 == r_count_17_io_out ? io_r_673_b : _GEN_13512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13514 = 10'h2a2 == r_count_17_io_out ? io_r_674_b : _GEN_13513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13515 = 10'h2a3 == r_count_17_io_out ? io_r_675_b : _GEN_13514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13516 = 10'h2a4 == r_count_17_io_out ? io_r_676_b : _GEN_13515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13517 = 10'h2a5 == r_count_17_io_out ? io_r_677_b : _GEN_13516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13518 = 10'h2a6 == r_count_17_io_out ? io_r_678_b : _GEN_13517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13519 = 10'h2a7 == r_count_17_io_out ? io_r_679_b : _GEN_13518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13520 = 10'h2a8 == r_count_17_io_out ? io_r_680_b : _GEN_13519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13521 = 10'h2a9 == r_count_17_io_out ? io_r_681_b : _GEN_13520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13522 = 10'h2aa == r_count_17_io_out ? io_r_682_b : _GEN_13521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13523 = 10'h2ab == r_count_17_io_out ? io_r_683_b : _GEN_13522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13524 = 10'h2ac == r_count_17_io_out ? io_r_684_b : _GEN_13523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13525 = 10'h2ad == r_count_17_io_out ? io_r_685_b : _GEN_13524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13526 = 10'h2ae == r_count_17_io_out ? io_r_686_b : _GEN_13525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13527 = 10'h2af == r_count_17_io_out ? io_r_687_b : _GEN_13526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13528 = 10'h2b0 == r_count_17_io_out ? io_r_688_b : _GEN_13527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13529 = 10'h2b1 == r_count_17_io_out ? io_r_689_b : _GEN_13528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13530 = 10'h2b2 == r_count_17_io_out ? io_r_690_b : _GEN_13529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13531 = 10'h2b3 == r_count_17_io_out ? io_r_691_b : _GEN_13530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13532 = 10'h2b4 == r_count_17_io_out ? io_r_692_b : _GEN_13531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13533 = 10'h2b5 == r_count_17_io_out ? io_r_693_b : _GEN_13532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13534 = 10'h2b6 == r_count_17_io_out ? io_r_694_b : _GEN_13533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13535 = 10'h2b7 == r_count_17_io_out ? io_r_695_b : _GEN_13534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13536 = 10'h2b8 == r_count_17_io_out ? io_r_696_b : _GEN_13535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13537 = 10'h2b9 == r_count_17_io_out ? io_r_697_b : _GEN_13536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13538 = 10'h2ba == r_count_17_io_out ? io_r_698_b : _GEN_13537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13539 = 10'h2bb == r_count_17_io_out ? io_r_699_b : _GEN_13538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13540 = 10'h2bc == r_count_17_io_out ? io_r_700_b : _GEN_13539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13541 = 10'h2bd == r_count_17_io_out ? io_r_701_b : _GEN_13540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13542 = 10'h2be == r_count_17_io_out ? io_r_702_b : _GEN_13541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13543 = 10'h2bf == r_count_17_io_out ? io_r_703_b : _GEN_13542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13544 = 10'h2c0 == r_count_17_io_out ? io_r_704_b : _GEN_13543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13545 = 10'h2c1 == r_count_17_io_out ? io_r_705_b : _GEN_13544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13546 = 10'h2c2 == r_count_17_io_out ? io_r_706_b : _GEN_13545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13547 = 10'h2c3 == r_count_17_io_out ? io_r_707_b : _GEN_13546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13548 = 10'h2c4 == r_count_17_io_out ? io_r_708_b : _GEN_13547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13549 = 10'h2c5 == r_count_17_io_out ? io_r_709_b : _GEN_13548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13550 = 10'h2c6 == r_count_17_io_out ? io_r_710_b : _GEN_13549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13551 = 10'h2c7 == r_count_17_io_out ? io_r_711_b : _GEN_13550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13552 = 10'h2c8 == r_count_17_io_out ? io_r_712_b : _GEN_13551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13553 = 10'h2c9 == r_count_17_io_out ? io_r_713_b : _GEN_13552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13554 = 10'h2ca == r_count_17_io_out ? io_r_714_b : _GEN_13553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13555 = 10'h2cb == r_count_17_io_out ? io_r_715_b : _GEN_13554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13556 = 10'h2cc == r_count_17_io_out ? io_r_716_b : _GEN_13555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13557 = 10'h2cd == r_count_17_io_out ? io_r_717_b : _GEN_13556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13558 = 10'h2ce == r_count_17_io_out ? io_r_718_b : _GEN_13557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13559 = 10'h2cf == r_count_17_io_out ? io_r_719_b : _GEN_13558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13560 = 10'h2d0 == r_count_17_io_out ? io_r_720_b : _GEN_13559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13561 = 10'h2d1 == r_count_17_io_out ? io_r_721_b : _GEN_13560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13562 = 10'h2d2 == r_count_17_io_out ? io_r_722_b : _GEN_13561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13563 = 10'h2d3 == r_count_17_io_out ? io_r_723_b : _GEN_13562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13564 = 10'h2d4 == r_count_17_io_out ? io_r_724_b : _GEN_13563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13565 = 10'h2d5 == r_count_17_io_out ? io_r_725_b : _GEN_13564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13566 = 10'h2d6 == r_count_17_io_out ? io_r_726_b : _GEN_13565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13567 = 10'h2d7 == r_count_17_io_out ? io_r_727_b : _GEN_13566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13568 = 10'h2d8 == r_count_17_io_out ? io_r_728_b : _GEN_13567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13569 = 10'h2d9 == r_count_17_io_out ? io_r_729_b : _GEN_13568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13570 = 10'h2da == r_count_17_io_out ? io_r_730_b : _GEN_13569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13571 = 10'h2db == r_count_17_io_out ? io_r_731_b : _GEN_13570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13572 = 10'h2dc == r_count_17_io_out ? io_r_732_b : _GEN_13571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13573 = 10'h2dd == r_count_17_io_out ? io_r_733_b : _GEN_13572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13574 = 10'h2de == r_count_17_io_out ? io_r_734_b : _GEN_13573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13575 = 10'h2df == r_count_17_io_out ? io_r_735_b : _GEN_13574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13576 = 10'h2e0 == r_count_17_io_out ? io_r_736_b : _GEN_13575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13577 = 10'h2e1 == r_count_17_io_out ? io_r_737_b : _GEN_13576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13578 = 10'h2e2 == r_count_17_io_out ? io_r_738_b : _GEN_13577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13579 = 10'h2e3 == r_count_17_io_out ? io_r_739_b : _GEN_13578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13580 = 10'h2e4 == r_count_17_io_out ? io_r_740_b : _GEN_13579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13581 = 10'h2e5 == r_count_17_io_out ? io_r_741_b : _GEN_13580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13582 = 10'h2e6 == r_count_17_io_out ? io_r_742_b : _GEN_13581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13583 = 10'h2e7 == r_count_17_io_out ? io_r_743_b : _GEN_13582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13584 = 10'h2e8 == r_count_17_io_out ? io_r_744_b : _GEN_13583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13585 = 10'h2e9 == r_count_17_io_out ? io_r_745_b : _GEN_13584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13586 = 10'h2ea == r_count_17_io_out ? io_r_746_b : _GEN_13585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13587 = 10'h2eb == r_count_17_io_out ? io_r_747_b : _GEN_13586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13588 = 10'h2ec == r_count_17_io_out ? io_r_748_b : _GEN_13587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13591 = 10'h1 == r_count_18_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13592 = 10'h2 == r_count_18_io_out ? io_r_2_b : _GEN_13591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13593 = 10'h3 == r_count_18_io_out ? io_r_3_b : _GEN_13592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13594 = 10'h4 == r_count_18_io_out ? io_r_4_b : _GEN_13593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13595 = 10'h5 == r_count_18_io_out ? io_r_5_b : _GEN_13594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13596 = 10'h6 == r_count_18_io_out ? io_r_6_b : _GEN_13595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13597 = 10'h7 == r_count_18_io_out ? io_r_7_b : _GEN_13596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13598 = 10'h8 == r_count_18_io_out ? io_r_8_b : _GEN_13597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13599 = 10'h9 == r_count_18_io_out ? io_r_9_b : _GEN_13598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13600 = 10'ha == r_count_18_io_out ? io_r_10_b : _GEN_13599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13601 = 10'hb == r_count_18_io_out ? io_r_11_b : _GEN_13600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13602 = 10'hc == r_count_18_io_out ? io_r_12_b : _GEN_13601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13603 = 10'hd == r_count_18_io_out ? io_r_13_b : _GEN_13602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13604 = 10'he == r_count_18_io_out ? io_r_14_b : _GEN_13603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13605 = 10'hf == r_count_18_io_out ? io_r_15_b : _GEN_13604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13606 = 10'h10 == r_count_18_io_out ? io_r_16_b : _GEN_13605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13607 = 10'h11 == r_count_18_io_out ? io_r_17_b : _GEN_13606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13608 = 10'h12 == r_count_18_io_out ? io_r_18_b : _GEN_13607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13609 = 10'h13 == r_count_18_io_out ? io_r_19_b : _GEN_13608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13610 = 10'h14 == r_count_18_io_out ? io_r_20_b : _GEN_13609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13611 = 10'h15 == r_count_18_io_out ? io_r_21_b : _GEN_13610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13612 = 10'h16 == r_count_18_io_out ? io_r_22_b : _GEN_13611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13613 = 10'h17 == r_count_18_io_out ? io_r_23_b : _GEN_13612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13614 = 10'h18 == r_count_18_io_out ? io_r_24_b : _GEN_13613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13615 = 10'h19 == r_count_18_io_out ? io_r_25_b : _GEN_13614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13616 = 10'h1a == r_count_18_io_out ? io_r_26_b : _GEN_13615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13617 = 10'h1b == r_count_18_io_out ? io_r_27_b : _GEN_13616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13618 = 10'h1c == r_count_18_io_out ? io_r_28_b : _GEN_13617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13619 = 10'h1d == r_count_18_io_out ? io_r_29_b : _GEN_13618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13620 = 10'h1e == r_count_18_io_out ? io_r_30_b : _GEN_13619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13621 = 10'h1f == r_count_18_io_out ? io_r_31_b : _GEN_13620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13622 = 10'h20 == r_count_18_io_out ? io_r_32_b : _GEN_13621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13623 = 10'h21 == r_count_18_io_out ? io_r_33_b : _GEN_13622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13624 = 10'h22 == r_count_18_io_out ? io_r_34_b : _GEN_13623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13625 = 10'h23 == r_count_18_io_out ? io_r_35_b : _GEN_13624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13626 = 10'h24 == r_count_18_io_out ? io_r_36_b : _GEN_13625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13627 = 10'h25 == r_count_18_io_out ? io_r_37_b : _GEN_13626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13628 = 10'h26 == r_count_18_io_out ? io_r_38_b : _GEN_13627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13629 = 10'h27 == r_count_18_io_out ? io_r_39_b : _GEN_13628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13630 = 10'h28 == r_count_18_io_out ? io_r_40_b : _GEN_13629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13631 = 10'h29 == r_count_18_io_out ? io_r_41_b : _GEN_13630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13632 = 10'h2a == r_count_18_io_out ? io_r_42_b : _GEN_13631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13633 = 10'h2b == r_count_18_io_out ? io_r_43_b : _GEN_13632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13634 = 10'h2c == r_count_18_io_out ? io_r_44_b : _GEN_13633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13635 = 10'h2d == r_count_18_io_out ? io_r_45_b : _GEN_13634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13636 = 10'h2e == r_count_18_io_out ? io_r_46_b : _GEN_13635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13637 = 10'h2f == r_count_18_io_out ? io_r_47_b : _GEN_13636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13638 = 10'h30 == r_count_18_io_out ? io_r_48_b : _GEN_13637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13639 = 10'h31 == r_count_18_io_out ? io_r_49_b : _GEN_13638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13640 = 10'h32 == r_count_18_io_out ? io_r_50_b : _GEN_13639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13641 = 10'h33 == r_count_18_io_out ? io_r_51_b : _GEN_13640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13642 = 10'h34 == r_count_18_io_out ? io_r_52_b : _GEN_13641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13643 = 10'h35 == r_count_18_io_out ? io_r_53_b : _GEN_13642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13644 = 10'h36 == r_count_18_io_out ? io_r_54_b : _GEN_13643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13645 = 10'h37 == r_count_18_io_out ? io_r_55_b : _GEN_13644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13646 = 10'h38 == r_count_18_io_out ? io_r_56_b : _GEN_13645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13647 = 10'h39 == r_count_18_io_out ? io_r_57_b : _GEN_13646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13648 = 10'h3a == r_count_18_io_out ? io_r_58_b : _GEN_13647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13649 = 10'h3b == r_count_18_io_out ? io_r_59_b : _GEN_13648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13650 = 10'h3c == r_count_18_io_out ? io_r_60_b : _GEN_13649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13651 = 10'h3d == r_count_18_io_out ? io_r_61_b : _GEN_13650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13652 = 10'h3e == r_count_18_io_out ? io_r_62_b : _GEN_13651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13653 = 10'h3f == r_count_18_io_out ? io_r_63_b : _GEN_13652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13654 = 10'h40 == r_count_18_io_out ? io_r_64_b : _GEN_13653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13655 = 10'h41 == r_count_18_io_out ? io_r_65_b : _GEN_13654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13656 = 10'h42 == r_count_18_io_out ? io_r_66_b : _GEN_13655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13657 = 10'h43 == r_count_18_io_out ? io_r_67_b : _GEN_13656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13658 = 10'h44 == r_count_18_io_out ? io_r_68_b : _GEN_13657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13659 = 10'h45 == r_count_18_io_out ? io_r_69_b : _GEN_13658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13660 = 10'h46 == r_count_18_io_out ? io_r_70_b : _GEN_13659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13661 = 10'h47 == r_count_18_io_out ? io_r_71_b : _GEN_13660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13662 = 10'h48 == r_count_18_io_out ? io_r_72_b : _GEN_13661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13663 = 10'h49 == r_count_18_io_out ? io_r_73_b : _GEN_13662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13664 = 10'h4a == r_count_18_io_out ? io_r_74_b : _GEN_13663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13665 = 10'h4b == r_count_18_io_out ? io_r_75_b : _GEN_13664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13666 = 10'h4c == r_count_18_io_out ? io_r_76_b : _GEN_13665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13667 = 10'h4d == r_count_18_io_out ? io_r_77_b : _GEN_13666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13668 = 10'h4e == r_count_18_io_out ? io_r_78_b : _GEN_13667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13669 = 10'h4f == r_count_18_io_out ? io_r_79_b : _GEN_13668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13670 = 10'h50 == r_count_18_io_out ? io_r_80_b : _GEN_13669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13671 = 10'h51 == r_count_18_io_out ? io_r_81_b : _GEN_13670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13672 = 10'h52 == r_count_18_io_out ? io_r_82_b : _GEN_13671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13673 = 10'h53 == r_count_18_io_out ? io_r_83_b : _GEN_13672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13674 = 10'h54 == r_count_18_io_out ? io_r_84_b : _GEN_13673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13675 = 10'h55 == r_count_18_io_out ? io_r_85_b : _GEN_13674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13676 = 10'h56 == r_count_18_io_out ? io_r_86_b : _GEN_13675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13677 = 10'h57 == r_count_18_io_out ? io_r_87_b : _GEN_13676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13678 = 10'h58 == r_count_18_io_out ? io_r_88_b : _GEN_13677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13679 = 10'h59 == r_count_18_io_out ? io_r_89_b : _GEN_13678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13680 = 10'h5a == r_count_18_io_out ? io_r_90_b : _GEN_13679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13681 = 10'h5b == r_count_18_io_out ? io_r_91_b : _GEN_13680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13682 = 10'h5c == r_count_18_io_out ? io_r_92_b : _GEN_13681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13683 = 10'h5d == r_count_18_io_out ? io_r_93_b : _GEN_13682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13684 = 10'h5e == r_count_18_io_out ? io_r_94_b : _GEN_13683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13685 = 10'h5f == r_count_18_io_out ? io_r_95_b : _GEN_13684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13686 = 10'h60 == r_count_18_io_out ? io_r_96_b : _GEN_13685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13687 = 10'h61 == r_count_18_io_out ? io_r_97_b : _GEN_13686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13688 = 10'h62 == r_count_18_io_out ? io_r_98_b : _GEN_13687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13689 = 10'h63 == r_count_18_io_out ? io_r_99_b : _GEN_13688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13690 = 10'h64 == r_count_18_io_out ? io_r_100_b : _GEN_13689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13691 = 10'h65 == r_count_18_io_out ? io_r_101_b : _GEN_13690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13692 = 10'h66 == r_count_18_io_out ? io_r_102_b : _GEN_13691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13693 = 10'h67 == r_count_18_io_out ? io_r_103_b : _GEN_13692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13694 = 10'h68 == r_count_18_io_out ? io_r_104_b : _GEN_13693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13695 = 10'h69 == r_count_18_io_out ? io_r_105_b : _GEN_13694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13696 = 10'h6a == r_count_18_io_out ? io_r_106_b : _GEN_13695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13697 = 10'h6b == r_count_18_io_out ? io_r_107_b : _GEN_13696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13698 = 10'h6c == r_count_18_io_out ? io_r_108_b : _GEN_13697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13699 = 10'h6d == r_count_18_io_out ? io_r_109_b : _GEN_13698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13700 = 10'h6e == r_count_18_io_out ? io_r_110_b : _GEN_13699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13701 = 10'h6f == r_count_18_io_out ? io_r_111_b : _GEN_13700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13702 = 10'h70 == r_count_18_io_out ? io_r_112_b : _GEN_13701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13703 = 10'h71 == r_count_18_io_out ? io_r_113_b : _GEN_13702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13704 = 10'h72 == r_count_18_io_out ? io_r_114_b : _GEN_13703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13705 = 10'h73 == r_count_18_io_out ? io_r_115_b : _GEN_13704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13706 = 10'h74 == r_count_18_io_out ? io_r_116_b : _GEN_13705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13707 = 10'h75 == r_count_18_io_out ? io_r_117_b : _GEN_13706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13708 = 10'h76 == r_count_18_io_out ? io_r_118_b : _GEN_13707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13709 = 10'h77 == r_count_18_io_out ? io_r_119_b : _GEN_13708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13710 = 10'h78 == r_count_18_io_out ? io_r_120_b : _GEN_13709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13711 = 10'h79 == r_count_18_io_out ? io_r_121_b : _GEN_13710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13712 = 10'h7a == r_count_18_io_out ? io_r_122_b : _GEN_13711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13713 = 10'h7b == r_count_18_io_out ? io_r_123_b : _GEN_13712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13714 = 10'h7c == r_count_18_io_out ? io_r_124_b : _GEN_13713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13715 = 10'h7d == r_count_18_io_out ? io_r_125_b : _GEN_13714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13716 = 10'h7e == r_count_18_io_out ? io_r_126_b : _GEN_13715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13717 = 10'h7f == r_count_18_io_out ? io_r_127_b : _GEN_13716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13718 = 10'h80 == r_count_18_io_out ? io_r_128_b : _GEN_13717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13719 = 10'h81 == r_count_18_io_out ? io_r_129_b : _GEN_13718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13720 = 10'h82 == r_count_18_io_out ? io_r_130_b : _GEN_13719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13721 = 10'h83 == r_count_18_io_out ? io_r_131_b : _GEN_13720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13722 = 10'h84 == r_count_18_io_out ? io_r_132_b : _GEN_13721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13723 = 10'h85 == r_count_18_io_out ? io_r_133_b : _GEN_13722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13724 = 10'h86 == r_count_18_io_out ? io_r_134_b : _GEN_13723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13725 = 10'h87 == r_count_18_io_out ? io_r_135_b : _GEN_13724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13726 = 10'h88 == r_count_18_io_out ? io_r_136_b : _GEN_13725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13727 = 10'h89 == r_count_18_io_out ? io_r_137_b : _GEN_13726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13728 = 10'h8a == r_count_18_io_out ? io_r_138_b : _GEN_13727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13729 = 10'h8b == r_count_18_io_out ? io_r_139_b : _GEN_13728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13730 = 10'h8c == r_count_18_io_out ? io_r_140_b : _GEN_13729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13731 = 10'h8d == r_count_18_io_out ? io_r_141_b : _GEN_13730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13732 = 10'h8e == r_count_18_io_out ? io_r_142_b : _GEN_13731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13733 = 10'h8f == r_count_18_io_out ? io_r_143_b : _GEN_13732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13734 = 10'h90 == r_count_18_io_out ? io_r_144_b : _GEN_13733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13735 = 10'h91 == r_count_18_io_out ? io_r_145_b : _GEN_13734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13736 = 10'h92 == r_count_18_io_out ? io_r_146_b : _GEN_13735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13737 = 10'h93 == r_count_18_io_out ? io_r_147_b : _GEN_13736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13738 = 10'h94 == r_count_18_io_out ? io_r_148_b : _GEN_13737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13739 = 10'h95 == r_count_18_io_out ? io_r_149_b : _GEN_13738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13740 = 10'h96 == r_count_18_io_out ? io_r_150_b : _GEN_13739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13741 = 10'h97 == r_count_18_io_out ? io_r_151_b : _GEN_13740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13742 = 10'h98 == r_count_18_io_out ? io_r_152_b : _GEN_13741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13743 = 10'h99 == r_count_18_io_out ? io_r_153_b : _GEN_13742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13744 = 10'h9a == r_count_18_io_out ? io_r_154_b : _GEN_13743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13745 = 10'h9b == r_count_18_io_out ? io_r_155_b : _GEN_13744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13746 = 10'h9c == r_count_18_io_out ? io_r_156_b : _GEN_13745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13747 = 10'h9d == r_count_18_io_out ? io_r_157_b : _GEN_13746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13748 = 10'h9e == r_count_18_io_out ? io_r_158_b : _GEN_13747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13749 = 10'h9f == r_count_18_io_out ? io_r_159_b : _GEN_13748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13750 = 10'ha0 == r_count_18_io_out ? io_r_160_b : _GEN_13749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13751 = 10'ha1 == r_count_18_io_out ? io_r_161_b : _GEN_13750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13752 = 10'ha2 == r_count_18_io_out ? io_r_162_b : _GEN_13751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13753 = 10'ha3 == r_count_18_io_out ? io_r_163_b : _GEN_13752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13754 = 10'ha4 == r_count_18_io_out ? io_r_164_b : _GEN_13753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13755 = 10'ha5 == r_count_18_io_out ? io_r_165_b : _GEN_13754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13756 = 10'ha6 == r_count_18_io_out ? io_r_166_b : _GEN_13755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13757 = 10'ha7 == r_count_18_io_out ? io_r_167_b : _GEN_13756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13758 = 10'ha8 == r_count_18_io_out ? io_r_168_b : _GEN_13757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13759 = 10'ha9 == r_count_18_io_out ? io_r_169_b : _GEN_13758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13760 = 10'haa == r_count_18_io_out ? io_r_170_b : _GEN_13759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13761 = 10'hab == r_count_18_io_out ? io_r_171_b : _GEN_13760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13762 = 10'hac == r_count_18_io_out ? io_r_172_b : _GEN_13761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13763 = 10'had == r_count_18_io_out ? io_r_173_b : _GEN_13762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13764 = 10'hae == r_count_18_io_out ? io_r_174_b : _GEN_13763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13765 = 10'haf == r_count_18_io_out ? io_r_175_b : _GEN_13764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13766 = 10'hb0 == r_count_18_io_out ? io_r_176_b : _GEN_13765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13767 = 10'hb1 == r_count_18_io_out ? io_r_177_b : _GEN_13766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13768 = 10'hb2 == r_count_18_io_out ? io_r_178_b : _GEN_13767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13769 = 10'hb3 == r_count_18_io_out ? io_r_179_b : _GEN_13768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13770 = 10'hb4 == r_count_18_io_out ? io_r_180_b : _GEN_13769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13771 = 10'hb5 == r_count_18_io_out ? io_r_181_b : _GEN_13770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13772 = 10'hb6 == r_count_18_io_out ? io_r_182_b : _GEN_13771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13773 = 10'hb7 == r_count_18_io_out ? io_r_183_b : _GEN_13772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13774 = 10'hb8 == r_count_18_io_out ? io_r_184_b : _GEN_13773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13775 = 10'hb9 == r_count_18_io_out ? io_r_185_b : _GEN_13774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13776 = 10'hba == r_count_18_io_out ? io_r_186_b : _GEN_13775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13777 = 10'hbb == r_count_18_io_out ? io_r_187_b : _GEN_13776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13778 = 10'hbc == r_count_18_io_out ? io_r_188_b : _GEN_13777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13779 = 10'hbd == r_count_18_io_out ? io_r_189_b : _GEN_13778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13780 = 10'hbe == r_count_18_io_out ? io_r_190_b : _GEN_13779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13781 = 10'hbf == r_count_18_io_out ? io_r_191_b : _GEN_13780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13782 = 10'hc0 == r_count_18_io_out ? io_r_192_b : _GEN_13781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13783 = 10'hc1 == r_count_18_io_out ? io_r_193_b : _GEN_13782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13784 = 10'hc2 == r_count_18_io_out ? io_r_194_b : _GEN_13783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13785 = 10'hc3 == r_count_18_io_out ? io_r_195_b : _GEN_13784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13786 = 10'hc4 == r_count_18_io_out ? io_r_196_b : _GEN_13785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13787 = 10'hc5 == r_count_18_io_out ? io_r_197_b : _GEN_13786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13788 = 10'hc6 == r_count_18_io_out ? io_r_198_b : _GEN_13787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13789 = 10'hc7 == r_count_18_io_out ? io_r_199_b : _GEN_13788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13790 = 10'hc8 == r_count_18_io_out ? io_r_200_b : _GEN_13789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13791 = 10'hc9 == r_count_18_io_out ? io_r_201_b : _GEN_13790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13792 = 10'hca == r_count_18_io_out ? io_r_202_b : _GEN_13791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13793 = 10'hcb == r_count_18_io_out ? io_r_203_b : _GEN_13792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13794 = 10'hcc == r_count_18_io_out ? io_r_204_b : _GEN_13793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13795 = 10'hcd == r_count_18_io_out ? io_r_205_b : _GEN_13794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13796 = 10'hce == r_count_18_io_out ? io_r_206_b : _GEN_13795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13797 = 10'hcf == r_count_18_io_out ? io_r_207_b : _GEN_13796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13798 = 10'hd0 == r_count_18_io_out ? io_r_208_b : _GEN_13797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13799 = 10'hd1 == r_count_18_io_out ? io_r_209_b : _GEN_13798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13800 = 10'hd2 == r_count_18_io_out ? io_r_210_b : _GEN_13799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13801 = 10'hd3 == r_count_18_io_out ? io_r_211_b : _GEN_13800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13802 = 10'hd4 == r_count_18_io_out ? io_r_212_b : _GEN_13801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13803 = 10'hd5 == r_count_18_io_out ? io_r_213_b : _GEN_13802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13804 = 10'hd6 == r_count_18_io_out ? io_r_214_b : _GEN_13803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13805 = 10'hd7 == r_count_18_io_out ? io_r_215_b : _GEN_13804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13806 = 10'hd8 == r_count_18_io_out ? io_r_216_b : _GEN_13805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13807 = 10'hd9 == r_count_18_io_out ? io_r_217_b : _GEN_13806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13808 = 10'hda == r_count_18_io_out ? io_r_218_b : _GEN_13807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13809 = 10'hdb == r_count_18_io_out ? io_r_219_b : _GEN_13808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13810 = 10'hdc == r_count_18_io_out ? io_r_220_b : _GEN_13809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13811 = 10'hdd == r_count_18_io_out ? io_r_221_b : _GEN_13810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13812 = 10'hde == r_count_18_io_out ? io_r_222_b : _GEN_13811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13813 = 10'hdf == r_count_18_io_out ? io_r_223_b : _GEN_13812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13814 = 10'he0 == r_count_18_io_out ? io_r_224_b : _GEN_13813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13815 = 10'he1 == r_count_18_io_out ? io_r_225_b : _GEN_13814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13816 = 10'he2 == r_count_18_io_out ? io_r_226_b : _GEN_13815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13817 = 10'he3 == r_count_18_io_out ? io_r_227_b : _GEN_13816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13818 = 10'he4 == r_count_18_io_out ? io_r_228_b : _GEN_13817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13819 = 10'he5 == r_count_18_io_out ? io_r_229_b : _GEN_13818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13820 = 10'he6 == r_count_18_io_out ? io_r_230_b : _GEN_13819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13821 = 10'he7 == r_count_18_io_out ? io_r_231_b : _GEN_13820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13822 = 10'he8 == r_count_18_io_out ? io_r_232_b : _GEN_13821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13823 = 10'he9 == r_count_18_io_out ? io_r_233_b : _GEN_13822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13824 = 10'hea == r_count_18_io_out ? io_r_234_b : _GEN_13823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13825 = 10'heb == r_count_18_io_out ? io_r_235_b : _GEN_13824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13826 = 10'hec == r_count_18_io_out ? io_r_236_b : _GEN_13825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13827 = 10'hed == r_count_18_io_out ? io_r_237_b : _GEN_13826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13828 = 10'hee == r_count_18_io_out ? io_r_238_b : _GEN_13827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13829 = 10'hef == r_count_18_io_out ? io_r_239_b : _GEN_13828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13830 = 10'hf0 == r_count_18_io_out ? io_r_240_b : _GEN_13829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13831 = 10'hf1 == r_count_18_io_out ? io_r_241_b : _GEN_13830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13832 = 10'hf2 == r_count_18_io_out ? io_r_242_b : _GEN_13831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13833 = 10'hf3 == r_count_18_io_out ? io_r_243_b : _GEN_13832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13834 = 10'hf4 == r_count_18_io_out ? io_r_244_b : _GEN_13833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13835 = 10'hf5 == r_count_18_io_out ? io_r_245_b : _GEN_13834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13836 = 10'hf6 == r_count_18_io_out ? io_r_246_b : _GEN_13835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13837 = 10'hf7 == r_count_18_io_out ? io_r_247_b : _GEN_13836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13838 = 10'hf8 == r_count_18_io_out ? io_r_248_b : _GEN_13837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13839 = 10'hf9 == r_count_18_io_out ? io_r_249_b : _GEN_13838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13840 = 10'hfa == r_count_18_io_out ? io_r_250_b : _GEN_13839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13841 = 10'hfb == r_count_18_io_out ? io_r_251_b : _GEN_13840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13842 = 10'hfc == r_count_18_io_out ? io_r_252_b : _GEN_13841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13843 = 10'hfd == r_count_18_io_out ? io_r_253_b : _GEN_13842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13844 = 10'hfe == r_count_18_io_out ? io_r_254_b : _GEN_13843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13845 = 10'hff == r_count_18_io_out ? io_r_255_b : _GEN_13844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13846 = 10'h100 == r_count_18_io_out ? io_r_256_b : _GEN_13845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13847 = 10'h101 == r_count_18_io_out ? io_r_257_b : _GEN_13846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13848 = 10'h102 == r_count_18_io_out ? io_r_258_b : _GEN_13847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13849 = 10'h103 == r_count_18_io_out ? io_r_259_b : _GEN_13848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13850 = 10'h104 == r_count_18_io_out ? io_r_260_b : _GEN_13849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13851 = 10'h105 == r_count_18_io_out ? io_r_261_b : _GEN_13850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13852 = 10'h106 == r_count_18_io_out ? io_r_262_b : _GEN_13851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13853 = 10'h107 == r_count_18_io_out ? io_r_263_b : _GEN_13852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13854 = 10'h108 == r_count_18_io_out ? io_r_264_b : _GEN_13853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13855 = 10'h109 == r_count_18_io_out ? io_r_265_b : _GEN_13854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13856 = 10'h10a == r_count_18_io_out ? io_r_266_b : _GEN_13855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13857 = 10'h10b == r_count_18_io_out ? io_r_267_b : _GEN_13856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13858 = 10'h10c == r_count_18_io_out ? io_r_268_b : _GEN_13857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13859 = 10'h10d == r_count_18_io_out ? io_r_269_b : _GEN_13858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13860 = 10'h10e == r_count_18_io_out ? io_r_270_b : _GEN_13859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13861 = 10'h10f == r_count_18_io_out ? io_r_271_b : _GEN_13860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13862 = 10'h110 == r_count_18_io_out ? io_r_272_b : _GEN_13861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13863 = 10'h111 == r_count_18_io_out ? io_r_273_b : _GEN_13862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13864 = 10'h112 == r_count_18_io_out ? io_r_274_b : _GEN_13863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13865 = 10'h113 == r_count_18_io_out ? io_r_275_b : _GEN_13864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13866 = 10'h114 == r_count_18_io_out ? io_r_276_b : _GEN_13865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13867 = 10'h115 == r_count_18_io_out ? io_r_277_b : _GEN_13866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13868 = 10'h116 == r_count_18_io_out ? io_r_278_b : _GEN_13867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13869 = 10'h117 == r_count_18_io_out ? io_r_279_b : _GEN_13868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13870 = 10'h118 == r_count_18_io_out ? io_r_280_b : _GEN_13869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13871 = 10'h119 == r_count_18_io_out ? io_r_281_b : _GEN_13870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13872 = 10'h11a == r_count_18_io_out ? io_r_282_b : _GEN_13871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13873 = 10'h11b == r_count_18_io_out ? io_r_283_b : _GEN_13872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13874 = 10'h11c == r_count_18_io_out ? io_r_284_b : _GEN_13873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13875 = 10'h11d == r_count_18_io_out ? io_r_285_b : _GEN_13874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13876 = 10'h11e == r_count_18_io_out ? io_r_286_b : _GEN_13875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13877 = 10'h11f == r_count_18_io_out ? io_r_287_b : _GEN_13876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13878 = 10'h120 == r_count_18_io_out ? io_r_288_b : _GEN_13877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13879 = 10'h121 == r_count_18_io_out ? io_r_289_b : _GEN_13878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13880 = 10'h122 == r_count_18_io_out ? io_r_290_b : _GEN_13879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13881 = 10'h123 == r_count_18_io_out ? io_r_291_b : _GEN_13880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13882 = 10'h124 == r_count_18_io_out ? io_r_292_b : _GEN_13881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13883 = 10'h125 == r_count_18_io_out ? io_r_293_b : _GEN_13882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13884 = 10'h126 == r_count_18_io_out ? io_r_294_b : _GEN_13883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13885 = 10'h127 == r_count_18_io_out ? io_r_295_b : _GEN_13884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13886 = 10'h128 == r_count_18_io_out ? io_r_296_b : _GEN_13885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13887 = 10'h129 == r_count_18_io_out ? io_r_297_b : _GEN_13886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13888 = 10'h12a == r_count_18_io_out ? io_r_298_b : _GEN_13887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13889 = 10'h12b == r_count_18_io_out ? io_r_299_b : _GEN_13888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13890 = 10'h12c == r_count_18_io_out ? io_r_300_b : _GEN_13889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13891 = 10'h12d == r_count_18_io_out ? io_r_301_b : _GEN_13890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13892 = 10'h12e == r_count_18_io_out ? io_r_302_b : _GEN_13891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13893 = 10'h12f == r_count_18_io_out ? io_r_303_b : _GEN_13892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13894 = 10'h130 == r_count_18_io_out ? io_r_304_b : _GEN_13893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13895 = 10'h131 == r_count_18_io_out ? io_r_305_b : _GEN_13894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13896 = 10'h132 == r_count_18_io_out ? io_r_306_b : _GEN_13895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13897 = 10'h133 == r_count_18_io_out ? io_r_307_b : _GEN_13896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13898 = 10'h134 == r_count_18_io_out ? io_r_308_b : _GEN_13897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13899 = 10'h135 == r_count_18_io_out ? io_r_309_b : _GEN_13898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13900 = 10'h136 == r_count_18_io_out ? io_r_310_b : _GEN_13899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13901 = 10'h137 == r_count_18_io_out ? io_r_311_b : _GEN_13900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13902 = 10'h138 == r_count_18_io_out ? io_r_312_b : _GEN_13901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13903 = 10'h139 == r_count_18_io_out ? io_r_313_b : _GEN_13902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13904 = 10'h13a == r_count_18_io_out ? io_r_314_b : _GEN_13903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13905 = 10'h13b == r_count_18_io_out ? io_r_315_b : _GEN_13904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13906 = 10'h13c == r_count_18_io_out ? io_r_316_b : _GEN_13905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13907 = 10'h13d == r_count_18_io_out ? io_r_317_b : _GEN_13906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13908 = 10'h13e == r_count_18_io_out ? io_r_318_b : _GEN_13907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13909 = 10'h13f == r_count_18_io_out ? io_r_319_b : _GEN_13908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13910 = 10'h140 == r_count_18_io_out ? io_r_320_b : _GEN_13909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13911 = 10'h141 == r_count_18_io_out ? io_r_321_b : _GEN_13910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13912 = 10'h142 == r_count_18_io_out ? io_r_322_b : _GEN_13911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13913 = 10'h143 == r_count_18_io_out ? io_r_323_b : _GEN_13912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13914 = 10'h144 == r_count_18_io_out ? io_r_324_b : _GEN_13913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13915 = 10'h145 == r_count_18_io_out ? io_r_325_b : _GEN_13914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13916 = 10'h146 == r_count_18_io_out ? io_r_326_b : _GEN_13915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13917 = 10'h147 == r_count_18_io_out ? io_r_327_b : _GEN_13916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13918 = 10'h148 == r_count_18_io_out ? io_r_328_b : _GEN_13917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13919 = 10'h149 == r_count_18_io_out ? io_r_329_b : _GEN_13918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13920 = 10'h14a == r_count_18_io_out ? io_r_330_b : _GEN_13919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13921 = 10'h14b == r_count_18_io_out ? io_r_331_b : _GEN_13920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13922 = 10'h14c == r_count_18_io_out ? io_r_332_b : _GEN_13921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13923 = 10'h14d == r_count_18_io_out ? io_r_333_b : _GEN_13922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13924 = 10'h14e == r_count_18_io_out ? io_r_334_b : _GEN_13923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13925 = 10'h14f == r_count_18_io_out ? io_r_335_b : _GEN_13924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13926 = 10'h150 == r_count_18_io_out ? io_r_336_b : _GEN_13925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13927 = 10'h151 == r_count_18_io_out ? io_r_337_b : _GEN_13926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13928 = 10'h152 == r_count_18_io_out ? io_r_338_b : _GEN_13927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13929 = 10'h153 == r_count_18_io_out ? io_r_339_b : _GEN_13928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13930 = 10'h154 == r_count_18_io_out ? io_r_340_b : _GEN_13929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13931 = 10'h155 == r_count_18_io_out ? io_r_341_b : _GEN_13930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13932 = 10'h156 == r_count_18_io_out ? io_r_342_b : _GEN_13931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13933 = 10'h157 == r_count_18_io_out ? io_r_343_b : _GEN_13932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13934 = 10'h158 == r_count_18_io_out ? io_r_344_b : _GEN_13933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13935 = 10'h159 == r_count_18_io_out ? io_r_345_b : _GEN_13934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13936 = 10'h15a == r_count_18_io_out ? io_r_346_b : _GEN_13935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13937 = 10'h15b == r_count_18_io_out ? io_r_347_b : _GEN_13936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13938 = 10'h15c == r_count_18_io_out ? io_r_348_b : _GEN_13937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13939 = 10'h15d == r_count_18_io_out ? io_r_349_b : _GEN_13938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13940 = 10'h15e == r_count_18_io_out ? io_r_350_b : _GEN_13939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13941 = 10'h15f == r_count_18_io_out ? io_r_351_b : _GEN_13940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13942 = 10'h160 == r_count_18_io_out ? io_r_352_b : _GEN_13941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13943 = 10'h161 == r_count_18_io_out ? io_r_353_b : _GEN_13942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13944 = 10'h162 == r_count_18_io_out ? io_r_354_b : _GEN_13943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13945 = 10'h163 == r_count_18_io_out ? io_r_355_b : _GEN_13944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13946 = 10'h164 == r_count_18_io_out ? io_r_356_b : _GEN_13945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13947 = 10'h165 == r_count_18_io_out ? io_r_357_b : _GEN_13946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13948 = 10'h166 == r_count_18_io_out ? io_r_358_b : _GEN_13947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13949 = 10'h167 == r_count_18_io_out ? io_r_359_b : _GEN_13948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13950 = 10'h168 == r_count_18_io_out ? io_r_360_b : _GEN_13949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13951 = 10'h169 == r_count_18_io_out ? io_r_361_b : _GEN_13950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13952 = 10'h16a == r_count_18_io_out ? io_r_362_b : _GEN_13951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13953 = 10'h16b == r_count_18_io_out ? io_r_363_b : _GEN_13952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13954 = 10'h16c == r_count_18_io_out ? io_r_364_b : _GEN_13953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13955 = 10'h16d == r_count_18_io_out ? io_r_365_b : _GEN_13954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13956 = 10'h16e == r_count_18_io_out ? io_r_366_b : _GEN_13955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13957 = 10'h16f == r_count_18_io_out ? io_r_367_b : _GEN_13956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13958 = 10'h170 == r_count_18_io_out ? io_r_368_b : _GEN_13957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13959 = 10'h171 == r_count_18_io_out ? io_r_369_b : _GEN_13958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13960 = 10'h172 == r_count_18_io_out ? io_r_370_b : _GEN_13959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13961 = 10'h173 == r_count_18_io_out ? io_r_371_b : _GEN_13960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13962 = 10'h174 == r_count_18_io_out ? io_r_372_b : _GEN_13961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13963 = 10'h175 == r_count_18_io_out ? io_r_373_b : _GEN_13962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13964 = 10'h176 == r_count_18_io_out ? io_r_374_b : _GEN_13963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13965 = 10'h177 == r_count_18_io_out ? io_r_375_b : _GEN_13964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13966 = 10'h178 == r_count_18_io_out ? io_r_376_b : _GEN_13965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13967 = 10'h179 == r_count_18_io_out ? io_r_377_b : _GEN_13966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13968 = 10'h17a == r_count_18_io_out ? io_r_378_b : _GEN_13967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13969 = 10'h17b == r_count_18_io_out ? io_r_379_b : _GEN_13968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13970 = 10'h17c == r_count_18_io_out ? io_r_380_b : _GEN_13969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13971 = 10'h17d == r_count_18_io_out ? io_r_381_b : _GEN_13970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13972 = 10'h17e == r_count_18_io_out ? io_r_382_b : _GEN_13971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13973 = 10'h17f == r_count_18_io_out ? io_r_383_b : _GEN_13972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13974 = 10'h180 == r_count_18_io_out ? io_r_384_b : _GEN_13973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13975 = 10'h181 == r_count_18_io_out ? io_r_385_b : _GEN_13974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13976 = 10'h182 == r_count_18_io_out ? io_r_386_b : _GEN_13975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13977 = 10'h183 == r_count_18_io_out ? io_r_387_b : _GEN_13976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13978 = 10'h184 == r_count_18_io_out ? io_r_388_b : _GEN_13977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13979 = 10'h185 == r_count_18_io_out ? io_r_389_b : _GEN_13978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13980 = 10'h186 == r_count_18_io_out ? io_r_390_b : _GEN_13979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13981 = 10'h187 == r_count_18_io_out ? io_r_391_b : _GEN_13980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13982 = 10'h188 == r_count_18_io_out ? io_r_392_b : _GEN_13981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13983 = 10'h189 == r_count_18_io_out ? io_r_393_b : _GEN_13982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13984 = 10'h18a == r_count_18_io_out ? io_r_394_b : _GEN_13983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13985 = 10'h18b == r_count_18_io_out ? io_r_395_b : _GEN_13984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13986 = 10'h18c == r_count_18_io_out ? io_r_396_b : _GEN_13985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13987 = 10'h18d == r_count_18_io_out ? io_r_397_b : _GEN_13986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13988 = 10'h18e == r_count_18_io_out ? io_r_398_b : _GEN_13987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13989 = 10'h18f == r_count_18_io_out ? io_r_399_b : _GEN_13988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13990 = 10'h190 == r_count_18_io_out ? io_r_400_b : _GEN_13989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13991 = 10'h191 == r_count_18_io_out ? io_r_401_b : _GEN_13990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13992 = 10'h192 == r_count_18_io_out ? io_r_402_b : _GEN_13991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13993 = 10'h193 == r_count_18_io_out ? io_r_403_b : _GEN_13992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13994 = 10'h194 == r_count_18_io_out ? io_r_404_b : _GEN_13993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13995 = 10'h195 == r_count_18_io_out ? io_r_405_b : _GEN_13994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13996 = 10'h196 == r_count_18_io_out ? io_r_406_b : _GEN_13995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13997 = 10'h197 == r_count_18_io_out ? io_r_407_b : _GEN_13996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13998 = 10'h198 == r_count_18_io_out ? io_r_408_b : _GEN_13997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13999 = 10'h199 == r_count_18_io_out ? io_r_409_b : _GEN_13998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14000 = 10'h19a == r_count_18_io_out ? io_r_410_b : _GEN_13999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14001 = 10'h19b == r_count_18_io_out ? io_r_411_b : _GEN_14000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14002 = 10'h19c == r_count_18_io_out ? io_r_412_b : _GEN_14001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14003 = 10'h19d == r_count_18_io_out ? io_r_413_b : _GEN_14002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14004 = 10'h19e == r_count_18_io_out ? io_r_414_b : _GEN_14003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14005 = 10'h19f == r_count_18_io_out ? io_r_415_b : _GEN_14004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14006 = 10'h1a0 == r_count_18_io_out ? io_r_416_b : _GEN_14005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14007 = 10'h1a1 == r_count_18_io_out ? io_r_417_b : _GEN_14006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14008 = 10'h1a2 == r_count_18_io_out ? io_r_418_b : _GEN_14007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14009 = 10'h1a3 == r_count_18_io_out ? io_r_419_b : _GEN_14008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14010 = 10'h1a4 == r_count_18_io_out ? io_r_420_b : _GEN_14009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14011 = 10'h1a5 == r_count_18_io_out ? io_r_421_b : _GEN_14010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14012 = 10'h1a6 == r_count_18_io_out ? io_r_422_b : _GEN_14011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14013 = 10'h1a7 == r_count_18_io_out ? io_r_423_b : _GEN_14012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14014 = 10'h1a8 == r_count_18_io_out ? io_r_424_b : _GEN_14013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14015 = 10'h1a9 == r_count_18_io_out ? io_r_425_b : _GEN_14014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14016 = 10'h1aa == r_count_18_io_out ? io_r_426_b : _GEN_14015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14017 = 10'h1ab == r_count_18_io_out ? io_r_427_b : _GEN_14016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14018 = 10'h1ac == r_count_18_io_out ? io_r_428_b : _GEN_14017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14019 = 10'h1ad == r_count_18_io_out ? io_r_429_b : _GEN_14018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14020 = 10'h1ae == r_count_18_io_out ? io_r_430_b : _GEN_14019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14021 = 10'h1af == r_count_18_io_out ? io_r_431_b : _GEN_14020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14022 = 10'h1b0 == r_count_18_io_out ? io_r_432_b : _GEN_14021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14023 = 10'h1b1 == r_count_18_io_out ? io_r_433_b : _GEN_14022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14024 = 10'h1b2 == r_count_18_io_out ? io_r_434_b : _GEN_14023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14025 = 10'h1b3 == r_count_18_io_out ? io_r_435_b : _GEN_14024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14026 = 10'h1b4 == r_count_18_io_out ? io_r_436_b : _GEN_14025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14027 = 10'h1b5 == r_count_18_io_out ? io_r_437_b : _GEN_14026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14028 = 10'h1b6 == r_count_18_io_out ? io_r_438_b : _GEN_14027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14029 = 10'h1b7 == r_count_18_io_out ? io_r_439_b : _GEN_14028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14030 = 10'h1b8 == r_count_18_io_out ? io_r_440_b : _GEN_14029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14031 = 10'h1b9 == r_count_18_io_out ? io_r_441_b : _GEN_14030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14032 = 10'h1ba == r_count_18_io_out ? io_r_442_b : _GEN_14031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14033 = 10'h1bb == r_count_18_io_out ? io_r_443_b : _GEN_14032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14034 = 10'h1bc == r_count_18_io_out ? io_r_444_b : _GEN_14033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14035 = 10'h1bd == r_count_18_io_out ? io_r_445_b : _GEN_14034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14036 = 10'h1be == r_count_18_io_out ? io_r_446_b : _GEN_14035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14037 = 10'h1bf == r_count_18_io_out ? io_r_447_b : _GEN_14036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14038 = 10'h1c0 == r_count_18_io_out ? io_r_448_b : _GEN_14037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14039 = 10'h1c1 == r_count_18_io_out ? io_r_449_b : _GEN_14038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14040 = 10'h1c2 == r_count_18_io_out ? io_r_450_b : _GEN_14039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14041 = 10'h1c3 == r_count_18_io_out ? io_r_451_b : _GEN_14040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14042 = 10'h1c4 == r_count_18_io_out ? io_r_452_b : _GEN_14041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14043 = 10'h1c5 == r_count_18_io_out ? io_r_453_b : _GEN_14042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14044 = 10'h1c6 == r_count_18_io_out ? io_r_454_b : _GEN_14043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14045 = 10'h1c7 == r_count_18_io_out ? io_r_455_b : _GEN_14044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14046 = 10'h1c8 == r_count_18_io_out ? io_r_456_b : _GEN_14045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14047 = 10'h1c9 == r_count_18_io_out ? io_r_457_b : _GEN_14046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14048 = 10'h1ca == r_count_18_io_out ? io_r_458_b : _GEN_14047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14049 = 10'h1cb == r_count_18_io_out ? io_r_459_b : _GEN_14048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14050 = 10'h1cc == r_count_18_io_out ? io_r_460_b : _GEN_14049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14051 = 10'h1cd == r_count_18_io_out ? io_r_461_b : _GEN_14050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14052 = 10'h1ce == r_count_18_io_out ? io_r_462_b : _GEN_14051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14053 = 10'h1cf == r_count_18_io_out ? io_r_463_b : _GEN_14052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14054 = 10'h1d0 == r_count_18_io_out ? io_r_464_b : _GEN_14053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14055 = 10'h1d1 == r_count_18_io_out ? io_r_465_b : _GEN_14054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14056 = 10'h1d2 == r_count_18_io_out ? io_r_466_b : _GEN_14055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14057 = 10'h1d3 == r_count_18_io_out ? io_r_467_b : _GEN_14056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14058 = 10'h1d4 == r_count_18_io_out ? io_r_468_b : _GEN_14057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14059 = 10'h1d5 == r_count_18_io_out ? io_r_469_b : _GEN_14058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14060 = 10'h1d6 == r_count_18_io_out ? io_r_470_b : _GEN_14059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14061 = 10'h1d7 == r_count_18_io_out ? io_r_471_b : _GEN_14060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14062 = 10'h1d8 == r_count_18_io_out ? io_r_472_b : _GEN_14061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14063 = 10'h1d9 == r_count_18_io_out ? io_r_473_b : _GEN_14062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14064 = 10'h1da == r_count_18_io_out ? io_r_474_b : _GEN_14063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14065 = 10'h1db == r_count_18_io_out ? io_r_475_b : _GEN_14064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14066 = 10'h1dc == r_count_18_io_out ? io_r_476_b : _GEN_14065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14067 = 10'h1dd == r_count_18_io_out ? io_r_477_b : _GEN_14066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14068 = 10'h1de == r_count_18_io_out ? io_r_478_b : _GEN_14067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14069 = 10'h1df == r_count_18_io_out ? io_r_479_b : _GEN_14068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14070 = 10'h1e0 == r_count_18_io_out ? io_r_480_b : _GEN_14069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14071 = 10'h1e1 == r_count_18_io_out ? io_r_481_b : _GEN_14070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14072 = 10'h1e2 == r_count_18_io_out ? io_r_482_b : _GEN_14071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14073 = 10'h1e3 == r_count_18_io_out ? io_r_483_b : _GEN_14072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14074 = 10'h1e4 == r_count_18_io_out ? io_r_484_b : _GEN_14073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14075 = 10'h1e5 == r_count_18_io_out ? io_r_485_b : _GEN_14074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14076 = 10'h1e6 == r_count_18_io_out ? io_r_486_b : _GEN_14075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14077 = 10'h1e7 == r_count_18_io_out ? io_r_487_b : _GEN_14076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14078 = 10'h1e8 == r_count_18_io_out ? io_r_488_b : _GEN_14077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14079 = 10'h1e9 == r_count_18_io_out ? io_r_489_b : _GEN_14078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14080 = 10'h1ea == r_count_18_io_out ? io_r_490_b : _GEN_14079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14081 = 10'h1eb == r_count_18_io_out ? io_r_491_b : _GEN_14080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14082 = 10'h1ec == r_count_18_io_out ? io_r_492_b : _GEN_14081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14083 = 10'h1ed == r_count_18_io_out ? io_r_493_b : _GEN_14082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14084 = 10'h1ee == r_count_18_io_out ? io_r_494_b : _GEN_14083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14085 = 10'h1ef == r_count_18_io_out ? io_r_495_b : _GEN_14084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14086 = 10'h1f0 == r_count_18_io_out ? io_r_496_b : _GEN_14085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14087 = 10'h1f1 == r_count_18_io_out ? io_r_497_b : _GEN_14086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14088 = 10'h1f2 == r_count_18_io_out ? io_r_498_b : _GEN_14087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14089 = 10'h1f3 == r_count_18_io_out ? io_r_499_b : _GEN_14088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14090 = 10'h1f4 == r_count_18_io_out ? io_r_500_b : _GEN_14089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14091 = 10'h1f5 == r_count_18_io_out ? io_r_501_b : _GEN_14090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14092 = 10'h1f6 == r_count_18_io_out ? io_r_502_b : _GEN_14091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14093 = 10'h1f7 == r_count_18_io_out ? io_r_503_b : _GEN_14092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14094 = 10'h1f8 == r_count_18_io_out ? io_r_504_b : _GEN_14093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14095 = 10'h1f9 == r_count_18_io_out ? io_r_505_b : _GEN_14094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14096 = 10'h1fa == r_count_18_io_out ? io_r_506_b : _GEN_14095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14097 = 10'h1fb == r_count_18_io_out ? io_r_507_b : _GEN_14096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14098 = 10'h1fc == r_count_18_io_out ? io_r_508_b : _GEN_14097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14099 = 10'h1fd == r_count_18_io_out ? io_r_509_b : _GEN_14098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14100 = 10'h1fe == r_count_18_io_out ? io_r_510_b : _GEN_14099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14101 = 10'h1ff == r_count_18_io_out ? io_r_511_b : _GEN_14100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14102 = 10'h200 == r_count_18_io_out ? io_r_512_b : _GEN_14101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14103 = 10'h201 == r_count_18_io_out ? io_r_513_b : _GEN_14102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14104 = 10'h202 == r_count_18_io_out ? io_r_514_b : _GEN_14103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14105 = 10'h203 == r_count_18_io_out ? io_r_515_b : _GEN_14104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14106 = 10'h204 == r_count_18_io_out ? io_r_516_b : _GEN_14105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14107 = 10'h205 == r_count_18_io_out ? io_r_517_b : _GEN_14106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14108 = 10'h206 == r_count_18_io_out ? io_r_518_b : _GEN_14107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14109 = 10'h207 == r_count_18_io_out ? io_r_519_b : _GEN_14108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14110 = 10'h208 == r_count_18_io_out ? io_r_520_b : _GEN_14109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14111 = 10'h209 == r_count_18_io_out ? io_r_521_b : _GEN_14110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14112 = 10'h20a == r_count_18_io_out ? io_r_522_b : _GEN_14111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14113 = 10'h20b == r_count_18_io_out ? io_r_523_b : _GEN_14112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14114 = 10'h20c == r_count_18_io_out ? io_r_524_b : _GEN_14113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14115 = 10'h20d == r_count_18_io_out ? io_r_525_b : _GEN_14114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14116 = 10'h20e == r_count_18_io_out ? io_r_526_b : _GEN_14115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14117 = 10'h20f == r_count_18_io_out ? io_r_527_b : _GEN_14116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14118 = 10'h210 == r_count_18_io_out ? io_r_528_b : _GEN_14117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14119 = 10'h211 == r_count_18_io_out ? io_r_529_b : _GEN_14118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14120 = 10'h212 == r_count_18_io_out ? io_r_530_b : _GEN_14119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14121 = 10'h213 == r_count_18_io_out ? io_r_531_b : _GEN_14120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14122 = 10'h214 == r_count_18_io_out ? io_r_532_b : _GEN_14121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14123 = 10'h215 == r_count_18_io_out ? io_r_533_b : _GEN_14122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14124 = 10'h216 == r_count_18_io_out ? io_r_534_b : _GEN_14123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14125 = 10'h217 == r_count_18_io_out ? io_r_535_b : _GEN_14124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14126 = 10'h218 == r_count_18_io_out ? io_r_536_b : _GEN_14125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14127 = 10'h219 == r_count_18_io_out ? io_r_537_b : _GEN_14126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14128 = 10'h21a == r_count_18_io_out ? io_r_538_b : _GEN_14127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14129 = 10'h21b == r_count_18_io_out ? io_r_539_b : _GEN_14128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14130 = 10'h21c == r_count_18_io_out ? io_r_540_b : _GEN_14129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14131 = 10'h21d == r_count_18_io_out ? io_r_541_b : _GEN_14130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14132 = 10'h21e == r_count_18_io_out ? io_r_542_b : _GEN_14131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14133 = 10'h21f == r_count_18_io_out ? io_r_543_b : _GEN_14132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14134 = 10'h220 == r_count_18_io_out ? io_r_544_b : _GEN_14133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14135 = 10'h221 == r_count_18_io_out ? io_r_545_b : _GEN_14134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14136 = 10'h222 == r_count_18_io_out ? io_r_546_b : _GEN_14135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14137 = 10'h223 == r_count_18_io_out ? io_r_547_b : _GEN_14136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14138 = 10'h224 == r_count_18_io_out ? io_r_548_b : _GEN_14137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14139 = 10'h225 == r_count_18_io_out ? io_r_549_b : _GEN_14138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14140 = 10'h226 == r_count_18_io_out ? io_r_550_b : _GEN_14139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14141 = 10'h227 == r_count_18_io_out ? io_r_551_b : _GEN_14140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14142 = 10'h228 == r_count_18_io_out ? io_r_552_b : _GEN_14141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14143 = 10'h229 == r_count_18_io_out ? io_r_553_b : _GEN_14142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14144 = 10'h22a == r_count_18_io_out ? io_r_554_b : _GEN_14143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14145 = 10'h22b == r_count_18_io_out ? io_r_555_b : _GEN_14144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14146 = 10'h22c == r_count_18_io_out ? io_r_556_b : _GEN_14145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14147 = 10'h22d == r_count_18_io_out ? io_r_557_b : _GEN_14146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14148 = 10'h22e == r_count_18_io_out ? io_r_558_b : _GEN_14147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14149 = 10'h22f == r_count_18_io_out ? io_r_559_b : _GEN_14148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14150 = 10'h230 == r_count_18_io_out ? io_r_560_b : _GEN_14149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14151 = 10'h231 == r_count_18_io_out ? io_r_561_b : _GEN_14150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14152 = 10'h232 == r_count_18_io_out ? io_r_562_b : _GEN_14151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14153 = 10'h233 == r_count_18_io_out ? io_r_563_b : _GEN_14152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14154 = 10'h234 == r_count_18_io_out ? io_r_564_b : _GEN_14153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14155 = 10'h235 == r_count_18_io_out ? io_r_565_b : _GEN_14154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14156 = 10'h236 == r_count_18_io_out ? io_r_566_b : _GEN_14155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14157 = 10'h237 == r_count_18_io_out ? io_r_567_b : _GEN_14156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14158 = 10'h238 == r_count_18_io_out ? io_r_568_b : _GEN_14157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14159 = 10'h239 == r_count_18_io_out ? io_r_569_b : _GEN_14158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14160 = 10'h23a == r_count_18_io_out ? io_r_570_b : _GEN_14159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14161 = 10'h23b == r_count_18_io_out ? io_r_571_b : _GEN_14160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14162 = 10'h23c == r_count_18_io_out ? io_r_572_b : _GEN_14161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14163 = 10'h23d == r_count_18_io_out ? io_r_573_b : _GEN_14162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14164 = 10'h23e == r_count_18_io_out ? io_r_574_b : _GEN_14163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14165 = 10'h23f == r_count_18_io_out ? io_r_575_b : _GEN_14164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14166 = 10'h240 == r_count_18_io_out ? io_r_576_b : _GEN_14165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14167 = 10'h241 == r_count_18_io_out ? io_r_577_b : _GEN_14166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14168 = 10'h242 == r_count_18_io_out ? io_r_578_b : _GEN_14167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14169 = 10'h243 == r_count_18_io_out ? io_r_579_b : _GEN_14168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14170 = 10'h244 == r_count_18_io_out ? io_r_580_b : _GEN_14169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14171 = 10'h245 == r_count_18_io_out ? io_r_581_b : _GEN_14170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14172 = 10'h246 == r_count_18_io_out ? io_r_582_b : _GEN_14171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14173 = 10'h247 == r_count_18_io_out ? io_r_583_b : _GEN_14172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14174 = 10'h248 == r_count_18_io_out ? io_r_584_b : _GEN_14173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14175 = 10'h249 == r_count_18_io_out ? io_r_585_b : _GEN_14174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14176 = 10'h24a == r_count_18_io_out ? io_r_586_b : _GEN_14175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14177 = 10'h24b == r_count_18_io_out ? io_r_587_b : _GEN_14176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14178 = 10'h24c == r_count_18_io_out ? io_r_588_b : _GEN_14177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14179 = 10'h24d == r_count_18_io_out ? io_r_589_b : _GEN_14178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14180 = 10'h24e == r_count_18_io_out ? io_r_590_b : _GEN_14179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14181 = 10'h24f == r_count_18_io_out ? io_r_591_b : _GEN_14180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14182 = 10'h250 == r_count_18_io_out ? io_r_592_b : _GEN_14181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14183 = 10'h251 == r_count_18_io_out ? io_r_593_b : _GEN_14182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14184 = 10'h252 == r_count_18_io_out ? io_r_594_b : _GEN_14183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14185 = 10'h253 == r_count_18_io_out ? io_r_595_b : _GEN_14184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14186 = 10'h254 == r_count_18_io_out ? io_r_596_b : _GEN_14185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14187 = 10'h255 == r_count_18_io_out ? io_r_597_b : _GEN_14186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14188 = 10'h256 == r_count_18_io_out ? io_r_598_b : _GEN_14187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14189 = 10'h257 == r_count_18_io_out ? io_r_599_b : _GEN_14188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14190 = 10'h258 == r_count_18_io_out ? io_r_600_b : _GEN_14189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14191 = 10'h259 == r_count_18_io_out ? io_r_601_b : _GEN_14190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14192 = 10'h25a == r_count_18_io_out ? io_r_602_b : _GEN_14191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14193 = 10'h25b == r_count_18_io_out ? io_r_603_b : _GEN_14192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14194 = 10'h25c == r_count_18_io_out ? io_r_604_b : _GEN_14193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14195 = 10'h25d == r_count_18_io_out ? io_r_605_b : _GEN_14194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14196 = 10'h25e == r_count_18_io_out ? io_r_606_b : _GEN_14195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14197 = 10'h25f == r_count_18_io_out ? io_r_607_b : _GEN_14196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14198 = 10'h260 == r_count_18_io_out ? io_r_608_b : _GEN_14197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14199 = 10'h261 == r_count_18_io_out ? io_r_609_b : _GEN_14198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14200 = 10'h262 == r_count_18_io_out ? io_r_610_b : _GEN_14199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14201 = 10'h263 == r_count_18_io_out ? io_r_611_b : _GEN_14200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14202 = 10'h264 == r_count_18_io_out ? io_r_612_b : _GEN_14201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14203 = 10'h265 == r_count_18_io_out ? io_r_613_b : _GEN_14202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14204 = 10'h266 == r_count_18_io_out ? io_r_614_b : _GEN_14203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14205 = 10'h267 == r_count_18_io_out ? io_r_615_b : _GEN_14204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14206 = 10'h268 == r_count_18_io_out ? io_r_616_b : _GEN_14205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14207 = 10'h269 == r_count_18_io_out ? io_r_617_b : _GEN_14206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14208 = 10'h26a == r_count_18_io_out ? io_r_618_b : _GEN_14207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14209 = 10'h26b == r_count_18_io_out ? io_r_619_b : _GEN_14208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14210 = 10'h26c == r_count_18_io_out ? io_r_620_b : _GEN_14209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14211 = 10'h26d == r_count_18_io_out ? io_r_621_b : _GEN_14210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14212 = 10'h26e == r_count_18_io_out ? io_r_622_b : _GEN_14211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14213 = 10'h26f == r_count_18_io_out ? io_r_623_b : _GEN_14212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14214 = 10'h270 == r_count_18_io_out ? io_r_624_b : _GEN_14213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14215 = 10'h271 == r_count_18_io_out ? io_r_625_b : _GEN_14214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14216 = 10'h272 == r_count_18_io_out ? io_r_626_b : _GEN_14215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14217 = 10'h273 == r_count_18_io_out ? io_r_627_b : _GEN_14216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14218 = 10'h274 == r_count_18_io_out ? io_r_628_b : _GEN_14217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14219 = 10'h275 == r_count_18_io_out ? io_r_629_b : _GEN_14218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14220 = 10'h276 == r_count_18_io_out ? io_r_630_b : _GEN_14219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14221 = 10'h277 == r_count_18_io_out ? io_r_631_b : _GEN_14220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14222 = 10'h278 == r_count_18_io_out ? io_r_632_b : _GEN_14221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14223 = 10'h279 == r_count_18_io_out ? io_r_633_b : _GEN_14222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14224 = 10'h27a == r_count_18_io_out ? io_r_634_b : _GEN_14223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14225 = 10'h27b == r_count_18_io_out ? io_r_635_b : _GEN_14224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14226 = 10'h27c == r_count_18_io_out ? io_r_636_b : _GEN_14225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14227 = 10'h27d == r_count_18_io_out ? io_r_637_b : _GEN_14226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14228 = 10'h27e == r_count_18_io_out ? io_r_638_b : _GEN_14227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14229 = 10'h27f == r_count_18_io_out ? io_r_639_b : _GEN_14228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14230 = 10'h280 == r_count_18_io_out ? io_r_640_b : _GEN_14229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14231 = 10'h281 == r_count_18_io_out ? io_r_641_b : _GEN_14230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14232 = 10'h282 == r_count_18_io_out ? io_r_642_b : _GEN_14231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14233 = 10'h283 == r_count_18_io_out ? io_r_643_b : _GEN_14232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14234 = 10'h284 == r_count_18_io_out ? io_r_644_b : _GEN_14233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14235 = 10'h285 == r_count_18_io_out ? io_r_645_b : _GEN_14234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14236 = 10'h286 == r_count_18_io_out ? io_r_646_b : _GEN_14235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14237 = 10'h287 == r_count_18_io_out ? io_r_647_b : _GEN_14236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14238 = 10'h288 == r_count_18_io_out ? io_r_648_b : _GEN_14237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14239 = 10'h289 == r_count_18_io_out ? io_r_649_b : _GEN_14238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14240 = 10'h28a == r_count_18_io_out ? io_r_650_b : _GEN_14239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14241 = 10'h28b == r_count_18_io_out ? io_r_651_b : _GEN_14240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14242 = 10'h28c == r_count_18_io_out ? io_r_652_b : _GEN_14241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14243 = 10'h28d == r_count_18_io_out ? io_r_653_b : _GEN_14242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14244 = 10'h28e == r_count_18_io_out ? io_r_654_b : _GEN_14243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14245 = 10'h28f == r_count_18_io_out ? io_r_655_b : _GEN_14244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14246 = 10'h290 == r_count_18_io_out ? io_r_656_b : _GEN_14245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14247 = 10'h291 == r_count_18_io_out ? io_r_657_b : _GEN_14246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14248 = 10'h292 == r_count_18_io_out ? io_r_658_b : _GEN_14247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14249 = 10'h293 == r_count_18_io_out ? io_r_659_b : _GEN_14248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14250 = 10'h294 == r_count_18_io_out ? io_r_660_b : _GEN_14249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14251 = 10'h295 == r_count_18_io_out ? io_r_661_b : _GEN_14250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14252 = 10'h296 == r_count_18_io_out ? io_r_662_b : _GEN_14251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14253 = 10'h297 == r_count_18_io_out ? io_r_663_b : _GEN_14252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14254 = 10'h298 == r_count_18_io_out ? io_r_664_b : _GEN_14253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14255 = 10'h299 == r_count_18_io_out ? io_r_665_b : _GEN_14254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14256 = 10'h29a == r_count_18_io_out ? io_r_666_b : _GEN_14255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14257 = 10'h29b == r_count_18_io_out ? io_r_667_b : _GEN_14256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14258 = 10'h29c == r_count_18_io_out ? io_r_668_b : _GEN_14257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14259 = 10'h29d == r_count_18_io_out ? io_r_669_b : _GEN_14258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14260 = 10'h29e == r_count_18_io_out ? io_r_670_b : _GEN_14259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14261 = 10'h29f == r_count_18_io_out ? io_r_671_b : _GEN_14260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14262 = 10'h2a0 == r_count_18_io_out ? io_r_672_b : _GEN_14261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14263 = 10'h2a1 == r_count_18_io_out ? io_r_673_b : _GEN_14262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14264 = 10'h2a2 == r_count_18_io_out ? io_r_674_b : _GEN_14263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14265 = 10'h2a3 == r_count_18_io_out ? io_r_675_b : _GEN_14264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14266 = 10'h2a4 == r_count_18_io_out ? io_r_676_b : _GEN_14265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14267 = 10'h2a5 == r_count_18_io_out ? io_r_677_b : _GEN_14266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14268 = 10'h2a6 == r_count_18_io_out ? io_r_678_b : _GEN_14267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14269 = 10'h2a7 == r_count_18_io_out ? io_r_679_b : _GEN_14268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14270 = 10'h2a8 == r_count_18_io_out ? io_r_680_b : _GEN_14269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14271 = 10'h2a9 == r_count_18_io_out ? io_r_681_b : _GEN_14270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14272 = 10'h2aa == r_count_18_io_out ? io_r_682_b : _GEN_14271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14273 = 10'h2ab == r_count_18_io_out ? io_r_683_b : _GEN_14272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14274 = 10'h2ac == r_count_18_io_out ? io_r_684_b : _GEN_14273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14275 = 10'h2ad == r_count_18_io_out ? io_r_685_b : _GEN_14274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14276 = 10'h2ae == r_count_18_io_out ? io_r_686_b : _GEN_14275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14277 = 10'h2af == r_count_18_io_out ? io_r_687_b : _GEN_14276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14278 = 10'h2b0 == r_count_18_io_out ? io_r_688_b : _GEN_14277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14279 = 10'h2b1 == r_count_18_io_out ? io_r_689_b : _GEN_14278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14280 = 10'h2b2 == r_count_18_io_out ? io_r_690_b : _GEN_14279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14281 = 10'h2b3 == r_count_18_io_out ? io_r_691_b : _GEN_14280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14282 = 10'h2b4 == r_count_18_io_out ? io_r_692_b : _GEN_14281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14283 = 10'h2b5 == r_count_18_io_out ? io_r_693_b : _GEN_14282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14284 = 10'h2b6 == r_count_18_io_out ? io_r_694_b : _GEN_14283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14285 = 10'h2b7 == r_count_18_io_out ? io_r_695_b : _GEN_14284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14286 = 10'h2b8 == r_count_18_io_out ? io_r_696_b : _GEN_14285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14287 = 10'h2b9 == r_count_18_io_out ? io_r_697_b : _GEN_14286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14288 = 10'h2ba == r_count_18_io_out ? io_r_698_b : _GEN_14287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14289 = 10'h2bb == r_count_18_io_out ? io_r_699_b : _GEN_14288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14290 = 10'h2bc == r_count_18_io_out ? io_r_700_b : _GEN_14289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14291 = 10'h2bd == r_count_18_io_out ? io_r_701_b : _GEN_14290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14292 = 10'h2be == r_count_18_io_out ? io_r_702_b : _GEN_14291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14293 = 10'h2bf == r_count_18_io_out ? io_r_703_b : _GEN_14292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14294 = 10'h2c0 == r_count_18_io_out ? io_r_704_b : _GEN_14293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14295 = 10'h2c1 == r_count_18_io_out ? io_r_705_b : _GEN_14294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14296 = 10'h2c2 == r_count_18_io_out ? io_r_706_b : _GEN_14295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14297 = 10'h2c3 == r_count_18_io_out ? io_r_707_b : _GEN_14296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14298 = 10'h2c4 == r_count_18_io_out ? io_r_708_b : _GEN_14297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14299 = 10'h2c5 == r_count_18_io_out ? io_r_709_b : _GEN_14298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14300 = 10'h2c6 == r_count_18_io_out ? io_r_710_b : _GEN_14299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14301 = 10'h2c7 == r_count_18_io_out ? io_r_711_b : _GEN_14300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14302 = 10'h2c8 == r_count_18_io_out ? io_r_712_b : _GEN_14301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14303 = 10'h2c9 == r_count_18_io_out ? io_r_713_b : _GEN_14302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14304 = 10'h2ca == r_count_18_io_out ? io_r_714_b : _GEN_14303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14305 = 10'h2cb == r_count_18_io_out ? io_r_715_b : _GEN_14304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14306 = 10'h2cc == r_count_18_io_out ? io_r_716_b : _GEN_14305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14307 = 10'h2cd == r_count_18_io_out ? io_r_717_b : _GEN_14306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14308 = 10'h2ce == r_count_18_io_out ? io_r_718_b : _GEN_14307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14309 = 10'h2cf == r_count_18_io_out ? io_r_719_b : _GEN_14308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14310 = 10'h2d0 == r_count_18_io_out ? io_r_720_b : _GEN_14309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14311 = 10'h2d1 == r_count_18_io_out ? io_r_721_b : _GEN_14310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14312 = 10'h2d2 == r_count_18_io_out ? io_r_722_b : _GEN_14311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14313 = 10'h2d3 == r_count_18_io_out ? io_r_723_b : _GEN_14312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14314 = 10'h2d4 == r_count_18_io_out ? io_r_724_b : _GEN_14313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14315 = 10'h2d5 == r_count_18_io_out ? io_r_725_b : _GEN_14314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14316 = 10'h2d6 == r_count_18_io_out ? io_r_726_b : _GEN_14315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14317 = 10'h2d7 == r_count_18_io_out ? io_r_727_b : _GEN_14316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14318 = 10'h2d8 == r_count_18_io_out ? io_r_728_b : _GEN_14317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14319 = 10'h2d9 == r_count_18_io_out ? io_r_729_b : _GEN_14318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14320 = 10'h2da == r_count_18_io_out ? io_r_730_b : _GEN_14319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14321 = 10'h2db == r_count_18_io_out ? io_r_731_b : _GEN_14320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14322 = 10'h2dc == r_count_18_io_out ? io_r_732_b : _GEN_14321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14323 = 10'h2dd == r_count_18_io_out ? io_r_733_b : _GEN_14322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14324 = 10'h2de == r_count_18_io_out ? io_r_734_b : _GEN_14323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14325 = 10'h2df == r_count_18_io_out ? io_r_735_b : _GEN_14324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14326 = 10'h2e0 == r_count_18_io_out ? io_r_736_b : _GEN_14325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14327 = 10'h2e1 == r_count_18_io_out ? io_r_737_b : _GEN_14326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14328 = 10'h2e2 == r_count_18_io_out ? io_r_738_b : _GEN_14327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14329 = 10'h2e3 == r_count_18_io_out ? io_r_739_b : _GEN_14328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14330 = 10'h2e4 == r_count_18_io_out ? io_r_740_b : _GEN_14329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14331 = 10'h2e5 == r_count_18_io_out ? io_r_741_b : _GEN_14330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14332 = 10'h2e6 == r_count_18_io_out ? io_r_742_b : _GEN_14331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14333 = 10'h2e7 == r_count_18_io_out ? io_r_743_b : _GEN_14332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14334 = 10'h2e8 == r_count_18_io_out ? io_r_744_b : _GEN_14333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14335 = 10'h2e9 == r_count_18_io_out ? io_r_745_b : _GEN_14334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14336 = 10'h2ea == r_count_18_io_out ? io_r_746_b : _GEN_14335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14337 = 10'h2eb == r_count_18_io_out ? io_r_747_b : _GEN_14336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14338 = 10'h2ec == r_count_18_io_out ? io_r_748_b : _GEN_14337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14341 = 10'h1 == r_count_19_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14342 = 10'h2 == r_count_19_io_out ? io_r_2_b : _GEN_14341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14343 = 10'h3 == r_count_19_io_out ? io_r_3_b : _GEN_14342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14344 = 10'h4 == r_count_19_io_out ? io_r_4_b : _GEN_14343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14345 = 10'h5 == r_count_19_io_out ? io_r_5_b : _GEN_14344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14346 = 10'h6 == r_count_19_io_out ? io_r_6_b : _GEN_14345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14347 = 10'h7 == r_count_19_io_out ? io_r_7_b : _GEN_14346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14348 = 10'h8 == r_count_19_io_out ? io_r_8_b : _GEN_14347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14349 = 10'h9 == r_count_19_io_out ? io_r_9_b : _GEN_14348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14350 = 10'ha == r_count_19_io_out ? io_r_10_b : _GEN_14349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14351 = 10'hb == r_count_19_io_out ? io_r_11_b : _GEN_14350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14352 = 10'hc == r_count_19_io_out ? io_r_12_b : _GEN_14351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14353 = 10'hd == r_count_19_io_out ? io_r_13_b : _GEN_14352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14354 = 10'he == r_count_19_io_out ? io_r_14_b : _GEN_14353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14355 = 10'hf == r_count_19_io_out ? io_r_15_b : _GEN_14354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14356 = 10'h10 == r_count_19_io_out ? io_r_16_b : _GEN_14355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14357 = 10'h11 == r_count_19_io_out ? io_r_17_b : _GEN_14356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14358 = 10'h12 == r_count_19_io_out ? io_r_18_b : _GEN_14357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14359 = 10'h13 == r_count_19_io_out ? io_r_19_b : _GEN_14358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14360 = 10'h14 == r_count_19_io_out ? io_r_20_b : _GEN_14359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14361 = 10'h15 == r_count_19_io_out ? io_r_21_b : _GEN_14360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14362 = 10'h16 == r_count_19_io_out ? io_r_22_b : _GEN_14361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14363 = 10'h17 == r_count_19_io_out ? io_r_23_b : _GEN_14362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14364 = 10'h18 == r_count_19_io_out ? io_r_24_b : _GEN_14363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14365 = 10'h19 == r_count_19_io_out ? io_r_25_b : _GEN_14364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14366 = 10'h1a == r_count_19_io_out ? io_r_26_b : _GEN_14365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14367 = 10'h1b == r_count_19_io_out ? io_r_27_b : _GEN_14366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14368 = 10'h1c == r_count_19_io_out ? io_r_28_b : _GEN_14367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14369 = 10'h1d == r_count_19_io_out ? io_r_29_b : _GEN_14368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14370 = 10'h1e == r_count_19_io_out ? io_r_30_b : _GEN_14369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14371 = 10'h1f == r_count_19_io_out ? io_r_31_b : _GEN_14370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14372 = 10'h20 == r_count_19_io_out ? io_r_32_b : _GEN_14371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14373 = 10'h21 == r_count_19_io_out ? io_r_33_b : _GEN_14372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14374 = 10'h22 == r_count_19_io_out ? io_r_34_b : _GEN_14373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14375 = 10'h23 == r_count_19_io_out ? io_r_35_b : _GEN_14374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14376 = 10'h24 == r_count_19_io_out ? io_r_36_b : _GEN_14375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14377 = 10'h25 == r_count_19_io_out ? io_r_37_b : _GEN_14376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14378 = 10'h26 == r_count_19_io_out ? io_r_38_b : _GEN_14377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14379 = 10'h27 == r_count_19_io_out ? io_r_39_b : _GEN_14378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14380 = 10'h28 == r_count_19_io_out ? io_r_40_b : _GEN_14379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14381 = 10'h29 == r_count_19_io_out ? io_r_41_b : _GEN_14380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14382 = 10'h2a == r_count_19_io_out ? io_r_42_b : _GEN_14381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14383 = 10'h2b == r_count_19_io_out ? io_r_43_b : _GEN_14382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14384 = 10'h2c == r_count_19_io_out ? io_r_44_b : _GEN_14383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14385 = 10'h2d == r_count_19_io_out ? io_r_45_b : _GEN_14384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14386 = 10'h2e == r_count_19_io_out ? io_r_46_b : _GEN_14385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14387 = 10'h2f == r_count_19_io_out ? io_r_47_b : _GEN_14386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14388 = 10'h30 == r_count_19_io_out ? io_r_48_b : _GEN_14387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14389 = 10'h31 == r_count_19_io_out ? io_r_49_b : _GEN_14388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14390 = 10'h32 == r_count_19_io_out ? io_r_50_b : _GEN_14389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14391 = 10'h33 == r_count_19_io_out ? io_r_51_b : _GEN_14390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14392 = 10'h34 == r_count_19_io_out ? io_r_52_b : _GEN_14391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14393 = 10'h35 == r_count_19_io_out ? io_r_53_b : _GEN_14392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14394 = 10'h36 == r_count_19_io_out ? io_r_54_b : _GEN_14393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14395 = 10'h37 == r_count_19_io_out ? io_r_55_b : _GEN_14394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14396 = 10'h38 == r_count_19_io_out ? io_r_56_b : _GEN_14395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14397 = 10'h39 == r_count_19_io_out ? io_r_57_b : _GEN_14396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14398 = 10'h3a == r_count_19_io_out ? io_r_58_b : _GEN_14397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14399 = 10'h3b == r_count_19_io_out ? io_r_59_b : _GEN_14398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14400 = 10'h3c == r_count_19_io_out ? io_r_60_b : _GEN_14399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14401 = 10'h3d == r_count_19_io_out ? io_r_61_b : _GEN_14400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14402 = 10'h3e == r_count_19_io_out ? io_r_62_b : _GEN_14401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14403 = 10'h3f == r_count_19_io_out ? io_r_63_b : _GEN_14402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14404 = 10'h40 == r_count_19_io_out ? io_r_64_b : _GEN_14403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14405 = 10'h41 == r_count_19_io_out ? io_r_65_b : _GEN_14404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14406 = 10'h42 == r_count_19_io_out ? io_r_66_b : _GEN_14405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14407 = 10'h43 == r_count_19_io_out ? io_r_67_b : _GEN_14406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14408 = 10'h44 == r_count_19_io_out ? io_r_68_b : _GEN_14407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14409 = 10'h45 == r_count_19_io_out ? io_r_69_b : _GEN_14408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14410 = 10'h46 == r_count_19_io_out ? io_r_70_b : _GEN_14409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14411 = 10'h47 == r_count_19_io_out ? io_r_71_b : _GEN_14410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14412 = 10'h48 == r_count_19_io_out ? io_r_72_b : _GEN_14411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14413 = 10'h49 == r_count_19_io_out ? io_r_73_b : _GEN_14412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14414 = 10'h4a == r_count_19_io_out ? io_r_74_b : _GEN_14413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14415 = 10'h4b == r_count_19_io_out ? io_r_75_b : _GEN_14414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14416 = 10'h4c == r_count_19_io_out ? io_r_76_b : _GEN_14415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14417 = 10'h4d == r_count_19_io_out ? io_r_77_b : _GEN_14416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14418 = 10'h4e == r_count_19_io_out ? io_r_78_b : _GEN_14417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14419 = 10'h4f == r_count_19_io_out ? io_r_79_b : _GEN_14418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14420 = 10'h50 == r_count_19_io_out ? io_r_80_b : _GEN_14419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14421 = 10'h51 == r_count_19_io_out ? io_r_81_b : _GEN_14420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14422 = 10'h52 == r_count_19_io_out ? io_r_82_b : _GEN_14421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14423 = 10'h53 == r_count_19_io_out ? io_r_83_b : _GEN_14422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14424 = 10'h54 == r_count_19_io_out ? io_r_84_b : _GEN_14423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14425 = 10'h55 == r_count_19_io_out ? io_r_85_b : _GEN_14424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14426 = 10'h56 == r_count_19_io_out ? io_r_86_b : _GEN_14425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14427 = 10'h57 == r_count_19_io_out ? io_r_87_b : _GEN_14426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14428 = 10'h58 == r_count_19_io_out ? io_r_88_b : _GEN_14427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14429 = 10'h59 == r_count_19_io_out ? io_r_89_b : _GEN_14428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14430 = 10'h5a == r_count_19_io_out ? io_r_90_b : _GEN_14429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14431 = 10'h5b == r_count_19_io_out ? io_r_91_b : _GEN_14430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14432 = 10'h5c == r_count_19_io_out ? io_r_92_b : _GEN_14431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14433 = 10'h5d == r_count_19_io_out ? io_r_93_b : _GEN_14432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14434 = 10'h5e == r_count_19_io_out ? io_r_94_b : _GEN_14433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14435 = 10'h5f == r_count_19_io_out ? io_r_95_b : _GEN_14434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14436 = 10'h60 == r_count_19_io_out ? io_r_96_b : _GEN_14435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14437 = 10'h61 == r_count_19_io_out ? io_r_97_b : _GEN_14436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14438 = 10'h62 == r_count_19_io_out ? io_r_98_b : _GEN_14437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14439 = 10'h63 == r_count_19_io_out ? io_r_99_b : _GEN_14438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14440 = 10'h64 == r_count_19_io_out ? io_r_100_b : _GEN_14439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14441 = 10'h65 == r_count_19_io_out ? io_r_101_b : _GEN_14440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14442 = 10'h66 == r_count_19_io_out ? io_r_102_b : _GEN_14441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14443 = 10'h67 == r_count_19_io_out ? io_r_103_b : _GEN_14442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14444 = 10'h68 == r_count_19_io_out ? io_r_104_b : _GEN_14443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14445 = 10'h69 == r_count_19_io_out ? io_r_105_b : _GEN_14444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14446 = 10'h6a == r_count_19_io_out ? io_r_106_b : _GEN_14445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14447 = 10'h6b == r_count_19_io_out ? io_r_107_b : _GEN_14446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14448 = 10'h6c == r_count_19_io_out ? io_r_108_b : _GEN_14447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14449 = 10'h6d == r_count_19_io_out ? io_r_109_b : _GEN_14448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14450 = 10'h6e == r_count_19_io_out ? io_r_110_b : _GEN_14449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14451 = 10'h6f == r_count_19_io_out ? io_r_111_b : _GEN_14450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14452 = 10'h70 == r_count_19_io_out ? io_r_112_b : _GEN_14451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14453 = 10'h71 == r_count_19_io_out ? io_r_113_b : _GEN_14452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14454 = 10'h72 == r_count_19_io_out ? io_r_114_b : _GEN_14453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14455 = 10'h73 == r_count_19_io_out ? io_r_115_b : _GEN_14454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14456 = 10'h74 == r_count_19_io_out ? io_r_116_b : _GEN_14455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14457 = 10'h75 == r_count_19_io_out ? io_r_117_b : _GEN_14456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14458 = 10'h76 == r_count_19_io_out ? io_r_118_b : _GEN_14457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14459 = 10'h77 == r_count_19_io_out ? io_r_119_b : _GEN_14458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14460 = 10'h78 == r_count_19_io_out ? io_r_120_b : _GEN_14459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14461 = 10'h79 == r_count_19_io_out ? io_r_121_b : _GEN_14460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14462 = 10'h7a == r_count_19_io_out ? io_r_122_b : _GEN_14461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14463 = 10'h7b == r_count_19_io_out ? io_r_123_b : _GEN_14462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14464 = 10'h7c == r_count_19_io_out ? io_r_124_b : _GEN_14463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14465 = 10'h7d == r_count_19_io_out ? io_r_125_b : _GEN_14464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14466 = 10'h7e == r_count_19_io_out ? io_r_126_b : _GEN_14465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14467 = 10'h7f == r_count_19_io_out ? io_r_127_b : _GEN_14466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14468 = 10'h80 == r_count_19_io_out ? io_r_128_b : _GEN_14467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14469 = 10'h81 == r_count_19_io_out ? io_r_129_b : _GEN_14468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14470 = 10'h82 == r_count_19_io_out ? io_r_130_b : _GEN_14469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14471 = 10'h83 == r_count_19_io_out ? io_r_131_b : _GEN_14470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14472 = 10'h84 == r_count_19_io_out ? io_r_132_b : _GEN_14471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14473 = 10'h85 == r_count_19_io_out ? io_r_133_b : _GEN_14472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14474 = 10'h86 == r_count_19_io_out ? io_r_134_b : _GEN_14473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14475 = 10'h87 == r_count_19_io_out ? io_r_135_b : _GEN_14474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14476 = 10'h88 == r_count_19_io_out ? io_r_136_b : _GEN_14475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14477 = 10'h89 == r_count_19_io_out ? io_r_137_b : _GEN_14476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14478 = 10'h8a == r_count_19_io_out ? io_r_138_b : _GEN_14477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14479 = 10'h8b == r_count_19_io_out ? io_r_139_b : _GEN_14478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14480 = 10'h8c == r_count_19_io_out ? io_r_140_b : _GEN_14479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14481 = 10'h8d == r_count_19_io_out ? io_r_141_b : _GEN_14480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14482 = 10'h8e == r_count_19_io_out ? io_r_142_b : _GEN_14481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14483 = 10'h8f == r_count_19_io_out ? io_r_143_b : _GEN_14482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14484 = 10'h90 == r_count_19_io_out ? io_r_144_b : _GEN_14483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14485 = 10'h91 == r_count_19_io_out ? io_r_145_b : _GEN_14484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14486 = 10'h92 == r_count_19_io_out ? io_r_146_b : _GEN_14485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14487 = 10'h93 == r_count_19_io_out ? io_r_147_b : _GEN_14486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14488 = 10'h94 == r_count_19_io_out ? io_r_148_b : _GEN_14487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14489 = 10'h95 == r_count_19_io_out ? io_r_149_b : _GEN_14488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14490 = 10'h96 == r_count_19_io_out ? io_r_150_b : _GEN_14489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14491 = 10'h97 == r_count_19_io_out ? io_r_151_b : _GEN_14490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14492 = 10'h98 == r_count_19_io_out ? io_r_152_b : _GEN_14491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14493 = 10'h99 == r_count_19_io_out ? io_r_153_b : _GEN_14492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14494 = 10'h9a == r_count_19_io_out ? io_r_154_b : _GEN_14493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14495 = 10'h9b == r_count_19_io_out ? io_r_155_b : _GEN_14494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14496 = 10'h9c == r_count_19_io_out ? io_r_156_b : _GEN_14495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14497 = 10'h9d == r_count_19_io_out ? io_r_157_b : _GEN_14496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14498 = 10'h9e == r_count_19_io_out ? io_r_158_b : _GEN_14497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14499 = 10'h9f == r_count_19_io_out ? io_r_159_b : _GEN_14498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14500 = 10'ha0 == r_count_19_io_out ? io_r_160_b : _GEN_14499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14501 = 10'ha1 == r_count_19_io_out ? io_r_161_b : _GEN_14500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14502 = 10'ha2 == r_count_19_io_out ? io_r_162_b : _GEN_14501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14503 = 10'ha3 == r_count_19_io_out ? io_r_163_b : _GEN_14502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14504 = 10'ha4 == r_count_19_io_out ? io_r_164_b : _GEN_14503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14505 = 10'ha5 == r_count_19_io_out ? io_r_165_b : _GEN_14504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14506 = 10'ha6 == r_count_19_io_out ? io_r_166_b : _GEN_14505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14507 = 10'ha7 == r_count_19_io_out ? io_r_167_b : _GEN_14506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14508 = 10'ha8 == r_count_19_io_out ? io_r_168_b : _GEN_14507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14509 = 10'ha9 == r_count_19_io_out ? io_r_169_b : _GEN_14508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14510 = 10'haa == r_count_19_io_out ? io_r_170_b : _GEN_14509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14511 = 10'hab == r_count_19_io_out ? io_r_171_b : _GEN_14510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14512 = 10'hac == r_count_19_io_out ? io_r_172_b : _GEN_14511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14513 = 10'had == r_count_19_io_out ? io_r_173_b : _GEN_14512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14514 = 10'hae == r_count_19_io_out ? io_r_174_b : _GEN_14513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14515 = 10'haf == r_count_19_io_out ? io_r_175_b : _GEN_14514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14516 = 10'hb0 == r_count_19_io_out ? io_r_176_b : _GEN_14515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14517 = 10'hb1 == r_count_19_io_out ? io_r_177_b : _GEN_14516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14518 = 10'hb2 == r_count_19_io_out ? io_r_178_b : _GEN_14517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14519 = 10'hb3 == r_count_19_io_out ? io_r_179_b : _GEN_14518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14520 = 10'hb4 == r_count_19_io_out ? io_r_180_b : _GEN_14519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14521 = 10'hb5 == r_count_19_io_out ? io_r_181_b : _GEN_14520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14522 = 10'hb6 == r_count_19_io_out ? io_r_182_b : _GEN_14521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14523 = 10'hb7 == r_count_19_io_out ? io_r_183_b : _GEN_14522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14524 = 10'hb8 == r_count_19_io_out ? io_r_184_b : _GEN_14523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14525 = 10'hb9 == r_count_19_io_out ? io_r_185_b : _GEN_14524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14526 = 10'hba == r_count_19_io_out ? io_r_186_b : _GEN_14525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14527 = 10'hbb == r_count_19_io_out ? io_r_187_b : _GEN_14526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14528 = 10'hbc == r_count_19_io_out ? io_r_188_b : _GEN_14527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14529 = 10'hbd == r_count_19_io_out ? io_r_189_b : _GEN_14528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14530 = 10'hbe == r_count_19_io_out ? io_r_190_b : _GEN_14529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14531 = 10'hbf == r_count_19_io_out ? io_r_191_b : _GEN_14530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14532 = 10'hc0 == r_count_19_io_out ? io_r_192_b : _GEN_14531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14533 = 10'hc1 == r_count_19_io_out ? io_r_193_b : _GEN_14532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14534 = 10'hc2 == r_count_19_io_out ? io_r_194_b : _GEN_14533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14535 = 10'hc3 == r_count_19_io_out ? io_r_195_b : _GEN_14534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14536 = 10'hc4 == r_count_19_io_out ? io_r_196_b : _GEN_14535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14537 = 10'hc5 == r_count_19_io_out ? io_r_197_b : _GEN_14536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14538 = 10'hc6 == r_count_19_io_out ? io_r_198_b : _GEN_14537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14539 = 10'hc7 == r_count_19_io_out ? io_r_199_b : _GEN_14538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14540 = 10'hc8 == r_count_19_io_out ? io_r_200_b : _GEN_14539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14541 = 10'hc9 == r_count_19_io_out ? io_r_201_b : _GEN_14540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14542 = 10'hca == r_count_19_io_out ? io_r_202_b : _GEN_14541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14543 = 10'hcb == r_count_19_io_out ? io_r_203_b : _GEN_14542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14544 = 10'hcc == r_count_19_io_out ? io_r_204_b : _GEN_14543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14545 = 10'hcd == r_count_19_io_out ? io_r_205_b : _GEN_14544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14546 = 10'hce == r_count_19_io_out ? io_r_206_b : _GEN_14545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14547 = 10'hcf == r_count_19_io_out ? io_r_207_b : _GEN_14546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14548 = 10'hd0 == r_count_19_io_out ? io_r_208_b : _GEN_14547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14549 = 10'hd1 == r_count_19_io_out ? io_r_209_b : _GEN_14548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14550 = 10'hd2 == r_count_19_io_out ? io_r_210_b : _GEN_14549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14551 = 10'hd3 == r_count_19_io_out ? io_r_211_b : _GEN_14550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14552 = 10'hd4 == r_count_19_io_out ? io_r_212_b : _GEN_14551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14553 = 10'hd5 == r_count_19_io_out ? io_r_213_b : _GEN_14552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14554 = 10'hd6 == r_count_19_io_out ? io_r_214_b : _GEN_14553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14555 = 10'hd7 == r_count_19_io_out ? io_r_215_b : _GEN_14554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14556 = 10'hd8 == r_count_19_io_out ? io_r_216_b : _GEN_14555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14557 = 10'hd9 == r_count_19_io_out ? io_r_217_b : _GEN_14556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14558 = 10'hda == r_count_19_io_out ? io_r_218_b : _GEN_14557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14559 = 10'hdb == r_count_19_io_out ? io_r_219_b : _GEN_14558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14560 = 10'hdc == r_count_19_io_out ? io_r_220_b : _GEN_14559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14561 = 10'hdd == r_count_19_io_out ? io_r_221_b : _GEN_14560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14562 = 10'hde == r_count_19_io_out ? io_r_222_b : _GEN_14561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14563 = 10'hdf == r_count_19_io_out ? io_r_223_b : _GEN_14562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14564 = 10'he0 == r_count_19_io_out ? io_r_224_b : _GEN_14563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14565 = 10'he1 == r_count_19_io_out ? io_r_225_b : _GEN_14564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14566 = 10'he2 == r_count_19_io_out ? io_r_226_b : _GEN_14565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14567 = 10'he3 == r_count_19_io_out ? io_r_227_b : _GEN_14566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14568 = 10'he4 == r_count_19_io_out ? io_r_228_b : _GEN_14567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14569 = 10'he5 == r_count_19_io_out ? io_r_229_b : _GEN_14568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14570 = 10'he6 == r_count_19_io_out ? io_r_230_b : _GEN_14569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14571 = 10'he7 == r_count_19_io_out ? io_r_231_b : _GEN_14570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14572 = 10'he8 == r_count_19_io_out ? io_r_232_b : _GEN_14571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14573 = 10'he9 == r_count_19_io_out ? io_r_233_b : _GEN_14572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14574 = 10'hea == r_count_19_io_out ? io_r_234_b : _GEN_14573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14575 = 10'heb == r_count_19_io_out ? io_r_235_b : _GEN_14574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14576 = 10'hec == r_count_19_io_out ? io_r_236_b : _GEN_14575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14577 = 10'hed == r_count_19_io_out ? io_r_237_b : _GEN_14576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14578 = 10'hee == r_count_19_io_out ? io_r_238_b : _GEN_14577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14579 = 10'hef == r_count_19_io_out ? io_r_239_b : _GEN_14578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14580 = 10'hf0 == r_count_19_io_out ? io_r_240_b : _GEN_14579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14581 = 10'hf1 == r_count_19_io_out ? io_r_241_b : _GEN_14580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14582 = 10'hf2 == r_count_19_io_out ? io_r_242_b : _GEN_14581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14583 = 10'hf3 == r_count_19_io_out ? io_r_243_b : _GEN_14582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14584 = 10'hf4 == r_count_19_io_out ? io_r_244_b : _GEN_14583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14585 = 10'hf5 == r_count_19_io_out ? io_r_245_b : _GEN_14584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14586 = 10'hf6 == r_count_19_io_out ? io_r_246_b : _GEN_14585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14587 = 10'hf7 == r_count_19_io_out ? io_r_247_b : _GEN_14586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14588 = 10'hf8 == r_count_19_io_out ? io_r_248_b : _GEN_14587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14589 = 10'hf9 == r_count_19_io_out ? io_r_249_b : _GEN_14588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14590 = 10'hfa == r_count_19_io_out ? io_r_250_b : _GEN_14589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14591 = 10'hfb == r_count_19_io_out ? io_r_251_b : _GEN_14590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14592 = 10'hfc == r_count_19_io_out ? io_r_252_b : _GEN_14591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14593 = 10'hfd == r_count_19_io_out ? io_r_253_b : _GEN_14592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14594 = 10'hfe == r_count_19_io_out ? io_r_254_b : _GEN_14593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14595 = 10'hff == r_count_19_io_out ? io_r_255_b : _GEN_14594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14596 = 10'h100 == r_count_19_io_out ? io_r_256_b : _GEN_14595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14597 = 10'h101 == r_count_19_io_out ? io_r_257_b : _GEN_14596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14598 = 10'h102 == r_count_19_io_out ? io_r_258_b : _GEN_14597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14599 = 10'h103 == r_count_19_io_out ? io_r_259_b : _GEN_14598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14600 = 10'h104 == r_count_19_io_out ? io_r_260_b : _GEN_14599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14601 = 10'h105 == r_count_19_io_out ? io_r_261_b : _GEN_14600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14602 = 10'h106 == r_count_19_io_out ? io_r_262_b : _GEN_14601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14603 = 10'h107 == r_count_19_io_out ? io_r_263_b : _GEN_14602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14604 = 10'h108 == r_count_19_io_out ? io_r_264_b : _GEN_14603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14605 = 10'h109 == r_count_19_io_out ? io_r_265_b : _GEN_14604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14606 = 10'h10a == r_count_19_io_out ? io_r_266_b : _GEN_14605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14607 = 10'h10b == r_count_19_io_out ? io_r_267_b : _GEN_14606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14608 = 10'h10c == r_count_19_io_out ? io_r_268_b : _GEN_14607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14609 = 10'h10d == r_count_19_io_out ? io_r_269_b : _GEN_14608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14610 = 10'h10e == r_count_19_io_out ? io_r_270_b : _GEN_14609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14611 = 10'h10f == r_count_19_io_out ? io_r_271_b : _GEN_14610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14612 = 10'h110 == r_count_19_io_out ? io_r_272_b : _GEN_14611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14613 = 10'h111 == r_count_19_io_out ? io_r_273_b : _GEN_14612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14614 = 10'h112 == r_count_19_io_out ? io_r_274_b : _GEN_14613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14615 = 10'h113 == r_count_19_io_out ? io_r_275_b : _GEN_14614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14616 = 10'h114 == r_count_19_io_out ? io_r_276_b : _GEN_14615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14617 = 10'h115 == r_count_19_io_out ? io_r_277_b : _GEN_14616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14618 = 10'h116 == r_count_19_io_out ? io_r_278_b : _GEN_14617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14619 = 10'h117 == r_count_19_io_out ? io_r_279_b : _GEN_14618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14620 = 10'h118 == r_count_19_io_out ? io_r_280_b : _GEN_14619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14621 = 10'h119 == r_count_19_io_out ? io_r_281_b : _GEN_14620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14622 = 10'h11a == r_count_19_io_out ? io_r_282_b : _GEN_14621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14623 = 10'h11b == r_count_19_io_out ? io_r_283_b : _GEN_14622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14624 = 10'h11c == r_count_19_io_out ? io_r_284_b : _GEN_14623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14625 = 10'h11d == r_count_19_io_out ? io_r_285_b : _GEN_14624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14626 = 10'h11e == r_count_19_io_out ? io_r_286_b : _GEN_14625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14627 = 10'h11f == r_count_19_io_out ? io_r_287_b : _GEN_14626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14628 = 10'h120 == r_count_19_io_out ? io_r_288_b : _GEN_14627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14629 = 10'h121 == r_count_19_io_out ? io_r_289_b : _GEN_14628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14630 = 10'h122 == r_count_19_io_out ? io_r_290_b : _GEN_14629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14631 = 10'h123 == r_count_19_io_out ? io_r_291_b : _GEN_14630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14632 = 10'h124 == r_count_19_io_out ? io_r_292_b : _GEN_14631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14633 = 10'h125 == r_count_19_io_out ? io_r_293_b : _GEN_14632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14634 = 10'h126 == r_count_19_io_out ? io_r_294_b : _GEN_14633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14635 = 10'h127 == r_count_19_io_out ? io_r_295_b : _GEN_14634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14636 = 10'h128 == r_count_19_io_out ? io_r_296_b : _GEN_14635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14637 = 10'h129 == r_count_19_io_out ? io_r_297_b : _GEN_14636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14638 = 10'h12a == r_count_19_io_out ? io_r_298_b : _GEN_14637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14639 = 10'h12b == r_count_19_io_out ? io_r_299_b : _GEN_14638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14640 = 10'h12c == r_count_19_io_out ? io_r_300_b : _GEN_14639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14641 = 10'h12d == r_count_19_io_out ? io_r_301_b : _GEN_14640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14642 = 10'h12e == r_count_19_io_out ? io_r_302_b : _GEN_14641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14643 = 10'h12f == r_count_19_io_out ? io_r_303_b : _GEN_14642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14644 = 10'h130 == r_count_19_io_out ? io_r_304_b : _GEN_14643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14645 = 10'h131 == r_count_19_io_out ? io_r_305_b : _GEN_14644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14646 = 10'h132 == r_count_19_io_out ? io_r_306_b : _GEN_14645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14647 = 10'h133 == r_count_19_io_out ? io_r_307_b : _GEN_14646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14648 = 10'h134 == r_count_19_io_out ? io_r_308_b : _GEN_14647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14649 = 10'h135 == r_count_19_io_out ? io_r_309_b : _GEN_14648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14650 = 10'h136 == r_count_19_io_out ? io_r_310_b : _GEN_14649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14651 = 10'h137 == r_count_19_io_out ? io_r_311_b : _GEN_14650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14652 = 10'h138 == r_count_19_io_out ? io_r_312_b : _GEN_14651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14653 = 10'h139 == r_count_19_io_out ? io_r_313_b : _GEN_14652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14654 = 10'h13a == r_count_19_io_out ? io_r_314_b : _GEN_14653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14655 = 10'h13b == r_count_19_io_out ? io_r_315_b : _GEN_14654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14656 = 10'h13c == r_count_19_io_out ? io_r_316_b : _GEN_14655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14657 = 10'h13d == r_count_19_io_out ? io_r_317_b : _GEN_14656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14658 = 10'h13e == r_count_19_io_out ? io_r_318_b : _GEN_14657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14659 = 10'h13f == r_count_19_io_out ? io_r_319_b : _GEN_14658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14660 = 10'h140 == r_count_19_io_out ? io_r_320_b : _GEN_14659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14661 = 10'h141 == r_count_19_io_out ? io_r_321_b : _GEN_14660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14662 = 10'h142 == r_count_19_io_out ? io_r_322_b : _GEN_14661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14663 = 10'h143 == r_count_19_io_out ? io_r_323_b : _GEN_14662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14664 = 10'h144 == r_count_19_io_out ? io_r_324_b : _GEN_14663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14665 = 10'h145 == r_count_19_io_out ? io_r_325_b : _GEN_14664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14666 = 10'h146 == r_count_19_io_out ? io_r_326_b : _GEN_14665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14667 = 10'h147 == r_count_19_io_out ? io_r_327_b : _GEN_14666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14668 = 10'h148 == r_count_19_io_out ? io_r_328_b : _GEN_14667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14669 = 10'h149 == r_count_19_io_out ? io_r_329_b : _GEN_14668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14670 = 10'h14a == r_count_19_io_out ? io_r_330_b : _GEN_14669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14671 = 10'h14b == r_count_19_io_out ? io_r_331_b : _GEN_14670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14672 = 10'h14c == r_count_19_io_out ? io_r_332_b : _GEN_14671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14673 = 10'h14d == r_count_19_io_out ? io_r_333_b : _GEN_14672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14674 = 10'h14e == r_count_19_io_out ? io_r_334_b : _GEN_14673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14675 = 10'h14f == r_count_19_io_out ? io_r_335_b : _GEN_14674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14676 = 10'h150 == r_count_19_io_out ? io_r_336_b : _GEN_14675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14677 = 10'h151 == r_count_19_io_out ? io_r_337_b : _GEN_14676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14678 = 10'h152 == r_count_19_io_out ? io_r_338_b : _GEN_14677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14679 = 10'h153 == r_count_19_io_out ? io_r_339_b : _GEN_14678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14680 = 10'h154 == r_count_19_io_out ? io_r_340_b : _GEN_14679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14681 = 10'h155 == r_count_19_io_out ? io_r_341_b : _GEN_14680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14682 = 10'h156 == r_count_19_io_out ? io_r_342_b : _GEN_14681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14683 = 10'h157 == r_count_19_io_out ? io_r_343_b : _GEN_14682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14684 = 10'h158 == r_count_19_io_out ? io_r_344_b : _GEN_14683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14685 = 10'h159 == r_count_19_io_out ? io_r_345_b : _GEN_14684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14686 = 10'h15a == r_count_19_io_out ? io_r_346_b : _GEN_14685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14687 = 10'h15b == r_count_19_io_out ? io_r_347_b : _GEN_14686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14688 = 10'h15c == r_count_19_io_out ? io_r_348_b : _GEN_14687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14689 = 10'h15d == r_count_19_io_out ? io_r_349_b : _GEN_14688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14690 = 10'h15e == r_count_19_io_out ? io_r_350_b : _GEN_14689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14691 = 10'h15f == r_count_19_io_out ? io_r_351_b : _GEN_14690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14692 = 10'h160 == r_count_19_io_out ? io_r_352_b : _GEN_14691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14693 = 10'h161 == r_count_19_io_out ? io_r_353_b : _GEN_14692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14694 = 10'h162 == r_count_19_io_out ? io_r_354_b : _GEN_14693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14695 = 10'h163 == r_count_19_io_out ? io_r_355_b : _GEN_14694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14696 = 10'h164 == r_count_19_io_out ? io_r_356_b : _GEN_14695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14697 = 10'h165 == r_count_19_io_out ? io_r_357_b : _GEN_14696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14698 = 10'h166 == r_count_19_io_out ? io_r_358_b : _GEN_14697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14699 = 10'h167 == r_count_19_io_out ? io_r_359_b : _GEN_14698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14700 = 10'h168 == r_count_19_io_out ? io_r_360_b : _GEN_14699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14701 = 10'h169 == r_count_19_io_out ? io_r_361_b : _GEN_14700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14702 = 10'h16a == r_count_19_io_out ? io_r_362_b : _GEN_14701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14703 = 10'h16b == r_count_19_io_out ? io_r_363_b : _GEN_14702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14704 = 10'h16c == r_count_19_io_out ? io_r_364_b : _GEN_14703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14705 = 10'h16d == r_count_19_io_out ? io_r_365_b : _GEN_14704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14706 = 10'h16e == r_count_19_io_out ? io_r_366_b : _GEN_14705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14707 = 10'h16f == r_count_19_io_out ? io_r_367_b : _GEN_14706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14708 = 10'h170 == r_count_19_io_out ? io_r_368_b : _GEN_14707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14709 = 10'h171 == r_count_19_io_out ? io_r_369_b : _GEN_14708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14710 = 10'h172 == r_count_19_io_out ? io_r_370_b : _GEN_14709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14711 = 10'h173 == r_count_19_io_out ? io_r_371_b : _GEN_14710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14712 = 10'h174 == r_count_19_io_out ? io_r_372_b : _GEN_14711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14713 = 10'h175 == r_count_19_io_out ? io_r_373_b : _GEN_14712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14714 = 10'h176 == r_count_19_io_out ? io_r_374_b : _GEN_14713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14715 = 10'h177 == r_count_19_io_out ? io_r_375_b : _GEN_14714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14716 = 10'h178 == r_count_19_io_out ? io_r_376_b : _GEN_14715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14717 = 10'h179 == r_count_19_io_out ? io_r_377_b : _GEN_14716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14718 = 10'h17a == r_count_19_io_out ? io_r_378_b : _GEN_14717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14719 = 10'h17b == r_count_19_io_out ? io_r_379_b : _GEN_14718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14720 = 10'h17c == r_count_19_io_out ? io_r_380_b : _GEN_14719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14721 = 10'h17d == r_count_19_io_out ? io_r_381_b : _GEN_14720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14722 = 10'h17e == r_count_19_io_out ? io_r_382_b : _GEN_14721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14723 = 10'h17f == r_count_19_io_out ? io_r_383_b : _GEN_14722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14724 = 10'h180 == r_count_19_io_out ? io_r_384_b : _GEN_14723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14725 = 10'h181 == r_count_19_io_out ? io_r_385_b : _GEN_14724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14726 = 10'h182 == r_count_19_io_out ? io_r_386_b : _GEN_14725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14727 = 10'h183 == r_count_19_io_out ? io_r_387_b : _GEN_14726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14728 = 10'h184 == r_count_19_io_out ? io_r_388_b : _GEN_14727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14729 = 10'h185 == r_count_19_io_out ? io_r_389_b : _GEN_14728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14730 = 10'h186 == r_count_19_io_out ? io_r_390_b : _GEN_14729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14731 = 10'h187 == r_count_19_io_out ? io_r_391_b : _GEN_14730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14732 = 10'h188 == r_count_19_io_out ? io_r_392_b : _GEN_14731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14733 = 10'h189 == r_count_19_io_out ? io_r_393_b : _GEN_14732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14734 = 10'h18a == r_count_19_io_out ? io_r_394_b : _GEN_14733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14735 = 10'h18b == r_count_19_io_out ? io_r_395_b : _GEN_14734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14736 = 10'h18c == r_count_19_io_out ? io_r_396_b : _GEN_14735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14737 = 10'h18d == r_count_19_io_out ? io_r_397_b : _GEN_14736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14738 = 10'h18e == r_count_19_io_out ? io_r_398_b : _GEN_14737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14739 = 10'h18f == r_count_19_io_out ? io_r_399_b : _GEN_14738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14740 = 10'h190 == r_count_19_io_out ? io_r_400_b : _GEN_14739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14741 = 10'h191 == r_count_19_io_out ? io_r_401_b : _GEN_14740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14742 = 10'h192 == r_count_19_io_out ? io_r_402_b : _GEN_14741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14743 = 10'h193 == r_count_19_io_out ? io_r_403_b : _GEN_14742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14744 = 10'h194 == r_count_19_io_out ? io_r_404_b : _GEN_14743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14745 = 10'h195 == r_count_19_io_out ? io_r_405_b : _GEN_14744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14746 = 10'h196 == r_count_19_io_out ? io_r_406_b : _GEN_14745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14747 = 10'h197 == r_count_19_io_out ? io_r_407_b : _GEN_14746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14748 = 10'h198 == r_count_19_io_out ? io_r_408_b : _GEN_14747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14749 = 10'h199 == r_count_19_io_out ? io_r_409_b : _GEN_14748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14750 = 10'h19a == r_count_19_io_out ? io_r_410_b : _GEN_14749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14751 = 10'h19b == r_count_19_io_out ? io_r_411_b : _GEN_14750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14752 = 10'h19c == r_count_19_io_out ? io_r_412_b : _GEN_14751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14753 = 10'h19d == r_count_19_io_out ? io_r_413_b : _GEN_14752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14754 = 10'h19e == r_count_19_io_out ? io_r_414_b : _GEN_14753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14755 = 10'h19f == r_count_19_io_out ? io_r_415_b : _GEN_14754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14756 = 10'h1a0 == r_count_19_io_out ? io_r_416_b : _GEN_14755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14757 = 10'h1a1 == r_count_19_io_out ? io_r_417_b : _GEN_14756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14758 = 10'h1a2 == r_count_19_io_out ? io_r_418_b : _GEN_14757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14759 = 10'h1a3 == r_count_19_io_out ? io_r_419_b : _GEN_14758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14760 = 10'h1a4 == r_count_19_io_out ? io_r_420_b : _GEN_14759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14761 = 10'h1a5 == r_count_19_io_out ? io_r_421_b : _GEN_14760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14762 = 10'h1a6 == r_count_19_io_out ? io_r_422_b : _GEN_14761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14763 = 10'h1a7 == r_count_19_io_out ? io_r_423_b : _GEN_14762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14764 = 10'h1a8 == r_count_19_io_out ? io_r_424_b : _GEN_14763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14765 = 10'h1a9 == r_count_19_io_out ? io_r_425_b : _GEN_14764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14766 = 10'h1aa == r_count_19_io_out ? io_r_426_b : _GEN_14765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14767 = 10'h1ab == r_count_19_io_out ? io_r_427_b : _GEN_14766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14768 = 10'h1ac == r_count_19_io_out ? io_r_428_b : _GEN_14767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14769 = 10'h1ad == r_count_19_io_out ? io_r_429_b : _GEN_14768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14770 = 10'h1ae == r_count_19_io_out ? io_r_430_b : _GEN_14769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14771 = 10'h1af == r_count_19_io_out ? io_r_431_b : _GEN_14770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14772 = 10'h1b0 == r_count_19_io_out ? io_r_432_b : _GEN_14771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14773 = 10'h1b1 == r_count_19_io_out ? io_r_433_b : _GEN_14772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14774 = 10'h1b2 == r_count_19_io_out ? io_r_434_b : _GEN_14773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14775 = 10'h1b3 == r_count_19_io_out ? io_r_435_b : _GEN_14774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14776 = 10'h1b4 == r_count_19_io_out ? io_r_436_b : _GEN_14775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14777 = 10'h1b5 == r_count_19_io_out ? io_r_437_b : _GEN_14776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14778 = 10'h1b6 == r_count_19_io_out ? io_r_438_b : _GEN_14777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14779 = 10'h1b7 == r_count_19_io_out ? io_r_439_b : _GEN_14778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14780 = 10'h1b8 == r_count_19_io_out ? io_r_440_b : _GEN_14779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14781 = 10'h1b9 == r_count_19_io_out ? io_r_441_b : _GEN_14780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14782 = 10'h1ba == r_count_19_io_out ? io_r_442_b : _GEN_14781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14783 = 10'h1bb == r_count_19_io_out ? io_r_443_b : _GEN_14782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14784 = 10'h1bc == r_count_19_io_out ? io_r_444_b : _GEN_14783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14785 = 10'h1bd == r_count_19_io_out ? io_r_445_b : _GEN_14784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14786 = 10'h1be == r_count_19_io_out ? io_r_446_b : _GEN_14785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14787 = 10'h1bf == r_count_19_io_out ? io_r_447_b : _GEN_14786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14788 = 10'h1c0 == r_count_19_io_out ? io_r_448_b : _GEN_14787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14789 = 10'h1c1 == r_count_19_io_out ? io_r_449_b : _GEN_14788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14790 = 10'h1c2 == r_count_19_io_out ? io_r_450_b : _GEN_14789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14791 = 10'h1c3 == r_count_19_io_out ? io_r_451_b : _GEN_14790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14792 = 10'h1c4 == r_count_19_io_out ? io_r_452_b : _GEN_14791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14793 = 10'h1c5 == r_count_19_io_out ? io_r_453_b : _GEN_14792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14794 = 10'h1c6 == r_count_19_io_out ? io_r_454_b : _GEN_14793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14795 = 10'h1c7 == r_count_19_io_out ? io_r_455_b : _GEN_14794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14796 = 10'h1c8 == r_count_19_io_out ? io_r_456_b : _GEN_14795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14797 = 10'h1c9 == r_count_19_io_out ? io_r_457_b : _GEN_14796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14798 = 10'h1ca == r_count_19_io_out ? io_r_458_b : _GEN_14797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14799 = 10'h1cb == r_count_19_io_out ? io_r_459_b : _GEN_14798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14800 = 10'h1cc == r_count_19_io_out ? io_r_460_b : _GEN_14799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14801 = 10'h1cd == r_count_19_io_out ? io_r_461_b : _GEN_14800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14802 = 10'h1ce == r_count_19_io_out ? io_r_462_b : _GEN_14801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14803 = 10'h1cf == r_count_19_io_out ? io_r_463_b : _GEN_14802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14804 = 10'h1d0 == r_count_19_io_out ? io_r_464_b : _GEN_14803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14805 = 10'h1d1 == r_count_19_io_out ? io_r_465_b : _GEN_14804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14806 = 10'h1d2 == r_count_19_io_out ? io_r_466_b : _GEN_14805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14807 = 10'h1d3 == r_count_19_io_out ? io_r_467_b : _GEN_14806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14808 = 10'h1d4 == r_count_19_io_out ? io_r_468_b : _GEN_14807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14809 = 10'h1d5 == r_count_19_io_out ? io_r_469_b : _GEN_14808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14810 = 10'h1d6 == r_count_19_io_out ? io_r_470_b : _GEN_14809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14811 = 10'h1d7 == r_count_19_io_out ? io_r_471_b : _GEN_14810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14812 = 10'h1d8 == r_count_19_io_out ? io_r_472_b : _GEN_14811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14813 = 10'h1d9 == r_count_19_io_out ? io_r_473_b : _GEN_14812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14814 = 10'h1da == r_count_19_io_out ? io_r_474_b : _GEN_14813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14815 = 10'h1db == r_count_19_io_out ? io_r_475_b : _GEN_14814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14816 = 10'h1dc == r_count_19_io_out ? io_r_476_b : _GEN_14815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14817 = 10'h1dd == r_count_19_io_out ? io_r_477_b : _GEN_14816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14818 = 10'h1de == r_count_19_io_out ? io_r_478_b : _GEN_14817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14819 = 10'h1df == r_count_19_io_out ? io_r_479_b : _GEN_14818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14820 = 10'h1e0 == r_count_19_io_out ? io_r_480_b : _GEN_14819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14821 = 10'h1e1 == r_count_19_io_out ? io_r_481_b : _GEN_14820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14822 = 10'h1e2 == r_count_19_io_out ? io_r_482_b : _GEN_14821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14823 = 10'h1e3 == r_count_19_io_out ? io_r_483_b : _GEN_14822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14824 = 10'h1e4 == r_count_19_io_out ? io_r_484_b : _GEN_14823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14825 = 10'h1e5 == r_count_19_io_out ? io_r_485_b : _GEN_14824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14826 = 10'h1e6 == r_count_19_io_out ? io_r_486_b : _GEN_14825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14827 = 10'h1e7 == r_count_19_io_out ? io_r_487_b : _GEN_14826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14828 = 10'h1e8 == r_count_19_io_out ? io_r_488_b : _GEN_14827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14829 = 10'h1e9 == r_count_19_io_out ? io_r_489_b : _GEN_14828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14830 = 10'h1ea == r_count_19_io_out ? io_r_490_b : _GEN_14829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14831 = 10'h1eb == r_count_19_io_out ? io_r_491_b : _GEN_14830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14832 = 10'h1ec == r_count_19_io_out ? io_r_492_b : _GEN_14831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14833 = 10'h1ed == r_count_19_io_out ? io_r_493_b : _GEN_14832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14834 = 10'h1ee == r_count_19_io_out ? io_r_494_b : _GEN_14833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14835 = 10'h1ef == r_count_19_io_out ? io_r_495_b : _GEN_14834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14836 = 10'h1f0 == r_count_19_io_out ? io_r_496_b : _GEN_14835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14837 = 10'h1f1 == r_count_19_io_out ? io_r_497_b : _GEN_14836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14838 = 10'h1f2 == r_count_19_io_out ? io_r_498_b : _GEN_14837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14839 = 10'h1f3 == r_count_19_io_out ? io_r_499_b : _GEN_14838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14840 = 10'h1f4 == r_count_19_io_out ? io_r_500_b : _GEN_14839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14841 = 10'h1f5 == r_count_19_io_out ? io_r_501_b : _GEN_14840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14842 = 10'h1f6 == r_count_19_io_out ? io_r_502_b : _GEN_14841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14843 = 10'h1f7 == r_count_19_io_out ? io_r_503_b : _GEN_14842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14844 = 10'h1f8 == r_count_19_io_out ? io_r_504_b : _GEN_14843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14845 = 10'h1f9 == r_count_19_io_out ? io_r_505_b : _GEN_14844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14846 = 10'h1fa == r_count_19_io_out ? io_r_506_b : _GEN_14845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14847 = 10'h1fb == r_count_19_io_out ? io_r_507_b : _GEN_14846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14848 = 10'h1fc == r_count_19_io_out ? io_r_508_b : _GEN_14847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14849 = 10'h1fd == r_count_19_io_out ? io_r_509_b : _GEN_14848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14850 = 10'h1fe == r_count_19_io_out ? io_r_510_b : _GEN_14849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14851 = 10'h1ff == r_count_19_io_out ? io_r_511_b : _GEN_14850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14852 = 10'h200 == r_count_19_io_out ? io_r_512_b : _GEN_14851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14853 = 10'h201 == r_count_19_io_out ? io_r_513_b : _GEN_14852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14854 = 10'h202 == r_count_19_io_out ? io_r_514_b : _GEN_14853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14855 = 10'h203 == r_count_19_io_out ? io_r_515_b : _GEN_14854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14856 = 10'h204 == r_count_19_io_out ? io_r_516_b : _GEN_14855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14857 = 10'h205 == r_count_19_io_out ? io_r_517_b : _GEN_14856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14858 = 10'h206 == r_count_19_io_out ? io_r_518_b : _GEN_14857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14859 = 10'h207 == r_count_19_io_out ? io_r_519_b : _GEN_14858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14860 = 10'h208 == r_count_19_io_out ? io_r_520_b : _GEN_14859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14861 = 10'h209 == r_count_19_io_out ? io_r_521_b : _GEN_14860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14862 = 10'h20a == r_count_19_io_out ? io_r_522_b : _GEN_14861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14863 = 10'h20b == r_count_19_io_out ? io_r_523_b : _GEN_14862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14864 = 10'h20c == r_count_19_io_out ? io_r_524_b : _GEN_14863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14865 = 10'h20d == r_count_19_io_out ? io_r_525_b : _GEN_14864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14866 = 10'h20e == r_count_19_io_out ? io_r_526_b : _GEN_14865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14867 = 10'h20f == r_count_19_io_out ? io_r_527_b : _GEN_14866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14868 = 10'h210 == r_count_19_io_out ? io_r_528_b : _GEN_14867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14869 = 10'h211 == r_count_19_io_out ? io_r_529_b : _GEN_14868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14870 = 10'h212 == r_count_19_io_out ? io_r_530_b : _GEN_14869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14871 = 10'h213 == r_count_19_io_out ? io_r_531_b : _GEN_14870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14872 = 10'h214 == r_count_19_io_out ? io_r_532_b : _GEN_14871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14873 = 10'h215 == r_count_19_io_out ? io_r_533_b : _GEN_14872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14874 = 10'h216 == r_count_19_io_out ? io_r_534_b : _GEN_14873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14875 = 10'h217 == r_count_19_io_out ? io_r_535_b : _GEN_14874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14876 = 10'h218 == r_count_19_io_out ? io_r_536_b : _GEN_14875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14877 = 10'h219 == r_count_19_io_out ? io_r_537_b : _GEN_14876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14878 = 10'h21a == r_count_19_io_out ? io_r_538_b : _GEN_14877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14879 = 10'h21b == r_count_19_io_out ? io_r_539_b : _GEN_14878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14880 = 10'h21c == r_count_19_io_out ? io_r_540_b : _GEN_14879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14881 = 10'h21d == r_count_19_io_out ? io_r_541_b : _GEN_14880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14882 = 10'h21e == r_count_19_io_out ? io_r_542_b : _GEN_14881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14883 = 10'h21f == r_count_19_io_out ? io_r_543_b : _GEN_14882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14884 = 10'h220 == r_count_19_io_out ? io_r_544_b : _GEN_14883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14885 = 10'h221 == r_count_19_io_out ? io_r_545_b : _GEN_14884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14886 = 10'h222 == r_count_19_io_out ? io_r_546_b : _GEN_14885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14887 = 10'h223 == r_count_19_io_out ? io_r_547_b : _GEN_14886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14888 = 10'h224 == r_count_19_io_out ? io_r_548_b : _GEN_14887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14889 = 10'h225 == r_count_19_io_out ? io_r_549_b : _GEN_14888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14890 = 10'h226 == r_count_19_io_out ? io_r_550_b : _GEN_14889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14891 = 10'h227 == r_count_19_io_out ? io_r_551_b : _GEN_14890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14892 = 10'h228 == r_count_19_io_out ? io_r_552_b : _GEN_14891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14893 = 10'h229 == r_count_19_io_out ? io_r_553_b : _GEN_14892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14894 = 10'h22a == r_count_19_io_out ? io_r_554_b : _GEN_14893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14895 = 10'h22b == r_count_19_io_out ? io_r_555_b : _GEN_14894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14896 = 10'h22c == r_count_19_io_out ? io_r_556_b : _GEN_14895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14897 = 10'h22d == r_count_19_io_out ? io_r_557_b : _GEN_14896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14898 = 10'h22e == r_count_19_io_out ? io_r_558_b : _GEN_14897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14899 = 10'h22f == r_count_19_io_out ? io_r_559_b : _GEN_14898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14900 = 10'h230 == r_count_19_io_out ? io_r_560_b : _GEN_14899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14901 = 10'h231 == r_count_19_io_out ? io_r_561_b : _GEN_14900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14902 = 10'h232 == r_count_19_io_out ? io_r_562_b : _GEN_14901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14903 = 10'h233 == r_count_19_io_out ? io_r_563_b : _GEN_14902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14904 = 10'h234 == r_count_19_io_out ? io_r_564_b : _GEN_14903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14905 = 10'h235 == r_count_19_io_out ? io_r_565_b : _GEN_14904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14906 = 10'h236 == r_count_19_io_out ? io_r_566_b : _GEN_14905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14907 = 10'h237 == r_count_19_io_out ? io_r_567_b : _GEN_14906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14908 = 10'h238 == r_count_19_io_out ? io_r_568_b : _GEN_14907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14909 = 10'h239 == r_count_19_io_out ? io_r_569_b : _GEN_14908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14910 = 10'h23a == r_count_19_io_out ? io_r_570_b : _GEN_14909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14911 = 10'h23b == r_count_19_io_out ? io_r_571_b : _GEN_14910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14912 = 10'h23c == r_count_19_io_out ? io_r_572_b : _GEN_14911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14913 = 10'h23d == r_count_19_io_out ? io_r_573_b : _GEN_14912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14914 = 10'h23e == r_count_19_io_out ? io_r_574_b : _GEN_14913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14915 = 10'h23f == r_count_19_io_out ? io_r_575_b : _GEN_14914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14916 = 10'h240 == r_count_19_io_out ? io_r_576_b : _GEN_14915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14917 = 10'h241 == r_count_19_io_out ? io_r_577_b : _GEN_14916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14918 = 10'h242 == r_count_19_io_out ? io_r_578_b : _GEN_14917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14919 = 10'h243 == r_count_19_io_out ? io_r_579_b : _GEN_14918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14920 = 10'h244 == r_count_19_io_out ? io_r_580_b : _GEN_14919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14921 = 10'h245 == r_count_19_io_out ? io_r_581_b : _GEN_14920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14922 = 10'h246 == r_count_19_io_out ? io_r_582_b : _GEN_14921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14923 = 10'h247 == r_count_19_io_out ? io_r_583_b : _GEN_14922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14924 = 10'h248 == r_count_19_io_out ? io_r_584_b : _GEN_14923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14925 = 10'h249 == r_count_19_io_out ? io_r_585_b : _GEN_14924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14926 = 10'h24a == r_count_19_io_out ? io_r_586_b : _GEN_14925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14927 = 10'h24b == r_count_19_io_out ? io_r_587_b : _GEN_14926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14928 = 10'h24c == r_count_19_io_out ? io_r_588_b : _GEN_14927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14929 = 10'h24d == r_count_19_io_out ? io_r_589_b : _GEN_14928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14930 = 10'h24e == r_count_19_io_out ? io_r_590_b : _GEN_14929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14931 = 10'h24f == r_count_19_io_out ? io_r_591_b : _GEN_14930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14932 = 10'h250 == r_count_19_io_out ? io_r_592_b : _GEN_14931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14933 = 10'h251 == r_count_19_io_out ? io_r_593_b : _GEN_14932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14934 = 10'h252 == r_count_19_io_out ? io_r_594_b : _GEN_14933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14935 = 10'h253 == r_count_19_io_out ? io_r_595_b : _GEN_14934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14936 = 10'h254 == r_count_19_io_out ? io_r_596_b : _GEN_14935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14937 = 10'h255 == r_count_19_io_out ? io_r_597_b : _GEN_14936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14938 = 10'h256 == r_count_19_io_out ? io_r_598_b : _GEN_14937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14939 = 10'h257 == r_count_19_io_out ? io_r_599_b : _GEN_14938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14940 = 10'h258 == r_count_19_io_out ? io_r_600_b : _GEN_14939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14941 = 10'h259 == r_count_19_io_out ? io_r_601_b : _GEN_14940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14942 = 10'h25a == r_count_19_io_out ? io_r_602_b : _GEN_14941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14943 = 10'h25b == r_count_19_io_out ? io_r_603_b : _GEN_14942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14944 = 10'h25c == r_count_19_io_out ? io_r_604_b : _GEN_14943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14945 = 10'h25d == r_count_19_io_out ? io_r_605_b : _GEN_14944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14946 = 10'h25e == r_count_19_io_out ? io_r_606_b : _GEN_14945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14947 = 10'h25f == r_count_19_io_out ? io_r_607_b : _GEN_14946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14948 = 10'h260 == r_count_19_io_out ? io_r_608_b : _GEN_14947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14949 = 10'h261 == r_count_19_io_out ? io_r_609_b : _GEN_14948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14950 = 10'h262 == r_count_19_io_out ? io_r_610_b : _GEN_14949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14951 = 10'h263 == r_count_19_io_out ? io_r_611_b : _GEN_14950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14952 = 10'h264 == r_count_19_io_out ? io_r_612_b : _GEN_14951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14953 = 10'h265 == r_count_19_io_out ? io_r_613_b : _GEN_14952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14954 = 10'h266 == r_count_19_io_out ? io_r_614_b : _GEN_14953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14955 = 10'h267 == r_count_19_io_out ? io_r_615_b : _GEN_14954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14956 = 10'h268 == r_count_19_io_out ? io_r_616_b : _GEN_14955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14957 = 10'h269 == r_count_19_io_out ? io_r_617_b : _GEN_14956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14958 = 10'h26a == r_count_19_io_out ? io_r_618_b : _GEN_14957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14959 = 10'h26b == r_count_19_io_out ? io_r_619_b : _GEN_14958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14960 = 10'h26c == r_count_19_io_out ? io_r_620_b : _GEN_14959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14961 = 10'h26d == r_count_19_io_out ? io_r_621_b : _GEN_14960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14962 = 10'h26e == r_count_19_io_out ? io_r_622_b : _GEN_14961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14963 = 10'h26f == r_count_19_io_out ? io_r_623_b : _GEN_14962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14964 = 10'h270 == r_count_19_io_out ? io_r_624_b : _GEN_14963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14965 = 10'h271 == r_count_19_io_out ? io_r_625_b : _GEN_14964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14966 = 10'h272 == r_count_19_io_out ? io_r_626_b : _GEN_14965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14967 = 10'h273 == r_count_19_io_out ? io_r_627_b : _GEN_14966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14968 = 10'h274 == r_count_19_io_out ? io_r_628_b : _GEN_14967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14969 = 10'h275 == r_count_19_io_out ? io_r_629_b : _GEN_14968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14970 = 10'h276 == r_count_19_io_out ? io_r_630_b : _GEN_14969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14971 = 10'h277 == r_count_19_io_out ? io_r_631_b : _GEN_14970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14972 = 10'h278 == r_count_19_io_out ? io_r_632_b : _GEN_14971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14973 = 10'h279 == r_count_19_io_out ? io_r_633_b : _GEN_14972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14974 = 10'h27a == r_count_19_io_out ? io_r_634_b : _GEN_14973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14975 = 10'h27b == r_count_19_io_out ? io_r_635_b : _GEN_14974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14976 = 10'h27c == r_count_19_io_out ? io_r_636_b : _GEN_14975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14977 = 10'h27d == r_count_19_io_out ? io_r_637_b : _GEN_14976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14978 = 10'h27e == r_count_19_io_out ? io_r_638_b : _GEN_14977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14979 = 10'h27f == r_count_19_io_out ? io_r_639_b : _GEN_14978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14980 = 10'h280 == r_count_19_io_out ? io_r_640_b : _GEN_14979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14981 = 10'h281 == r_count_19_io_out ? io_r_641_b : _GEN_14980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14982 = 10'h282 == r_count_19_io_out ? io_r_642_b : _GEN_14981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14983 = 10'h283 == r_count_19_io_out ? io_r_643_b : _GEN_14982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14984 = 10'h284 == r_count_19_io_out ? io_r_644_b : _GEN_14983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14985 = 10'h285 == r_count_19_io_out ? io_r_645_b : _GEN_14984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14986 = 10'h286 == r_count_19_io_out ? io_r_646_b : _GEN_14985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14987 = 10'h287 == r_count_19_io_out ? io_r_647_b : _GEN_14986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14988 = 10'h288 == r_count_19_io_out ? io_r_648_b : _GEN_14987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14989 = 10'h289 == r_count_19_io_out ? io_r_649_b : _GEN_14988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14990 = 10'h28a == r_count_19_io_out ? io_r_650_b : _GEN_14989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14991 = 10'h28b == r_count_19_io_out ? io_r_651_b : _GEN_14990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14992 = 10'h28c == r_count_19_io_out ? io_r_652_b : _GEN_14991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14993 = 10'h28d == r_count_19_io_out ? io_r_653_b : _GEN_14992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14994 = 10'h28e == r_count_19_io_out ? io_r_654_b : _GEN_14993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14995 = 10'h28f == r_count_19_io_out ? io_r_655_b : _GEN_14994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14996 = 10'h290 == r_count_19_io_out ? io_r_656_b : _GEN_14995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14997 = 10'h291 == r_count_19_io_out ? io_r_657_b : _GEN_14996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14998 = 10'h292 == r_count_19_io_out ? io_r_658_b : _GEN_14997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14999 = 10'h293 == r_count_19_io_out ? io_r_659_b : _GEN_14998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15000 = 10'h294 == r_count_19_io_out ? io_r_660_b : _GEN_14999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15001 = 10'h295 == r_count_19_io_out ? io_r_661_b : _GEN_15000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15002 = 10'h296 == r_count_19_io_out ? io_r_662_b : _GEN_15001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15003 = 10'h297 == r_count_19_io_out ? io_r_663_b : _GEN_15002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15004 = 10'h298 == r_count_19_io_out ? io_r_664_b : _GEN_15003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15005 = 10'h299 == r_count_19_io_out ? io_r_665_b : _GEN_15004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15006 = 10'h29a == r_count_19_io_out ? io_r_666_b : _GEN_15005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15007 = 10'h29b == r_count_19_io_out ? io_r_667_b : _GEN_15006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15008 = 10'h29c == r_count_19_io_out ? io_r_668_b : _GEN_15007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15009 = 10'h29d == r_count_19_io_out ? io_r_669_b : _GEN_15008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15010 = 10'h29e == r_count_19_io_out ? io_r_670_b : _GEN_15009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15011 = 10'h29f == r_count_19_io_out ? io_r_671_b : _GEN_15010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15012 = 10'h2a0 == r_count_19_io_out ? io_r_672_b : _GEN_15011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15013 = 10'h2a1 == r_count_19_io_out ? io_r_673_b : _GEN_15012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15014 = 10'h2a2 == r_count_19_io_out ? io_r_674_b : _GEN_15013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15015 = 10'h2a3 == r_count_19_io_out ? io_r_675_b : _GEN_15014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15016 = 10'h2a4 == r_count_19_io_out ? io_r_676_b : _GEN_15015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15017 = 10'h2a5 == r_count_19_io_out ? io_r_677_b : _GEN_15016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15018 = 10'h2a6 == r_count_19_io_out ? io_r_678_b : _GEN_15017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15019 = 10'h2a7 == r_count_19_io_out ? io_r_679_b : _GEN_15018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15020 = 10'h2a8 == r_count_19_io_out ? io_r_680_b : _GEN_15019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15021 = 10'h2a9 == r_count_19_io_out ? io_r_681_b : _GEN_15020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15022 = 10'h2aa == r_count_19_io_out ? io_r_682_b : _GEN_15021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15023 = 10'h2ab == r_count_19_io_out ? io_r_683_b : _GEN_15022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15024 = 10'h2ac == r_count_19_io_out ? io_r_684_b : _GEN_15023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15025 = 10'h2ad == r_count_19_io_out ? io_r_685_b : _GEN_15024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15026 = 10'h2ae == r_count_19_io_out ? io_r_686_b : _GEN_15025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15027 = 10'h2af == r_count_19_io_out ? io_r_687_b : _GEN_15026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15028 = 10'h2b0 == r_count_19_io_out ? io_r_688_b : _GEN_15027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15029 = 10'h2b1 == r_count_19_io_out ? io_r_689_b : _GEN_15028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15030 = 10'h2b2 == r_count_19_io_out ? io_r_690_b : _GEN_15029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15031 = 10'h2b3 == r_count_19_io_out ? io_r_691_b : _GEN_15030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15032 = 10'h2b4 == r_count_19_io_out ? io_r_692_b : _GEN_15031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15033 = 10'h2b5 == r_count_19_io_out ? io_r_693_b : _GEN_15032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15034 = 10'h2b6 == r_count_19_io_out ? io_r_694_b : _GEN_15033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15035 = 10'h2b7 == r_count_19_io_out ? io_r_695_b : _GEN_15034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15036 = 10'h2b8 == r_count_19_io_out ? io_r_696_b : _GEN_15035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15037 = 10'h2b9 == r_count_19_io_out ? io_r_697_b : _GEN_15036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15038 = 10'h2ba == r_count_19_io_out ? io_r_698_b : _GEN_15037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15039 = 10'h2bb == r_count_19_io_out ? io_r_699_b : _GEN_15038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15040 = 10'h2bc == r_count_19_io_out ? io_r_700_b : _GEN_15039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15041 = 10'h2bd == r_count_19_io_out ? io_r_701_b : _GEN_15040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15042 = 10'h2be == r_count_19_io_out ? io_r_702_b : _GEN_15041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15043 = 10'h2bf == r_count_19_io_out ? io_r_703_b : _GEN_15042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15044 = 10'h2c0 == r_count_19_io_out ? io_r_704_b : _GEN_15043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15045 = 10'h2c1 == r_count_19_io_out ? io_r_705_b : _GEN_15044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15046 = 10'h2c2 == r_count_19_io_out ? io_r_706_b : _GEN_15045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15047 = 10'h2c3 == r_count_19_io_out ? io_r_707_b : _GEN_15046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15048 = 10'h2c4 == r_count_19_io_out ? io_r_708_b : _GEN_15047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15049 = 10'h2c5 == r_count_19_io_out ? io_r_709_b : _GEN_15048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15050 = 10'h2c6 == r_count_19_io_out ? io_r_710_b : _GEN_15049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15051 = 10'h2c7 == r_count_19_io_out ? io_r_711_b : _GEN_15050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15052 = 10'h2c8 == r_count_19_io_out ? io_r_712_b : _GEN_15051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15053 = 10'h2c9 == r_count_19_io_out ? io_r_713_b : _GEN_15052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15054 = 10'h2ca == r_count_19_io_out ? io_r_714_b : _GEN_15053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15055 = 10'h2cb == r_count_19_io_out ? io_r_715_b : _GEN_15054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15056 = 10'h2cc == r_count_19_io_out ? io_r_716_b : _GEN_15055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15057 = 10'h2cd == r_count_19_io_out ? io_r_717_b : _GEN_15056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15058 = 10'h2ce == r_count_19_io_out ? io_r_718_b : _GEN_15057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15059 = 10'h2cf == r_count_19_io_out ? io_r_719_b : _GEN_15058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15060 = 10'h2d0 == r_count_19_io_out ? io_r_720_b : _GEN_15059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15061 = 10'h2d1 == r_count_19_io_out ? io_r_721_b : _GEN_15060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15062 = 10'h2d2 == r_count_19_io_out ? io_r_722_b : _GEN_15061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15063 = 10'h2d3 == r_count_19_io_out ? io_r_723_b : _GEN_15062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15064 = 10'h2d4 == r_count_19_io_out ? io_r_724_b : _GEN_15063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15065 = 10'h2d5 == r_count_19_io_out ? io_r_725_b : _GEN_15064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15066 = 10'h2d6 == r_count_19_io_out ? io_r_726_b : _GEN_15065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15067 = 10'h2d7 == r_count_19_io_out ? io_r_727_b : _GEN_15066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15068 = 10'h2d8 == r_count_19_io_out ? io_r_728_b : _GEN_15067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15069 = 10'h2d9 == r_count_19_io_out ? io_r_729_b : _GEN_15068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15070 = 10'h2da == r_count_19_io_out ? io_r_730_b : _GEN_15069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15071 = 10'h2db == r_count_19_io_out ? io_r_731_b : _GEN_15070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15072 = 10'h2dc == r_count_19_io_out ? io_r_732_b : _GEN_15071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15073 = 10'h2dd == r_count_19_io_out ? io_r_733_b : _GEN_15072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15074 = 10'h2de == r_count_19_io_out ? io_r_734_b : _GEN_15073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15075 = 10'h2df == r_count_19_io_out ? io_r_735_b : _GEN_15074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15076 = 10'h2e0 == r_count_19_io_out ? io_r_736_b : _GEN_15075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15077 = 10'h2e1 == r_count_19_io_out ? io_r_737_b : _GEN_15076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15078 = 10'h2e2 == r_count_19_io_out ? io_r_738_b : _GEN_15077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15079 = 10'h2e3 == r_count_19_io_out ? io_r_739_b : _GEN_15078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15080 = 10'h2e4 == r_count_19_io_out ? io_r_740_b : _GEN_15079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15081 = 10'h2e5 == r_count_19_io_out ? io_r_741_b : _GEN_15080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15082 = 10'h2e6 == r_count_19_io_out ? io_r_742_b : _GEN_15081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15083 = 10'h2e7 == r_count_19_io_out ? io_r_743_b : _GEN_15082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15084 = 10'h2e8 == r_count_19_io_out ? io_r_744_b : _GEN_15083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15085 = 10'h2e9 == r_count_19_io_out ? io_r_745_b : _GEN_15084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15086 = 10'h2ea == r_count_19_io_out ? io_r_746_b : _GEN_15085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15087 = 10'h2eb == r_count_19_io_out ? io_r_747_b : _GEN_15086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15088 = 10'h2ec == r_count_19_io_out ? io_r_748_b : _GEN_15087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15091 = 10'h1 == r_count_20_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15092 = 10'h2 == r_count_20_io_out ? io_r_2_b : _GEN_15091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15093 = 10'h3 == r_count_20_io_out ? io_r_3_b : _GEN_15092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15094 = 10'h4 == r_count_20_io_out ? io_r_4_b : _GEN_15093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15095 = 10'h5 == r_count_20_io_out ? io_r_5_b : _GEN_15094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15096 = 10'h6 == r_count_20_io_out ? io_r_6_b : _GEN_15095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15097 = 10'h7 == r_count_20_io_out ? io_r_7_b : _GEN_15096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15098 = 10'h8 == r_count_20_io_out ? io_r_8_b : _GEN_15097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15099 = 10'h9 == r_count_20_io_out ? io_r_9_b : _GEN_15098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15100 = 10'ha == r_count_20_io_out ? io_r_10_b : _GEN_15099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15101 = 10'hb == r_count_20_io_out ? io_r_11_b : _GEN_15100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15102 = 10'hc == r_count_20_io_out ? io_r_12_b : _GEN_15101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15103 = 10'hd == r_count_20_io_out ? io_r_13_b : _GEN_15102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15104 = 10'he == r_count_20_io_out ? io_r_14_b : _GEN_15103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15105 = 10'hf == r_count_20_io_out ? io_r_15_b : _GEN_15104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15106 = 10'h10 == r_count_20_io_out ? io_r_16_b : _GEN_15105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15107 = 10'h11 == r_count_20_io_out ? io_r_17_b : _GEN_15106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15108 = 10'h12 == r_count_20_io_out ? io_r_18_b : _GEN_15107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15109 = 10'h13 == r_count_20_io_out ? io_r_19_b : _GEN_15108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15110 = 10'h14 == r_count_20_io_out ? io_r_20_b : _GEN_15109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15111 = 10'h15 == r_count_20_io_out ? io_r_21_b : _GEN_15110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15112 = 10'h16 == r_count_20_io_out ? io_r_22_b : _GEN_15111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15113 = 10'h17 == r_count_20_io_out ? io_r_23_b : _GEN_15112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15114 = 10'h18 == r_count_20_io_out ? io_r_24_b : _GEN_15113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15115 = 10'h19 == r_count_20_io_out ? io_r_25_b : _GEN_15114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15116 = 10'h1a == r_count_20_io_out ? io_r_26_b : _GEN_15115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15117 = 10'h1b == r_count_20_io_out ? io_r_27_b : _GEN_15116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15118 = 10'h1c == r_count_20_io_out ? io_r_28_b : _GEN_15117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15119 = 10'h1d == r_count_20_io_out ? io_r_29_b : _GEN_15118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15120 = 10'h1e == r_count_20_io_out ? io_r_30_b : _GEN_15119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15121 = 10'h1f == r_count_20_io_out ? io_r_31_b : _GEN_15120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15122 = 10'h20 == r_count_20_io_out ? io_r_32_b : _GEN_15121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15123 = 10'h21 == r_count_20_io_out ? io_r_33_b : _GEN_15122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15124 = 10'h22 == r_count_20_io_out ? io_r_34_b : _GEN_15123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15125 = 10'h23 == r_count_20_io_out ? io_r_35_b : _GEN_15124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15126 = 10'h24 == r_count_20_io_out ? io_r_36_b : _GEN_15125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15127 = 10'h25 == r_count_20_io_out ? io_r_37_b : _GEN_15126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15128 = 10'h26 == r_count_20_io_out ? io_r_38_b : _GEN_15127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15129 = 10'h27 == r_count_20_io_out ? io_r_39_b : _GEN_15128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15130 = 10'h28 == r_count_20_io_out ? io_r_40_b : _GEN_15129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15131 = 10'h29 == r_count_20_io_out ? io_r_41_b : _GEN_15130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15132 = 10'h2a == r_count_20_io_out ? io_r_42_b : _GEN_15131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15133 = 10'h2b == r_count_20_io_out ? io_r_43_b : _GEN_15132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15134 = 10'h2c == r_count_20_io_out ? io_r_44_b : _GEN_15133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15135 = 10'h2d == r_count_20_io_out ? io_r_45_b : _GEN_15134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15136 = 10'h2e == r_count_20_io_out ? io_r_46_b : _GEN_15135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15137 = 10'h2f == r_count_20_io_out ? io_r_47_b : _GEN_15136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15138 = 10'h30 == r_count_20_io_out ? io_r_48_b : _GEN_15137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15139 = 10'h31 == r_count_20_io_out ? io_r_49_b : _GEN_15138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15140 = 10'h32 == r_count_20_io_out ? io_r_50_b : _GEN_15139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15141 = 10'h33 == r_count_20_io_out ? io_r_51_b : _GEN_15140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15142 = 10'h34 == r_count_20_io_out ? io_r_52_b : _GEN_15141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15143 = 10'h35 == r_count_20_io_out ? io_r_53_b : _GEN_15142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15144 = 10'h36 == r_count_20_io_out ? io_r_54_b : _GEN_15143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15145 = 10'h37 == r_count_20_io_out ? io_r_55_b : _GEN_15144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15146 = 10'h38 == r_count_20_io_out ? io_r_56_b : _GEN_15145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15147 = 10'h39 == r_count_20_io_out ? io_r_57_b : _GEN_15146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15148 = 10'h3a == r_count_20_io_out ? io_r_58_b : _GEN_15147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15149 = 10'h3b == r_count_20_io_out ? io_r_59_b : _GEN_15148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15150 = 10'h3c == r_count_20_io_out ? io_r_60_b : _GEN_15149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15151 = 10'h3d == r_count_20_io_out ? io_r_61_b : _GEN_15150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15152 = 10'h3e == r_count_20_io_out ? io_r_62_b : _GEN_15151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15153 = 10'h3f == r_count_20_io_out ? io_r_63_b : _GEN_15152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15154 = 10'h40 == r_count_20_io_out ? io_r_64_b : _GEN_15153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15155 = 10'h41 == r_count_20_io_out ? io_r_65_b : _GEN_15154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15156 = 10'h42 == r_count_20_io_out ? io_r_66_b : _GEN_15155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15157 = 10'h43 == r_count_20_io_out ? io_r_67_b : _GEN_15156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15158 = 10'h44 == r_count_20_io_out ? io_r_68_b : _GEN_15157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15159 = 10'h45 == r_count_20_io_out ? io_r_69_b : _GEN_15158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15160 = 10'h46 == r_count_20_io_out ? io_r_70_b : _GEN_15159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15161 = 10'h47 == r_count_20_io_out ? io_r_71_b : _GEN_15160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15162 = 10'h48 == r_count_20_io_out ? io_r_72_b : _GEN_15161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15163 = 10'h49 == r_count_20_io_out ? io_r_73_b : _GEN_15162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15164 = 10'h4a == r_count_20_io_out ? io_r_74_b : _GEN_15163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15165 = 10'h4b == r_count_20_io_out ? io_r_75_b : _GEN_15164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15166 = 10'h4c == r_count_20_io_out ? io_r_76_b : _GEN_15165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15167 = 10'h4d == r_count_20_io_out ? io_r_77_b : _GEN_15166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15168 = 10'h4e == r_count_20_io_out ? io_r_78_b : _GEN_15167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15169 = 10'h4f == r_count_20_io_out ? io_r_79_b : _GEN_15168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15170 = 10'h50 == r_count_20_io_out ? io_r_80_b : _GEN_15169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15171 = 10'h51 == r_count_20_io_out ? io_r_81_b : _GEN_15170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15172 = 10'h52 == r_count_20_io_out ? io_r_82_b : _GEN_15171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15173 = 10'h53 == r_count_20_io_out ? io_r_83_b : _GEN_15172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15174 = 10'h54 == r_count_20_io_out ? io_r_84_b : _GEN_15173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15175 = 10'h55 == r_count_20_io_out ? io_r_85_b : _GEN_15174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15176 = 10'h56 == r_count_20_io_out ? io_r_86_b : _GEN_15175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15177 = 10'h57 == r_count_20_io_out ? io_r_87_b : _GEN_15176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15178 = 10'h58 == r_count_20_io_out ? io_r_88_b : _GEN_15177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15179 = 10'h59 == r_count_20_io_out ? io_r_89_b : _GEN_15178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15180 = 10'h5a == r_count_20_io_out ? io_r_90_b : _GEN_15179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15181 = 10'h5b == r_count_20_io_out ? io_r_91_b : _GEN_15180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15182 = 10'h5c == r_count_20_io_out ? io_r_92_b : _GEN_15181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15183 = 10'h5d == r_count_20_io_out ? io_r_93_b : _GEN_15182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15184 = 10'h5e == r_count_20_io_out ? io_r_94_b : _GEN_15183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15185 = 10'h5f == r_count_20_io_out ? io_r_95_b : _GEN_15184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15186 = 10'h60 == r_count_20_io_out ? io_r_96_b : _GEN_15185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15187 = 10'h61 == r_count_20_io_out ? io_r_97_b : _GEN_15186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15188 = 10'h62 == r_count_20_io_out ? io_r_98_b : _GEN_15187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15189 = 10'h63 == r_count_20_io_out ? io_r_99_b : _GEN_15188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15190 = 10'h64 == r_count_20_io_out ? io_r_100_b : _GEN_15189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15191 = 10'h65 == r_count_20_io_out ? io_r_101_b : _GEN_15190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15192 = 10'h66 == r_count_20_io_out ? io_r_102_b : _GEN_15191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15193 = 10'h67 == r_count_20_io_out ? io_r_103_b : _GEN_15192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15194 = 10'h68 == r_count_20_io_out ? io_r_104_b : _GEN_15193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15195 = 10'h69 == r_count_20_io_out ? io_r_105_b : _GEN_15194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15196 = 10'h6a == r_count_20_io_out ? io_r_106_b : _GEN_15195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15197 = 10'h6b == r_count_20_io_out ? io_r_107_b : _GEN_15196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15198 = 10'h6c == r_count_20_io_out ? io_r_108_b : _GEN_15197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15199 = 10'h6d == r_count_20_io_out ? io_r_109_b : _GEN_15198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15200 = 10'h6e == r_count_20_io_out ? io_r_110_b : _GEN_15199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15201 = 10'h6f == r_count_20_io_out ? io_r_111_b : _GEN_15200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15202 = 10'h70 == r_count_20_io_out ? io_r_112_b : _GEN_15201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15203 = 10'h71 == r_count_20_io_out ? io_r_113_b : _GEN_15202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15204 = 10'h72 == r_count_20_io_out ? io_r_114_b : _GEN_15203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15205 = 10'h73 == r_count_20_io_out ? io_r_115_b : _GEN_15204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15206 = 10'h74 == r_count_20_io_out ? io_r_116_b : _GEN_15205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15207 = 10'h75 == r_count_20_io_out ? io_r_117_b : _GEN_15206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15208 = 10'h76 == r_count_20_io_out ? io_r_118_b : _GEN_15207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15209 = 10'h77 == r_count_20_io_out ? io_r_119_b : _GEN_15208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15210 = 10'h78 == r_count_20_io_out ? io_r_120_b : _GEN_15209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15211 = 10'h79 == r_count_20_io_out ? io_r_121_b : _GEN_15210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15212 = 10'h7a == r_count_20_io_out ? io_r_122_b : _GEN_15211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15213 = 10'h7b == r_count_20_io_out ? io_r_123_b : _GEN_15212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15214 = 10'h7c == r_count_20_io_out ? io_r_124_b : _GEN_15213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15215 = 10'h7d == r_count_20_io_out ? io_r_125_b : _GEN_15214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15216 = 10'h7e == r_count_20_io_out ? io_r_126_b : _GEN_15215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15217 = 10'h7f == r_count_20_io_out ? io_r_127_b : _GEN_15216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15218 = 10'h80 == r_count_20_io_out ? io_r_128_b : _GEN_15217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15219 = 10'h81 == r_count_20_io_out ? io_r_129_b : _GEN_15218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15220 = 10'h82 == r_count_20_io_out ? io_r_130_b : _GEN_15219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15221 = 10'h83 == r_count_20_io_out ? io_r_131_b : _GEN_15220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15222 = 10'h84 == r_count_20_io_out ? io_r_132_b : _GEN_15221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15223 = 10'h85 == r_count_20_io_out ? io_r_133_b : _GEN_15222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15224 = 10'h86 == r_count_20_io_out ? io_r_134_b : _GEN_15223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15225 = 10'h87 == r_count_20_io_out ? io_r_135_b : _GEN_15224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15226 = 10'h88 == r_count_20_io_out ? io_r_136_b : _GEN_15225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15227 = 10'h89 == r_count_20_io_out ? io_r_137_b : _GEN_15226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15228 = 10'h8a == r_count_20_io_out ? io_r_138_b : _GEN_15227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15229 = 10'h8b == r_count_20_io_out ? io_r_139_b : _GEN_15228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15230 = 10'h8c == r_count_20_io_out ? io_r_140_b : _GEN_15229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15231 = 10'h8d == r_count_20_io_out ? io_r_141_b : _GEN_15230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15232 = 10'h8e == r_count_20_io_out ? io_r_142_b : _GEN_15231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15233 = 10'h8f == r_count_20_io_out ? io_r_143_b : _GEN_15232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15234 = 10'h90 == r_count_20_io_out ? io_r_144_b : _GEN_15233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15235 = 10'h91 == r_count_20_io_out ? io_r_145_b : _GEN_15234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15236 = 10'h92 == r_count_20_io_out ? io_r_146_b : _GEN_15235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15237 = 10'h93 == r_count_20_io_out ? io_r_147_b : _GEN_15236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15238 = 10'h94 == r_count_20_io_out ? io_r_148_b : _GEN_15237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15239 = 10'h95 == r_count_20_io_out ? io_r_149_b : _GEN_15238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15240 = 10'h96 == r_count_20_io_out ? io_r_150_b : _GEN_15239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15241 = 10'h97 == r_count_20_io_out ? io_r_151_b : _GEN_15240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15242 = 10'h98 == r_count_20_io_out ? io_r_152_b : _GEN_15241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15243 = 10'h99 == r_count_20_io_out ? io_r_153_b : _GEN_15242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15244 = 10'h9a == r_count_20_io_out ? io_r_154_b : _GEN_15243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15245 = 10'h9b == r_count_20_io_out ? io_r_155_b : _GEN_15244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15246 = 10'h9c == r_count_20_io_out ? io_r_156_b : _GEN_15245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15247 = 10'h9d == r_count_20_io_out ? io_r_157_b : _GEN_15246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15248 = 10'h9e == r_count_20_io_out ? io_r_158_b : _GEN_15247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15249 = 10'h9f == r_count_20_io_out ? io_r_159_b : _GEN_15248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15250 = 10'ha0 == r_count_20_io_out ? io_r_160_b : _GEN_15249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15251 = 10'ha1 == r_count_20_io_out ? io_r_161_b : _GEN_15250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15252 = 10'ha2 == r_count_20_io_out ? io_r_162_b : _GEN_15251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15253 = 10'ha3 == r_count_20_io_out ? io_r_163_b : _GEN_15252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15254 = 10'ha4 == r_count_20_io_out ? io_r_164_b : _GEN_15253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15255 = 10'ha5 == r_count_20_io_out ? io_r_165_b : _GEN_15254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15256 = 10'ha6 == r_count_20_io_out ? io_r_166_b : _GEN_15255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15257 = 10'ha7 == r_count_20_io_out ? io_r_167_b : _GEN_15256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15258 = 10'ha8 == r_count_20_io_out ? io_r_168_b : _GEN_15257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15259 = 10'ha9 == r_count_20_io_out ? io_r_169_b : _GEN_15258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15260 = 10'haa == r_count_20_io_out ? io_r_170_b : _GEN_15259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15261 = 10'hab == r_count_20_io_out ? io_r_171_b : _GEN_15260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15262 = 10'hac == r_count_20_io_out ? io_r_172_b : _GEN_15261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15263 = 10'had == r_count_20_io_out ? io_r_173_b : _GEN_15262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15264 = 10'hae == r_count_20_io_out ? io_r_174_b : _GEN_15263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15265 = 10'haf == r_count_20_io_out ? io_r_175_b : _GEN_15264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15266 = 10'hb0 == r_count_20_io_out ? io_r_176_b : _GEN_15265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15267 = 10'hb1 == r_count_20_io_out ? io_r_177_b : _GEN_15266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15268 = 10'hb2 == r_count_20_io_out ? io_r_178_b : _GEN_15267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15269 = 10'hb3 == r_count_20_io_out ? io_r_179_b : _GEN_15268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15270 = 10'hb4 == r_count_20_io_out ? io_r_180_b : _GEN_15269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15271 = 10'hb5 == r_count_20_io_out ? io_r_181_b : _GEN_15270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15272 = 10'hb6 == r_count_20_io_out ? io_r_182_b : _GEN_15271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15273 = 10'hb7 == r_count_20_io_out ? io_r_183_b : _GEN_15272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15274 = 10'hb8 == r_count_20_io_out ? io_r_184_b : _GEN_15273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15275 = 10'hb9 == r_count_20_io_out ? io_r_185_b : _GEN_15274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15276 = 10'hba == r_count_20_io_out ? io_r_186_b : _GEN_15275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15277 = 10'hbb == r_count_20_io_out ? io_r_187_b : _GEN_15276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15278 = 10'hbc == r_count_20_io_out ? io_r_188_b : _GEN_15277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15279 = 10'hbd == r_count_20_io_out ? io_r_189_b : _GEN_15278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15280 = 10'hbe == r_count_20_io_out ? io_r_190_b : _GEN_15279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15281 = 10'hbf == r_count_20_io_out ? io_r_191_b : _GEN_15280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15282 = 10'hc0 == r_count_20_io_out ? io_r_192_b : _GEN_15281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15283 = 10'hc1 == r_count_20_io_out ? io_r_193_b : _GEN_15282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15284 = 10'hc2 == r_count_20_io_out ? io_r_194_b : _GEN_15283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15285 = 10'hc3 == r_count_20_io_out ? io_r_195_b : _GEN_15284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15286 = 10'hc4 == r_count_20_io_out ? io_r_196_b : _GEN_15285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15287 = 10'hc5 == r_count_20_io_out ? io_r_197_b : _GEN_15286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15288 = 10'hc6 == r_count_20_io_out ? io_r_198_b : _GEN_15287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15289 = 10'hc7 == r_count_20_io_out ? io_r_199_b : _GEN_15288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15290 = 10'hc8 == r_count_20_io_out ? io_r_200_b : _GEN_15289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15291 = 10'hc9 == r_count_20_io_out ? io_r_201_b : _GEN_15290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15292 = 10'hca == r_count_20_io_out ? io_r_202_b : _GEN_15291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15293 = 10'hcb == r_count_20_io_out ? io_r_203_b : _GEN_15292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15294 = 10'hcc == r_count_20_io_out ? io_r_204_b : _GEN_15293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15295 = 10'hcd == r_count_20_io_out ? io_r_205_b : _GEN_15294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15296 = 10'hce == r_count_20_io_out ? io_r_206_b : _GEN_15295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15297 = 10'hcf == r_count_20_io_out ? io_r_207_b : _GEN_15296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15298 = 10'hd0 == r_count_20_io_out ? io_r_208_b : _GEN_15297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15299 = 10'hd1 == r_count_20_io_out ? io_r_209_b : _GEN_15298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15300 = 10'hd2 == r_count_20_io_out ? io_r_210_b : _GEN_15299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15301 = 10'hd3 == r_count_20_io_out ? io_r_211_b : _GEN_15300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15302 = 10'hd4 == r_count_20_io_out ? io_r_212_b : _GEN_15301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15303 = 10'hd5 == r_count_20_io_out ? io_r_213_b : _GEN_15302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15304 = 10'hd6 == r_count_20_io_out ? io_r_214_b : _GEN_15303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15305 = 10'hd7 == r_count_20_io_out ? io_r_215_b : _GEN_15304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15306 = 10'hd8 == r_count_20_io_out ? io_r_216_b : _GEN_15305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15307 = 10'hd9 == r_count_20_io_out ? io_r_217_b : _GEN_15306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15308 = 10'hda == r_count_20_io_out ? io_r_218_b : _GEN_15307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15309 = 10'hdb == r_count_20_io_out ? io_r_219_b : _GEN_15308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15310 = 10'hdc == r_count_20_io_out ? io_r_220_b : _GEN_15309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15311 = 10'hdd == r_count_20_io_out ? io_r_221_b : _GEN_15310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15312 = 10'hde == r_count_20_io_out ? io_r_222_b : _GEN_15311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15313 = 10'hdf == r_count_20_io_out ? io_r_223_b : _GEN_15312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15314 = 10'he0 == r_count_20_io_out ? io_r_224_b : _GEN_15313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15315 = 10'he1 == r_count_20_io_out ? io_r_225_b : _GEN_15314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15316 = 10'he2 == r_count_20_io_out ? io_r_226_b : _GEN_15315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15317 = 10'he3 == r_count_20_io_out ? io_r_227_b : _GEN_15316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15318 = 10'he4 == r_count_20_io_out ? io_r_228_b : _GEN_15317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15319 = 10'he5 == r_count_20_io_out ? io_r_229_b : _GEN_15318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15320 = 10'he6 == r_count_20_io_out ? io_r_230_b : _GEN_15319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15321 = 10'he7 == r_count_20_io_out ? io_r_231_b : _GEN_15320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15322 = 10'he8 == r_count_20_io_out ? io_r_232_b : _GEN_15321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15323 = 10'he9 == r_count_20_io_out ? io_r_233_b : _GEN_15322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15324 = 10'hea == r_count_20_io_out ? io_r_234_b : _GEN_15323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15325 = 10'heb == r_count_20_io_out ? io_r_235_b : _GEN_15324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15326 = 10'hec == r_count_20_io_out ? io_r_236_b : _GEN_15325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15327 = 10'hed == r_count_20_io_out ? io_r_237_b : _GEN_15326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15328 = 10'hee == r_count_20_io_out ? io_r_238_b : _GEN_15327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15329 = 10'hef == r_count_20_io_out ? io_r_239_b : _GEN_15328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15330 = 10'hf0 == r_count_20_io_out ? io_r_240_b : _GEN_15329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15331 = 10'hf1 == r_count_20_io_out ? io_r_241_b : _GEN_15330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15332 = 10'hf2 == r_count_20_io_out ? io_r_242_b : _GEN_15331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15333 = 10'hf3 == r_count_20_io_out ? io_r_243_b : _GEN_15332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15334 = 10'hf4 == r_count_20_io_out ? io_r_244_b : _GEN_15333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15335 = 10'hf5 == r_count_20_io_out ? io_r_245_b : _GEN_15334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15336 = 10'hf6 == r_count_20_io_out ? io_r_246_b : _GEN_15335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15337 = 10'hf7 == r_count_20_io_out ? io_r_247_b : _GEN_15336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15338 = 10'hf8 == r_count_20_io_out ? io_r_248_b : _GEN_15337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15339 = 10'hf9 == r_count_20_io_out ? io_r_249_b : _GEN_15338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15340 = 10'hfa == r_count_20_io_out ? io_r_250_b : _GEN_15339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15341 = 10'hfb == r_count_20_io_out ? io_r_251_b : _GEN_15340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15342 = 10'hfc == r_count_20_io_out ? io_r_252_b : _GEN_15341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15343 = 10'hfd == r_count_20_io_out ? io_r_253_b : _GEN_15342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15344 = 10'hfe == r_count_20_io_out ? io_r_254_b : _GEN_15343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15345 = 10'hff == r_count_20_io_out ? io_r_255_b : _GEN_15344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15346 = 10'h100 == r_count_20_io_out ? io_r_256_b : _GEN_15345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15347 = 10'h101 == r_count_20_io_out ? io_r_257_b : _GEN_15346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15348 = 10'h102 == r_count_20_io_out ? io_r_258_b : _GEN_15347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15349 = 10'h103 == r_count_20_io_out ? io_r_259_b : _GEN_15348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15350 = 10'h104 == r_count_20_io_out ? io_r_260_b : _GEN_15349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15351 = 10'h105 == r_count_20_io_out ? io_r_261_b : _GEN_15350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15352 = 10'h106 == r_count_20_io_out ? io_r_262_b : _GEN_15351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15353 = 10'h107 == r_count_20_io_out ? io_r_263_b : _GEN_15352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15354 = 10'h108 == r_count_20_io_out ? io_r_264_b : _GEN_15353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15355 = 10'h109 == r_count_20_io_out ? io_r_265_b : _GEN_15354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15356 = 10'h10a == r_count_20_io_out ? io_r_266_b : _GEN_15355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15357 = 10'h10b == r_count_20_io_out ? io_r_267_b : _GEN_15356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15358 = 10'h10c == r_count_20_io_out ? io_r_268_b : _GEN_15357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15359 = 10'h10d == r_count_20_io_out ? io_r_269_b : _GEN_15358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15360 = 10'h10e == r_count_20_io_out ? io_r_270_b : _GEN_15359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15361 = 10'h10f == r_count_20_io_out ? io_r_271_b : _GEN_15360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15362 = 10'h110 == r_count_20_io_out ? io_r_272_b : _GEN_15361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15363 = 10'h111 == r_count_20_io_out ? io_r_273_b : _GEN_15362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15364 = 10'h112 == r_count_20_io_out ? io_r_274_b : _GEN_15363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15365 = 10'h113 == r_count_20_io_out ? io_r_275_b : _GEN_15364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15366 = 10'h114 == r_count_20_io_out ? io_r_276_b : _GEN_15365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15367 = 10'h115 == r_count_20_io_out ? io_r_277_b : _GEN_15366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15368 = 10'h116 == r_count_20_io_out ? io_r_278_b : _GEN_15367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15369 = 10'h117 == r_count_20_io_out ? io_r_279_b : _GEN_15368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15370 = 10'h118 == r_count_20_io_out ? io_r_280_b : _GEN_15369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15371 = 10'h119 == r_count_20_io_out ? io_r_281_b : _GEN_15370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15372 = 10'h11a == r_count_20_io_out ? io_r_282_b : _GEN_15371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15373 = 10'h11b == r_count_20_io_out ? io_r_283_b : _GEN_15372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15374 = 10'h11c == r_count_20_io_out ? io_r_284_b : _GEN_15373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15375 = 10'h11d == r_count_20_io_out ? io_r_285_b : _GEN_15374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15376 = 10'h11e == r_count_20_io_out ? io_r_286_b : _GEN_15375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15377 = 10'h11f == r_count_20_io_out ? io_r_287_b : _GEN_15376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15378 = 10'h120 == r_count_20_io_out ? io_r_288_b : _GEN_15377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15379 = 10'h121 == r_count_20_io_out ? io_r_289_b : _GEN_15378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15380 = 10'h122 == r_count_20_io_out ? io_r_290_b : _GEN_15379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15381 = 10'h123 == r_count_20_io_out ? io_r_291_b : _GEN_15380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15382 = 10'h124 == r_count_20_io_out ? io_r_292_b : _GEN_15381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15383 = 10'h125 == r_count_20_io_out ? io_r_293_b : _GEN_15382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15384 = 10'h126 == r_count_20_io_out ? io_r_294_b : _GEN_15383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15385 = 10'h127 == r_count_20_io_out ? io_r_295_b : _GEN_15384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15386 = 10'h128 == r_count_20_io_out ? io_r_296_b : _GEN_15385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15387 = 10'h129 == r_count_20_io_out ? io_r_297_b : _GEN_15386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15388 = 10'h12a == r_count_20_io_out ? io_r_298_b : _GEN_15387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15389 = 10'h12b == r_count_20_io_out ? io_r_299_b : _GEN_15388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15390 = 10'h12c == r_count_20_io_out ? io_r_300_b : _GEN_15389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15391 = 10'h12d == r_count_20_io_out ? io_r_301_b : _GEN_15390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15392 = 10'h12e == r_count_20_io_out ? io_r_302_b : _GEN_15391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15393 = 10'h12f == r_count_20_io_out ? io_r_303_b : _GEN_15392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15394 = 10'h130 == r_count_20_io_out ? io_r_304_b : _GEN_15393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15395 = 10'h131 == r_count_20_io_out ? io_r_305_b : _GEN_15394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15396 = 10'h132 == r_count_20_io_out ? io_r_306_b : _GEN_15395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15397 = 10'h133 == r_count_20_io_out ? io_r_307_b : _GEN_15396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15398 = 10'h134 == r_count_20_io_out ? io_r_308_b : _GEN_15397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15399 = 10'h135 == r_count_20_io_out ? io_r_309_b : _GEN_15398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15400 = 10'h136 == r_count_20_io_out ? io_r_310_b : _GEN_15399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15401 = 10'h137 == r_count_20_io_out ? io_r_311_b : _GEN_15400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15402 = 10'h138 == r_count_20_io_out ? io_r_312_b : _GEN_15401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15403 = 10'h139 == r_count_20_io_out ? io_r_313_b : _GEN_15402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15404 = 10'h13a == r_count_20_io_out ? io_r_314_b : _GEN_15403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15405 = 10'h13b == r_count_20_io_out ? io_r_315_b : _GEN_15404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15406 = 10'h13c == r_count_20_io_out ? io_r_316_b : _GEN_15405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15407 = 10'h13d == r_count_20_io_out ? io_r_317_b : _GEN_15406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15408 = 10'h13e == r_count_20_io_out ? io_r_318_b : _GEN_15407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15409 = 10'h13f == r_count_20_io_out ? io_r_319_b : _GEN_15408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15410 = 10'h140 == r_count_20_io_out ? io_r_320_b : _GEN_15409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15411 = 10'h141 == r_count_20_io_out ? io_r_321_b : _GEN_15410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15412 = 10'h142 == r_count_20_io_out ? io_r_322_b : _GEN_15411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15413 = 10'h143 == r_count_20_io_out ? io_r_323_b : _GEN_15412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15414 = 10'h144 == r_count_20_io_out ? io_r_324_b : _GEN_15413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15415 = 10'h145 == r_count_20_io_out ? io_r_325_b : _GEN_15414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15416 = 10'h146 == r_count_20_io_out ? io_r_326_b : _GEN_15415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15417 = 10'h147 == r_count_20_io_out ? io_r_327_b : _GEN_15416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15418 = 10'h148 == r_count_20_io_out ? io_r_328_b : _GEN_15417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15419 = 10'h149 == r_count_20_io_out ? io_r_329_b : _GEN_15418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15420 = 10'h14a == r_count_20_io_out ? io_r_330_b : _GEN_15419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15421 = 10'h14b == r_count_20_io_out ? io_r_331_b : _GEN_15420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15422 = 10'h14c == r_count_20_io_out ? io_r_332_b : _GEN_15421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15423 = 10'h14d == r_count_20_io_out ? io_r_333_b : _GEN_15422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15424 = 10'h14e == r_count_20_io_out ? io_r_334_b : _GEN_15423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15425 = 10'h14f == r_count_20_io_out ? io_r_335_b : _GEN_15424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15426 = 10'h150 == r_count_20_io_out ? io_r_336_b : _GEN_15425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15427 = 10'h151 == r_count_20_io_out ? io_r_337_b : _GEN_15426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15428 = 10'h152 == r_count_20_io_out ? io_r_338_b : _GEN_15427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15429 = 10'h153 == r_count_20_io_out ? io_r_339_b : _GEN_15428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15430 = 10'h154 == r_count_20_io_out ? io_r_340_b : _GEN_15429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15431 = 10'h155 == r_count_20_io_out ? io_r_341_b : _GEN_15430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15432 = 10'h156 == r_count_20_io_out ? io_r_342_b : _GEN_15431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15433 = 10'h157 == r_count_20_io_out ? io_r_343_b : _GEN_15432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15434 = 10'h158 == r_count_20_io_out ? io_r_344_b : _GEN_15433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15435 = 10'h159 == r_count_20_io_out ? io_r_345_b : _GEN_15434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15436 = 10'h15a == r_count_20_io_out ? io_r_346_b : _GEN_15435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15437 = 10'h15b == r_count_20_io_out ? io_r_347_b : _GEN_15436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15438 = 10'h15c == r_count_20_io_out ? io_r_348_b : _GEN_15437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15439 = 10'h15d == r_count_20_io_out ? io_r_349_b : _GEN_15438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15440 = 10'h15e == r_count_20_io_out ? io_r_350_b : _GEN_15439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15441 = 10'h15f == r_count_20_io_out ? io_r_351_b : _GEN_15440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15442 = 10'h160 == r_count_20_io_out ? io_r_352_b : _GEN_15441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15443 = 10'h161 == r_count_20_io_out ? io_r_353_b : _GEN_15442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15444 = 10'h162 == r_count_20_io_out ? io_r_354_b : _GEN_15443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15445 = 10'h163 == r_count_20_io_out ? io_r_355_b : _GEN_15444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15446 = 10'h164 == r_count_20_io_out ? io_r_356_b : _GEN_15445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15447 = 10'h165 == r_count_20_io_out ? io_r_357_b : _GEN_15446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15448 = 10'h166 == r_count_20_io_out ? io_r_358_b : _GEN_15447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15449 = 10'h167 == r_count_20_io_out ? io_r_359_b : _GEN_15448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15450 = 10'h168 == r_count_20_io_out ? io_r_360_b : _GEN_15449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15451 = 10'h169 == r_count_20_io_out ? io_r_361_b : _GEN_15450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15452 = 10'h16a == r_count_20_io_out ? io_r_362_b : _GEN_15451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15453 = 10'h16b == r_count_20_io_out ? io_r_363_b : _GEN_15452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15454 = 10'h16c == r_count_20_io_out ? io_r_364_b : _GEN_15453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15455 = 10'h16d == r_count_20_io_out ? io_r_365_b : _GEN_15454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15456 = 10'h16e == r_count_20_io_out ? io_r_366_b : _GEN_15455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15457 = 10'h16f == r_count_20_io_out ? io_r_367_b : _GEN_15456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15458 = 10'h170 == r_count_20_io_out ? io_r_368_b : _GEN_15457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15459 = 10'h171 == r_count_20_io_out ? io_r_369_b : _GEN_15458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15460 = 10'h172 == r_count_20_io_out ? io_r_370_b : _GEN_15459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15461 = 10'h173 == r_count_20_io_out ? io_r_371_b : _GEN_15460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15462 = 10'h174 == r_count_20_io_out ? io_r_372_b : _GEN_15461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15463 = 10'h175 == r_count_20_io_out ? io_r_373_b : _GEN_15462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15464 = 10'h176 == r_count_20_io_out ? io_r_374_b : _GEN_15463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15465 = 10'h177 == r_count_20_io_out ? io_r_375_b : _GEN_15464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15466 = 10'h178 == r_count_20_io_out ? io_r_376_b : _GEN_15465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15467 = 10'h179 == r_count_20_io_out ? io_r_377_b : _GEN_15466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15468 = 10'h17a == r_count_20_io_out ? io_r_378_b : _GEN_15467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15469 = 10'h17b == r_count_20_io_out ? io_r_379_b : _GEN_15468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15470 = 10'h17c == r_count_20_io_out ? io_r_380_b : _GEN_15469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15471 = 10'h17d == r_count_20_io_out ? io_r_381_b : _GEN_15470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15472 = 10'h17e == r_count_20_io_out ? io_r_382_b : _GEN_15471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15473 = 10'h17f == r_count_20_io_out ? io_r_383_b : _GEN_15472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15474 = 10'h180 == r_count_20_io_out ? io_r_384_b : _GEN_15473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15475 = 10'h181 == r_count_20_io_out ? io_r_385_b : _GEN_15474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15476 = 10'h182 == r_count_20_io_out ? io_r_386_b : _GEN_15475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15477 = 10'h183 == r_count_20_io_out ? io_r_387_b : _GEN_15476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15478 = 10'h184 == r_count_20_io_out ? io_r_388_b : _GEN_15477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15479 = 10'h185 == r_count_20_io_out ? io_r_389_b : _GEN_15478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15480 = 10'h186 == r_count_20_io_out ? io_r_390_b : _GEN_15479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15481 = 10'h187 == r_count_20_io_out ? io_r_391_b : _GEN_15480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15482 = 10'h188 == r_count_20_io_out ? io_r_392_b : _GEN_15481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15483 = 10'h189 == r_count_20_io_out ? io_r_393_b : _GEN_15482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15484 = 10'h18a == r_count_20_io_out ? io_r_394_b : _GEN_15483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15485 = 10'h18b == r_count_20_io_out ? io_r_395_b : _GEN_15484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15486 = 10'h18c == r_count_20_io_out ? io_r_396_b : _GEN_15485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15487 = 10'h18d == r_count_20_io_out ? io_r_397_b : _GEN_15486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15488 = 10'h18e == r_count_20_io_out ? io_r_398_b : _GEN_15487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15489 = 10'h18f == r_count_20_io_out ? io_r_399_b : _GEN_15488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15490 = 10'h190 == r_count_20_io_out ? io_r_400_b : _GEN_15489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15491 = 10'h191 == r_count_20_io_out ? io_r_401_b : _GEN_15490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15492 = 10'h192 == r_count_20_io_out ? io_r_402_b : _GEN_15491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15493 = 10'h193 == r_count_20_io_out ? io_r_403_b : _GEN_15492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15494 = 10'h194 == r_count_20_io_out ? io_r_404_b : _GEN_15493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15495 = 10'h195 == r_count_20_io_out ? io_r_405_b : _GEN_15494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15496 = 10'h196 == r_count_20_io_out ? io_r_406_b : _GEN_15495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15497 = 10'h197 == r_count_20_io_out ? io_r_407_b : _GEN_15496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15498 = 10'h198 == r_count_20_io_out ? io_r_408_b : _GEN_15497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15499 = 10'h199 == r_count_20_io_out ? io_r_409_b : _GEN_15498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15500 = 10'h19a == r_count_20_io_out ? io_r_410_b : _GEN_15499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15501 = 10'h19b == r_count_20_io_out ? io_r_411_b : _GEN_15500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15502 = 10'h19c == r_count_20_io_out ? io_r_412_b : _GEN_15501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15503 = 10'h19d == r_count_20_io_out ? io_r_413_b : _GEN_15502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15504 = 10'h19e == r_count_20_io_out ? io_r_414_b : _GEN_15503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15505 = 10'h19f == r_count_20_io_out ? io_r_415_b : _GEN_15504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15506 = 10'h1a0 == r_count_20_io_out ? io_r_416_b : _GEN_15505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15507 = 10'h1a1 == r_count_20_io_out ? io_r_417_b : _GEN_15506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15508 = 10'h1a2 == r_count_20_io_out ? io_r_418_b : _GEN_15507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15509 = 10'h1a3 == r_count_20_io_out ? io_r_419_b : _GEN_15508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15510 = 10'h1a4 == r_count_20_io_out ? io_r_420_b : _GEN_15509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15511 = 10'h1a5 == r_count_20_io_out ? io_r_421_b : _GEN_15510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15512 = 10'h1a6 == r_count_20_io_out ? io_r_422_b : _GEN_15511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15513 = 10'h1a7 == r_count_20_io_out ? io_r_423_b : _GEN_15512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15514 = 10'h1a8 == r_count_20_io_out ? io_r_424_b : _GEN_15513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15515 = 10'h1a9 == r_count_20_io_out ? io_r_425_b : _GEN_15514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15516 = 10'h1aa == r_count_20_io_out ? io_r_426_b : _GEN_15515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15517 = 10'h1ab == r_count_20_io_out ? io_r_427_b : _GEN_15516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15518 = 10'h1ac == r_count_20_io_out ? io_r_428_b : _GEN_15517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15519 = 10'h1ad == r_count_20_io_out ? io_r_429_b : _GEN_15518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15520 = 10'h1ae == r_count_20_io_out ? io_r_430_b : _GEN_15519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15521 = 10'h1af == r_count_20_io_out ? io_r_431_b : _GEN_15520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15522 = 10'h1b0 == r_count_20_io_out ? io_r_432_b : _GEN_15521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15523 = 10'h1b1 == r_count_20_io_out ? io_r_433_b : _GEN_15522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15524 = 10'h1b2 == r_count_20_io_out ? io_r_434_b : _GEN_15523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15525 = 10'h1b3 == r_count_20_io_out ? io_r_435_b : _GEN_15524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15526 = 10'h1b4 == r_count_20_io_out ? io_r_436_b : _GEN_15525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15527 = 10'h1b5 == r_count_20_io_out ? io_r_437_b : _GEN_15526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15528 = 10'h1b6 == r_count_20_io_out ? io_r_438_b : _GEN_15527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15529 = 10'h1b7 == r_count_20_io_out ? io_r_439_b : _GEN_15528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15530 = 10'h1b8 == r_count_20_io_out ? io_r_440_b : _GEN_15529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15531 = 10'h1b9 == r_count_20_io_out ? io_r_441_b : _GEN_15530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15532 = 10'h1ba == r_count_20_io_out ? io_r_442_b : _GEN_15531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15533 = 10'h1bb == r_count_20_io_out ? io_r_443_b : _GEN_15532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15534 = 10'h1bc == r_count_20_io_out ? io_r_444_b : _GEN_15533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15535 = 10'h1bd == r_count_20_io_out ? io_r_445_b : _GEN_15534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15536 = 10'h1be == r_count_20_io_out ? io_r_446_b : _GEN_15535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15537 = 10'h1bf == r_count_20_io_out ? io_r_447_b : _GEN_15536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15538 = 10'h1c0 == r_count_20_io_out ? io_r_448_b : _GEN_15537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15539 = 10'h1c1 == r_count_20_io_out ? io_r_449_b : _GEN_15538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15540 = 10'h1c2 == r_count_20_io_out ? io_r_450_b : _GEN_15539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15541 = 10'h1c3 == r_count_20_io_out ? io_r_451_b : _GEN_15540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15542 = 10'h1c4 == r_count_20_io_out ? io_r_452_b : _GEN_15541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15543 = 10'h1c5 == r_count_20_io_out ? io_r_453_b : _GEN_15542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15544 = 10'h1c6 == r_count_20_io_out ? io_r_454_b : _GEN_15543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15545 = 10'h1c7 == r_count_20_io_out ? io_r_455_b : _GEN_15544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15546 = 10'h1c8 == r_count_20_io_out ? io_r_456_b : _GEN_15545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15547 = 10'h1c9 == r_count_20_io_out ? io_r_457_b : _GEN_15546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15548 = 10'h1ca == r_count_20_io_out ? io_r_458_b : _GEN_15547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15549 = 10'h1cb == r_count_20_io_out ? io_r_459_b : _GEN_15548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15550 = 10'h1cc == r_count_20_io_out ? io_r_460_b : _GEN_15549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15551 = 10'h1cd == r_count_20_io_out ? io_r_461_b : _GEN_15550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15552 = 10'h1ce == r_count_20_io_out ? io_r_462_b : _GEN_15551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15553 = 10'h1cf == r_count_20_io_out ? io_r_463_b : _GEN_15552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15554 = 10'h1d0 == r_count_20_io_out ? io_r_464_b : _GEN_15553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15555 = 10'h1d1 == r_count_20_io_out ? io_r_465_b : _GEN_15554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15556 = 10'h1d2 == r_count_20_io_out ? io_r_466_b : _GEN_15555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15557 = 10'h1d3 == r_count_20_io_out ? io_r_467_b : _GEN_15556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15558 = 10'h1d4 == r_count_20_io_out ? io_r_468_b : _GEN_15557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15559 = 10'h1d5 == r_count_20_io_out ? io_r_469_b : _GEN_15558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15560 = 10'h1d6 == r_count_20_io_out ? io_r_470_b : _GEN_15559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15561 = 10'h1d7 == r_count_20_io_out ? io_r_471_b : _GEN_15560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15562 = 10'h1d8 == r_count_20_io_out ? io_r_472_b : _GEN_15561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15563 = 10'h1d9 == r_count_20_io_out ? io_r_473_b : _GEN_15562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15564 = 10'h1da == r_count_20_io_out ? io_r_474_b : _GEN_15563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15565 = 10'h1db == r_count_20_io_out ? io_r_475_b : _GEN_15564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15566 = 10'h1dc == r_count_20_io_out ? io_r_476_b : _GEN_15565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15567 = 10'h1dd == r_count_20_io_out ? io_r_477_b : _GEN_15566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15568 = 10'h1de == r_count_20_io_out ? io_r_478_b : _GEN_15567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15569 = 10'h1df == r_count_20_io_out ? io_r_479_b : _GEN_15568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15570 = 10'h1e0 == r_count_20_io_out ? io_r_480_b : _GEN_15569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15571 = 10'h1e1 == r_count_20_io_out ? io_r_481_b : _GEN_15570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15572 = 10'h1e2 == r_count_20_io_out ? io_r_482_b : _GEN_15571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15573 = 10'h1e3 == r_count_20_io_out ? io_r_483_b : _GEN_15572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15574 = 10'h1e4 == r_count_20_io_out ? io_r_484_b : _GEN_15573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15575 = 10'h1e5 == r_count_20_io_out ? io_r_485_b : _GEN_15574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15576 = 10'h1e6 == r_count_20_io_out ? io_r_486_b : _GEN_15575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15577 = 10'h1e7 == r_count_20_io_out ? io_r_487_b : _GEN_15576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15578 = 10'h1e8 == r_count_20_io_out ? io_r_488_b : _GEN_15577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15579 = 10'h1e9 == r_count_20_io_out ? io_r_489_b : _GEN_15578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15580 = 10'h1ea == r_count_20_io_out ? io_r_490_b : _GEN_15579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15581 = 10'h1eb == r_count_20_io_out ? io_r_491_b : _GEN_15580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15582 = 10'h1ec == r_count_20_io_out ? io_r_492_b : _GEN_15581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15583 = 10'h1ed == r_count_20_io_out ? io_r_493_b : _GEN_15582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15584 = 10'h1ee == r_count_20_io_out ? io_r_494_b : _GEN_15583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15585 = 10'h1ef == r_count_20_io_out ? io_r_495_b : _GEN_15584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15586 = 10'h1f0 == r_count_20_io_out ? io_r_496_b : _GEN_15585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15587 = 10'h1f1 == r_count_20_io_out ? io_r_497_b : _GEN_15586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15588 = 10'h1f2 == r_count_20_io_out ? io_r_498_b : _GEN_15587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15589 = 10'h1f3 == r_count_20_io_out ? io_r_499_b : _GEN_15588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15590 = 10'h1f4 == r_count_20_io_out ? io_r_500_b : _GEN_15589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15591 = 10'h1f5 == r_count_20_io_out ? io_r_501_b : _GEN_15590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15592 = 10'h1f6 == r_count_20_io_out ? io_r_502_b : _GEN_15591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15593 = 10'h1f7 == r_count_20_io_out ? io_r_503_b : _GEN_15592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15594 = 10'h1f8 == r_count_20_io_out ? io_r_504_b : _GEN_15593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15595 = 10'h1f9 == r_count_20_io_out ? io_r_505_b : _GEN_15594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15596 = 10'h1fa == r_count_20_io_out ? io_r_506_b : _GEN_15595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15597 = 10'h1fb == r_count_20_io_out ? io_r_507_b : _GEN_15596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15598 = 10'h1fc == r_count_20_io_out ? io_r_508_b : _GEN_15597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15599 = 10'h1fd == r_count_20_io_out ? io_r_509_b : _GEN_15598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15600 = 10'h1fe == r_count_20_io_out ? io_r_510_b : _GEN_15599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15601 = 10'h1ff == r_count_20_io_out ? io_r_511_b : _GEN_15600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15602 = 10'h200 == r_count_20_io_out ? io_r_512_b : _GEN_15601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15603 = 10'h201 == r_count_20_io_out ? io_r_513_b : _GEN_15602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15604 = 10'h202 == r_count_20_io_out ? io_r_514_b : _GEN_15603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15605 = 10'h203 == r_count_20_io_out ? io_r_515_b : _GEN_15604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15606 = 10'h204 == r_count_20_io_out ? io_r_516_b : _GEN_15605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15607 = 10'h205 == r_count_20_io_out ? io_r_517_b : _GEN_15606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15608 = 10'h206 == r_count_20_io_out ? io_r_518_b : _GEN_15607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15609 = 10'h207 == r_count_20_io_out ? io_r_519_b : _GEN_15608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15610 = 10'h208 == r_count_20_io_out ? io_r_520_b : _GEN_15609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15611 = 10'h209 == r_count_20_io_out ? io_r_521_b : _GEN_15610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15612 = 10'h20a == r_count_20_io_out ? io_r_522_b : _GEN_15611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15613 = 10'h20b == r_count_20_io_out ? io_r_523_b : _GEN_15612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15614 = 10'h20c == r_count_20_io_out ? io_r_524_b : _GEN_15613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15615 = 10'h20d == r_count_20_io_out ? io_r_525_b : _GEN_15614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15616 = 10'h20e == r_count_20_io_out ? io_r_526_b : _GEN_15615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15617 = 10'h20f == r_count_20_io_out ? io_r_527_b : _GEN_15616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15618 = 10'h210 == r_count_20_io_out ? io_r_528_b : _GEN_15617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15619 = 10'h211 == r_count_20_io_out ? io_r_529_b : _GEN_15618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15620 = 10'h212 == r_count_20_io_out ? io_r_530_b : _GEN_15619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15621 = 10'h213 == r_count_20_io_out ? io_r_531_b : _GEN_15620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15622 = 10'h214 == r_count_20_io_out ? io_r_532_b : _GEN_15621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15623 = 10'h215 == r_count_20_io_out ? io_r_533_b : _GEN_15622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15624 = 10'h216 == r_count_20_io_out ? io_r_534_b : _GEN_15623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15625 = 10'h217 == r_count_20_io_out ? io_r_535_b : _GEN_15624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15626 = 10'h218 == r_count_20_io_out ? io_r_536_b : _GEN_15625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15627 = 10'h219 == r_count_20_io_out ? io_r_537_b : _GEN_15626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15628 = 10'h21a == r_count_20_io_out ? io_r_538_b : _GEN_15627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15629 = 10'h21b == r_count_20_io_out ? io_r_539_b : _GEN_15628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15630 = 10'h21c == r_count_20_io_out ? io_r_540_b : _GEN_15629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15631 = 10'h21d == r_count_20_io_out ? io_r_541_b : _GEN_15630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15632 = 10'h21e == r_count_20_io_out ? io_r_542_b : _GEN_15631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15633 = 10'h21f == r_count_20_io_out ? io_r_543_b : _GEN_15632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15634 = 10'h220 == r_count_20_io_out ? io_r_544_b : _GEN_15633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15635 = 10'h221 == r_count_20_io_out ? io_r_545_b : _GEN_15634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15636 = 10'h222 == r_count_20_io_out ? io_r_546_b : _GEN_15635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15637 = 10'h223 == r_count_20_io_out ? io_r_547_b : _GEN_15636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15638 = 10'h224 == r_count_20_io_out ? io_r_548_b : _GEN_15637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15639 = 10'h225 == r_count_20_io_out ? io_r_549_b : _GEN_15638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15640 = 10'h226 == r_count_20_io_out ? io_r_550_b : _GEN_15639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15641 = 10'h227 == r_count_20_io_out ? io_r_551_b : _GEN_15640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15642 = 10'h228 == r_count_20_io_out ? io_r_552_b : _GEN_15641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15643 = 10'h229 == r_count_20_io_out ? io_r_553_b : _GEN_15642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15644 = 10'h22a == r_count_20_io_out ? io_r_554_b : _GEN_15643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15645 = 10'h22b == r_count_20_io_out ? io_r_555_b : _GEN_15644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15646 = 10'h22c == r_count_20_io_out ? io_r_556_b : _GEN_15645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15647 = 10'h22d == r_count_20_io_out ? io_r_557_b : _GEN_15646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15648 = 10'h22e == r_count_20_io_out ? io_r_558_b : _GEN_15647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15649 = 10'h22f == r_count_20_io_out ? io_r_559_b : _GEN_15648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15650 = 10'h230 == r_count_20_io_out ? io_r_560_b : _GEN_15649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15651 = 10'h231 == r_count_20_io_out ? io_r_561_b : _GEN_15650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15652 = 10'h232 == r_count_20_io_out ? io_r_562_b : _GEN_15651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15653 = 10'h233 == r_count_20_io_out ? io_r_563_b : _GEN_15652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15654 = 10'h234 == r_count_20_io_out ? io_r_564_b : _GEN_15653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15655 = 10'h235 == r_count_20_io_out ? io_r_565_b : _GEN_15654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15656 = 10'h236 == r_count_20_io_out ? io_r_566_b : _GEN_15655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15657 = 10'h237 == r_count_20_io_out ? io_r_567_b : _GEN_15656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15658 = 10'h238 == r_count_20_io_out ? io_r_568_b : _GEN_15657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15659 = 10'h239 == r_count_20_io_out ? io_r_569_b : _GEN_15658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15660 = 10'h23a == r_count_20_io_out ? io_r_570_b : _GEN_15659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15661 = 10'h23b == r_count_20_io_out ? io_r_571_b : _GEN_15660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15662 = 10'h23c == r_count_20_io_out ? io_r_572_b : _GEN_15661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15663 = 10'h23d == r_count_20_io_out ? io_r_573_b : _GEN_15662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15664 = 10'h23e == r_count_20_io_out ? io_r_574_b : _GEN_15663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15665 = 10'h23f == r_count_20_io_out ? io_r_575_b : _GEN_15664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15666 = 10'h240 == r_count_20_io_out ? io_r_576_b : _GEN_15665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15667 = 10'h241 == r_count_20_io_out ? io_r_577_b : _GEN_15666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15668 = 10'h242 == r_count_20_io_out ? io_r_578_b : _GEN_15667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15669 = 10'h243 == r_count_20_io_out ? io_r_579_b : _GEN_15668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15670 = 10'h244 == r_count_20_io_out ? io_r_580_b : _GEN_15669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15671 = 10'h245 == r_count_20_io_out ? io_r_581_b : _GEN_15670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15672 = 10'h246 == r_count_20_io_out ? io_r_582_b : _GEN_15671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15673 = 10'h247 == r_count_20_io_out ? io_r_583_b : _GEN_15672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15674 = 10'h248 == r_count_20_io_out ? io_r_584_b : _GEN_15673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15675 = 10'h249 == r_count_20_io_out ? io_r_585_b : _GEN_15674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15676 = 10'h24a == r_count_20_io_out ? io_r_586_b : _GEN_15675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15677 = 10'h24b == r_count_20_io_out ? io_r_587_b : _GEN_15676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15678 = 10'h24c == r_count_20_io_out ? io_r_588_b : _GEN_15677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15679 = 10'h24d == r_count_20_io_out ? io_r_589_b : _GEN_15678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15680 = 10'h24e == r_count_20_io_out ? io_r_590_b : _GEN_15679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15681 = 10'h24f == r_count_20_io_out ? io_r_591_b : _GEN_15680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15682 = 10'h250 == r_count_20_io_out ? io_r_592_b : _GEN_15681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15683 = 10'h251 == r_count_20_io_out ? io_r_593_b : _GEN_15682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15684 = 10'h252 == r_count_20_io_out ? io_r_594_b : _GEN_15683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15685 = 10'h253 == r_count_20_io_out ? io_r_595_b : _GEN_15684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15686 = 10'h254 == r_count_20_io_out ? io_r_596_b : _GEN_15685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15687 = 10'h255 == r_count_20_io_out ? io_r_597_b : _GEN_15686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15688 = 10'h256 == r_count_20_io_out ? io_r_598_b : _GEN_15687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15689 = 10'h257 == r_count_20_io_out ? io_r_599_b : _GEN_15688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15690 = 10'h258 == r_count_20_io_out ? io_r_600_b : _GEN_15689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15691 = 10'h259 == r_count_20_io_out ? io_r_601_b : _GEN_15690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15692 = 10'h25a == r_count_20_io_out ? io_r_602_b : _GEN_15691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15693 = 10'h25b == r_count_20_io_out ? io_r_603_b : _GEN_15692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15694 = 10'h25c == r_count_20_io_out ? io_r_604_b : _GEN_15693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15695 = 10'h25d == r_count_20_io_out ? io_r_605_b : _GEN_15694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15696 = 10'h25e == r_count_20_io_out ? io_r_606_b : _GEN_15695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15697 = 10'h25f == r_count_20_io_out ? io_r_607_b : _GEN_15696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15698 = 10'h260 == r_count_20_io_out ? io_r_608_b : _GEN_15697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15699 = 10'h261 == r_count_20_io_out ? io_r_609_b : _GEN_15698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15700 = 10'h262 == r_count_20_io_out ? io_r_610_b : _GEN_15699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15701 = 10'h263 == r_count_20_io_out ? io_r_611_b : _GEN_15700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15702 = 10'h264 == r_count_20_io_out ? io_r_612_b : _GEN_15701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15703 = 10'h265 == r_count_20_io_out ? io_r_613_b : _GEN_15702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15704 = 10'h266 == r_count_20_io_out ? io_r_614_b : _GEN_15703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15705 = 10'h267 == r_count_20_io_out ? io_r_615_b : _GEN_15704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15706 = 10'h268 == r_count_20_io_out ? io_r_616_b : _GEN_15705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15707 = 10'h269 == r_count_20_io_out ? io_r_617_b : _GEN_15706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15708 = 10'h26a == r_count_20_io_out ? io_r_618_b : _GEN_15707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15709 = 10'h26b == r_count_20_io_out ? io_r_619_b : _GEN_15708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15710 = 10'h26c == r_count_20_io_out ? io_r_620_b : _GEN_15709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15711 = 10'h26d == r_count_20_io_out ? io_r_621_b : _GEN_15710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15712 = 10'h26e == r_count_20_io_out ? io_r_622_b : _GEN_15711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15713 = 10'h26f == r_count_20_io_out ? io_r_623_b : _GEN_15712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15714 = 10'h270 == r_count_20_io_out ? io_r_624_b : _GEN_15713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15715 = 10'h271 == r_count_20_io_out ? io_r_625_b : _GEN_15714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15716 = 10'h272 == r_count_20_io_out ? io_r_626_b : _GEN_15715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15717 = 10'h273 == r_count_20_io_out ? io_r_627_b : _GEN_15716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15718 = 10'h274 == r_count_20_io_out ? io_r_628_b : _GEN_15717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15719 = 10'h275 == r_count_20_io_out ? io_r_629_b : _GEN_15718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15720 = 10'h276 == r_count_20_io_out ? io_r_630_b : _GEN_15719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15721 = 10'h277 == r_count_20_io_out ? io_r_631_b : _GEN_15720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15722 = 10'h278 == r_count_20_io_out ? io_r_632_b : _GEN_15721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15723 = 10'h279 == r_count_20_io_out ? io_r_633_b : _GEN_15722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15724 = 10'h27a == r_count_20_io_out ? io_r_634_b : _GEN_15723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15725 = 10'h27b == r_count_20_io_out ? io_r_635_b : _GEN_15724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15726 = 10'h27c == r_count_20_io_out ? io_r_636_b : _GEN_15725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15727 = 10'h27d == r_count_20_io_out ? io_r_637_b : _GEN_15726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15728 = 10'h27e == r_count_20_io_out ? io_r_638_b : _GEN_15727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15729 = 10'h27f == r_count_20_io_out ? io_r_639_b : _GEN_15728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15730 = 10'h280 == r_count_20_io_out ? io_r_640_b : _GEN_15729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15731 = 10'h281 == r_count_20_io_out ? io_r_641_b : _GEN_15730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15732 = 10'h282 == r_count_20_io_out ? io_r_642_b : _GEN_15731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15733 = 10'h283 == r_count_20_io_out ? io_r_643_b : _GEN_15732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15734 = 10'h284 == r_count_20_io_out ? io_r_644_b : _GEN_15733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15735 = 10'h285 == r_count_20_io_out ? io_r_645_b : _GEN_15734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15736 = 10'h286 == r_count_20_io_out ? io_r_646_b : _GEN_15735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15737 = 10'h287 == r_count_20_io_out ? io_r_647_b : _GEN_15736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15738 = 10'h288 == r_count_20_io_out ? io_r_648_b : _GEN_15737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15739 = 10'h289 == r_count_20_io_out ? io_r_649_b : _GEN_15738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15740 = 10'h28a == r_count_20_io_out ? io_r_650_b : _GEN_15739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15741 = 10'h28b == r_count_20_io_out ? io_r_651_b : _GEN_15740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15742 = 10'h28c == r_count_20_io_out ? io_r_652_b : _GEN_15741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15743 = 10'h28d == r_count_20_io_out ? io_r_653_b : _GEN_15742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15744 = 10'h28e == r_count_20_io_out ? io_r_654_b : _GEN_15743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15745 = 10'h28f == r_count_20_io_out ? io_r_655_b : _GEN_15744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15746 = 10'h290 == r_count_20_io_out ? io_r_656_b : _GEN_15745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15747 = 10'h291 == r_count_20_io_out ? io_r_657_b : _GEN_15746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15748 = 10'h292 == r_count_20_io_out ? io_r_658_b : _GEN_15747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15749 = 10'h293 == r_count_20_io_out ? io_r_659_b : _GEN_15748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15750 = 10'h294 == r_count_20_io_out ? io_r_660_b : _GEN_15749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15751 = 10'h295 == r_count_20_io_out ? io_r_661_b : _GEN_15750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15752 = 10'h296 == r_count_20_io_out ? io_r_662_b : _GEN_15751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15753 = 10'h297 == r_count_20_io_out ? io_r_663_b : _GEN_15752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15754 = 10'h298 == r_count_20_io_out ? io_r_664_b : _GEN_15753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15755 = 10'h299 == r_count_20_io_out ? io_r_665_b : _GEN_15754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15756 = 10'h29a == r_count_20_io_out ? io_r_666_b : _GEN_15755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15757 = 10'h29b == r_count_20_io_out ? io_r_667_b : _GEN_15756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15758 = 10'h29c == r_count_20_io_out ? io_r_668_b : _GEN_15757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15759 = 10'h29d == r_count_20_io_out ? io_r_669_b : _GEN_15758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15760 = 10'h29e == r_count_20_io_out ? io_r_670_b : _GEN_15759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15761 = 10'h29f == r_count_20_io_out ? io_r_671_b : _GEN_15760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15762 = 10'h2a0 == r_count_20_io_out ? io_r_672_b : _GEN_15761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15763 = 10'h2a1 == r_count_20_io_out ? io_r_673_b : _GEN_15762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15764 = 10'h2a2 == r_count_20_io_out ? io_r_674_b : _GEN_15763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15765 = 10'h2a3 == r_count_20_io_out ? io_r_675_b : _GEN_15764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15766 = 10'h2a4 == r_count_20_io_out ? io_r_676_b : _GEN_15765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15767 = 10'h2a5 == r_count_20_io_out ? io_r_677_b : _GEN_15766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15768 = 10'h2a6 == r_count_20_io_out ? io_r_678_b : _GEN_15767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15769 = 10'h2a7 == r_count_20_io_out ? io_r_679_b : _GEN_15768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15770 = 10'h2a8 == r_count_20_io_out ? io_r_680_b : _GEN_15769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15771 = 10'h2a9 == r_count_20_io_out ? io_r_681_b : _GEN_15770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15772 = 10'h2aa == r_count_20_io_out ? io_r_682_b : _GEN_15771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15773 = 10'h2ab == r_count_20_io_out ? io_r_683_b : _GEN_15772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15774 = 10'h2ac == r_count_20_io_out ? io_r_684_b : _GEN_15773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15775 = 10'h2ad == r_count_20_io_out ? io_r_685_b : _GEN_15774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15776 = 10'h2ae == r_count_20_io_out ? io_r_686_b : _GEN_15775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15777 = 10'h2af == r_count_20_io_out ? io_r_687_b : _GEN_15776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15778 = 10'h2b0 == r_count_20_io_out ? io_r_688_b : _GEN_15777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15779 = 10'h2b1 == r_count_20_io_out ? io_r_689_b : _GEN_15778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15780 = 10'h2b2 == r_count_20_io_out ? io_r_690_b : _GEN_15779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15781 = 10'h2b3 == r_count_20_io_out ? io_r_691_b : _GEN_15780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15782 = 10'h2b4 == r_count_20_io_out ? io_r_692_b : _GEN_15781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15783 = 10'h2b5 == r_count_20_io_out ? io_r_693_b : _GEN_15782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15784 = 10'h2b6 == r_count_20_io_out ? io_r_694_b : _GEN_15783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15785 = 10'h2b7 == r_count_20_io_out ? io_r_695_b : _GEN_15784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15786 = 10'h2b8 == r_count_20_io_out ? io_r_696_b : _GEN_15785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15787 = 10'h2b9 == r_count_20_io_out ? io_r_697_b : _GEN_15786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15788 = 10'h2ba == r_count_20_io_out ? io_r_698_b : _GEN_15787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15789 = 10'h2bb == r_count_20_io_out ? io_r_699_b : _GEN_15788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15790 = 10'h2bc == r_count_20_io_out ? io_r_700_b : _GEN_15789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15791 = 10'h2bd == r_count_20_io_out ? io_r_701_b : _GEN_15790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15792 = 10'h2be == r_count_20_io_out ? io_r_702_b : _GEN_15791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15793 = 10'h2bf == r_count_20_io_out ? io_r_703_b : _GEN_15792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15794 = 10'h2c0 == r_count_20_io_out ? io_r_704_b : _GEN_15793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15795 = 10'h2c1 == r_count_20_io_out ? io_r_705_b : _GEN_15794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15796 = 10'h2c2 == r_count_20_io_out ? io_r_706_b : _GEN_15795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15797 = 10'h2c3 == r_count_20_io_out ? io_r_707_b : _GEN_15796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15798 = 10'h2c4 == r_count_20_io_out ? io_r_708_b : _GEN_15797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15799 = 10'h2c5 == r_count_20_io_out ? io_r_709_b : _GEN_15798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15800 = 10'h2c6 == r_count_20_io_out ? io_r_710_b : _GEN_15799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15801 = 10'h2c7 == r_count_20_io_out ? io_r_711_b : _GEN_15800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15802 = 10'h2c8 == r_count_20_io_out ? io_r_712_b : _GEN_15801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15803 = 10'h2c9 == r_count_20_io_out ? io_r_713_b : _GEN_15802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15804 = 10'h2ca == r_count_20_io_out ? io_r_714_b : _GEN_15803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15805 = 10'h2cb == r_count_20_io_out ? io_r_715_b : _GEN_15804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15806 = 10'h2cc == r_count_20_io_out ? io_r_716_b : _GEN_15805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15807 = 10'h2cd == r_count_20_io_out ? io_r_717_b : _GEN_15806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15808 = 10'h2ce == r_count_20_io_out ? io_r_718_b : _GEN_15807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15809 = 10'h2cf == r_count_20_io_out ? io_r_719_b : _GEN_15808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15810 = 10'h2d0 == r_count_20_io_out ? io_r_720_b : _GEN_15809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15811 = 10'h2d1 == r_count_20_io_out ? io_r_721_b : _GEN_15810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15812 = 10'h2d2 == r_count_20_io_out ? io_r_722_b : _GEN_15811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15813 = 10'h2d3 == r_count_20_io_out ? io_r_723_b : _GEN_15812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15814 = 10'h2d4 == r_count_20_io_out ? io_r_724_b : _GEN_15813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15815 = 10'h2d5 == r_count_20_io_out ? io_r_725_b : _GEN_15814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15816 = 10'h2d6 == r_count_20_io_out ? io_r_726_b : _GEN_15815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15817 = 10'h2d7 == r_count_20_io_out ? io_r_727_b : _GEN_15816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15818 = 10'h2d8 == r_count_20_io_out ? io_r_728_b : _GEN_15817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15819 = 10'h2d9 == r_count_20_io_out ? io_r_729_b : _GEN_15818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15820 = 10'h2da == r_count_20_io_out ? io_r_730_b : _GEN_15819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15821 = 10'h2db == r_count_20_io_out ? io_r_731_b : _GEN_15820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15822 = 10'h2dc == r_count_20_io_out ? io_r_732_b : _GEN_15821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15823 = 10'h2dd == r_count_20_io_out ? io_r_733_b : _GEN_15822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15824 = 10'h2de == r_count_20_io_out ? io_r_734_b : _GEN_15823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15825 = 10'h2df == r_count_20_io_out ? io_r_735_b : _GEN_15824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15826 = 10'h2e0 == r_count_20_io_out ? io_r_736_b : _GEN_15825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15827 = 10'h2e1 == r_count_20_io_out ? io_r_737_b : _GEN_15826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15828 = 10'h2e2 == r_count_20_io_out ? io_r_738_b : _GEN_15827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15829 = 10'h2e3 == r_count_20_io_out ? io_r_739_b : _GEN_15828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15830 = 10'h2e4 == r_count_20_io_out ? io_r_740_b : _GEN_15829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15831 = 10'h2e5 == r_count_20_io_out ? io_r_741_b : _GEN_15830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15832 = 10'h2e6 == r_count_20_io_out ? io_r_742_b : _GEN_15831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15833 = 10'h2e7 == r_count_20_io_out ? io_r_743_b : _GEN_15832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15834 = 10'h2e8 == r_count_20_io_out ? io_r_744_b : _GEN_15833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15835 = 10'h2e9 == r_count_20_io_out ? io_r_745_b : _GEN_15834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15836 = 10'h2ea == r_count_20_io_out ? io_r_746_b : _GEN_15835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15837 = 10'h2eb == r_count_20_io_out ? io_r_747_b : _GEN_15836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15838 = 10'h2ec == r_count_20_io_out ? io_r_748_b : _GEN_15837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15841 = 10'h1 == r_count_21_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15842 = 10'h2 == r_count_21_io_out ? io_r_2_b : _GEN_15841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15843 = 10'h3 == r_count_21_io_out ? io_r_3_b : _GEN_15842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15844 = 10'h4 == r_count_21_io_out ? io_r_4_b : _GEN_15843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15845 = 10'h5 == r_count_21_io_out ? io_r_5_b : _GEN_15844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15846 = 10'h6 == r_count_21_io_out ? io_r_6_b : _GEN_15845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15847 = 10'h7 == r_count_21_io_out ? io_r_7_b : _GEN_15846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15848 = 10'h8 == r_count_21_io_out ? io_r_8_b : _GEN_15847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15849 = 10'h9 == r_count_21_io_out ? io_r_9_b : _GEN_15848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15850 = 10'ha == r_count_21_io_out ? io_r_10_b : _GEN_15849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15851 = 10'hb == r_count_21_io_out ? io_r_11_b : _GEN_15850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15852 = 10'hc == r_count_21_io_out ? io_r_12_b : _GEN_15851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15853 = 10'hd == r_count_21_io_out ? io_r_13_b : _GEN_15852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15854 = 10'he == r_count_21_io_out ? io_r_14_b : _GEN_15853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15855 = 10'hf == r_count_21_io_out ? io_r_15_b : _GEN_15854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15856 = 10'h10 == r_count_21_io_out ? io_r_16_b : _GEN_15855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15857 = 10'h11 == r_count_21_io_out ? io_r_17_b : _GEN_15856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15858 = 10'h12 == r_count_21_io_out ? io_r_18_b : _GEN_15857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15859 = 10'h13 == r_count_21_io_out ? io_r_19_b : _GEN_15858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15860 = 10'h14 == r_count_21_io_out ? io_r_20_b : _GEN_15859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15861 = 10'h15 == r_count_21_io_out ? io_r_21_b : _GEN_15860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15862 = 10'h16 == r_count_21_io_out ? io_r_22_b : _GEN_15861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15863 = 10'h17 == r_count_21_io_out ? io_r_23_b : _GEN_15862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15864 = 10'h18 == r_count_21_io_out ? io_r_24_b : _GEN_15863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15865 = 10'h19 == r_count_21_io_out ? io_r_25_b : _GEN_15864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15866 = 10'h1a == r_count_21_io_out ? io_r_26_b : _GEN_15865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15867 = 10'h1b == r_count_21_io_out ? io_r_27_b : _GEN_15866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15868 = 10'h1c == r_count_21_io_out ? io_r_28_b : _GEN_15867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15869 = 10'h1d == r_count_21_io_out ? io_r_29_b : _GEN_15868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15870 = 10'h1e == r_count_21_io_out ? io_r_30_b : _GEN_15869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15871 = 10'h1f == r_count_21_io_out ? io_r_31_b : _GEN_15870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15872 = 10'h20 == r_count_21_io_out ? io_r_32_b : _GEN_15871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15873 = 10'h21 == r_count_21_io_out ? io_r_33_b : _GEN_15872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15874 = 10'h22 == r_count_21_io_out ? io_r_34_b : _GEN_15873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15875 = 10'h23 == r_count_21_io_out ? io_r_35_b : _GEN_15874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15876 = 10'h24 == r_count_21_io_out ? io_r_36_b : _GEN_15875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15877 = 10'h25 == r_count_21_io_out ? io_r_37_b : _GEN_15876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15878 = 10'h26 == r_count_21_io_out ? io_r_38_b : _GEN_15877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15879 = 10'h27 == r_count_21_io_out ? io_r_39_b : _GEN_15878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15880 = 10'h28 == r_count_21_io_out ? io_r_40_b : _GEN_15879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15881 = 10'h29 == r_count_21_io_out ? io_r_41_b : _GEN_15880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15882 = 10'h2a == r_count_21_io_out ? io_r_42_b : _GEN_15881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15883 = 10'h2b == r_count_21_io_out ? io_r_43_b : _GEN_15882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15884 = 10'h2c == r_count_21_io_out ? io_r_44_b : _GEN_15883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15885 = 10'h2d == r_count_21_io_out ? io_r_45_b : _GEN_15884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15886 = 10'h2e == r_count_21_io_out ? io_r_46_b : _GEN_15885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15887 = 10'h2f == r_count_21_io_out ? io_r_47_b : _GEN_15886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15888 = 10'h30 == r_count_21_io_out ? io_r_48_b : _GEN_15887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15889 = 10'h31 == r_count_21_io_out ? io_r_49_b : _GEN_15888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15890 = 10'h32 == r_count_21_io_out ? io_r_50_b : _GEN_15889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15891 = 10'h33 == r_count_21_io_out ? io_r_51_b : _GEN_15890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15892 = 10'h34 == r_count_21_io_out ? io_r_52_b : _GEN_15891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15893 = 10'h35 == r_count_21_io_out ? io_r_53_b : _GEN_15892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15894 = 10'h36 == r_count_21_io_out ? io_r_54_b : _GEN_15893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15895 = 10'h37 == r_count_21_io_out ? io_r_55_b : _GEN_15894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15896 = 10'h38 == r_count_21_io_out ? io_r_56_b : _GEN_15895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15897 = 10'h39 == r_count_21_io_out ? io_r_57_b : _GEN_15896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15898 = 10'h3a == r_count_21_io_out ? io_r_58_b : _GEN_15897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15899 = 10'h3b == r_count_21_io_out ? io_r_59_b : _GEN_15898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15900 = 10'h3c == r_count_21_io_out ? io_r_60_b : _GEN_15899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15901 = 10'h3d == r_count_21_io_out ? io_r_61_b : _GEN_15900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15902 = 10'h3e == r_count_21_io_out ? io_r_62_b : _GEN_15901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15903 = 10'h3f == r_count_21_io_out ? io_r_63_b : _GEN_15902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15904 = 10'h40 == r_count_21_io_out ? io_r_64_b : _GEN_15903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15905 = 10'h41 == r_count_21_io_out ? io_r_65_b : _GEN_15904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15906 = 10'h42 == r_count_21_io_out ? io_r_66_b : _GEN_15905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15907 = 10'h43 == r_count_21_io_out ? io_r_67_b : _GEN_15906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15908 = 10'h44 == r_count_21_io_out ? io_r_68_b : _GEN_15907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15909 = 10'h45 == r_count_21_io_out ? io_r_69_b : _GEN_15908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15910 = 10'h46 == r_count_21_io_out ? io_r_70_b : _GEN_15909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15911 = 10'h47 == r_count_21_io_out ? io_r_71_b : _GEN_15910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15912 = 10'h48 == r_count_21_io_out ? io_r_72_b : _GEN_15911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15913 = 10'h49 == r_count_21_io_out ? io_r_73_b : _GEN_15912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15914 = 10'h4a == r_count_21_io_out ? io_r_74_b : _GEN_15913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15915 = 10'h4b == r_count_21_io_out ? io_r_75_b : _GEN_15914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15916 = 10'h4c == r_count_21_io_out ? io_r_76_b : _GEN_15915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15917 = 10'h4d == r_count_21_io_out ? io_r_77_b : _GEN_15916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15918 = 10'h4e == r_count_21_io_out ? io_r_78_b : _GEN_15917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15919 = 10'h4f == r_count_21_io_out ? io_r_79_b : _GEN_15918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15920 = 10'h50 == r_count_21_io_out ? io_r_80_b : _GEN_15919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15921 = 10'h51 == r_count_21_io_out ? io_r_81_b : _GEN_15920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15922 = 10'h52 == r_count_21_io_out ? io_r_82_b : _GEN_15921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15923 = 10'h53 == r_count_21_io_out ? io_r_83_b : _GEN_15922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15924 = 10'h54 == r_count_21_io_out ? io_r_84_b : _GEN_15923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15925 = 10'h55 == r_count_21_io_out ? io_r_85_b : _GEN_15924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15926 = 10'h56 == r_count_21_io_out ? io_r_86_b : _GEN_15925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15927 = 10'h57 == r_count_21_io_out ? io_r_87_b : _GEN_15926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15928 = 10'h58 == r_count_21_io_out ? io_r_88_b : _GEN_15927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15929 = 10'h59 == r_count_21_io_out ? io_r_89_b : _GEN_15928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15930 = 10'h5a == r_count_21_io_out ? io_r_90_b : _GEN_15929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15931 = 10'h5b == r_count_21_io_out ? io_r_91_b : _GEN_15930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15932 = 10'h5c == r_count_21_io_out ? io_r_92_b : _GEN_15931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15933 = 10'h5d == r_count_21_io_out ? io_r_93_b : _GEN_15932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15934 = 10'h5e == r_count_21_io_out ? io_r_94_b : _GEN_15933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15935 = 10'h5f == r_count_21_io_out ? io_r_95_b : _GEN_15934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15936 = 10'h60 == r_count_21_io_out ? io_r_96_b : _GEN_15935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15937 = 10'h61 == r_count_21_io_out ? io_r_97_b : _GEN_15936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15938 = 10'h62 == r_count_21_io_out ? io_r_98_b : _GEN_15937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15939 = 10'h63 == r_count_21_io_out ? io_r_99_b : _GEN_15938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15940 = 10'h64 == r_count_21_io_out ? io_r_100_b : _GEN_15939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15941 = 10'h65 == r_count_21_io_out ? io_r_101_b : _GEN_15940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15942 = 10'h66 == r_count_21_io_out ? io_r_102_b : _GEN_15941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15943 = 10'h67 == r_count_21_io_out ? io_r_103_b : _GEN_15942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15944 = 10'h68 == r_count_21_io_out ? io_r_104_b : _GEN_15943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15945 = 10'h69 == r_count_21_io_out ? io_r_105_b : _GEN_15944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15946 = 10'h6a == r_count_21_io_out ? io_r_106_b : _GEN_15945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15947 = 10'h6b == r_count_21_io_out ? io_r_107_b : _GEN_15946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15948 = 10'h6c == r_count_21_io_out ? io_r_108_b : _GEN_15947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15949 = 10'h6d == r_count_21_io_out ? io_r_109_b : _GEN_15948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15950 = 10'h6e == r_count_21_io_out ? io_r_110_b : _GEN_15949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15951 = 10'h6f == r_count_21_io_out ? io_r_111_b : _GEN_15950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15952 = 10'h70 == r_count_21_io_out ? io_r_112_b : _GEN_15951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15953 = 10'h71 == r_count_21_io_out ? io_r_113_b : _GEN_15952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15954 = 10'h72 == r_count_21_io_out ? io_r_114_b : _GEN_15953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15955 = 10'h73 == r_count_21_io_out ? io_r_115_b : _GEN_15954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15956 = 10'h74 == r_count_21_io_out ? io_r_116_b : _GEN_15955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15957 = 10'h75 == r_count_21_io_out ? io_r_117_b : _GEN_15956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15958 = 10'h76 == r_count_21_io_out ? io_r_118_b : _GEN_15957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15959 = 10'h77 == r_count_21_io_out ? io_r_119_b : _GEN_15958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15960 = 10'h78 == r_count_21_io_out ? io_r_120_b : _GEN_15959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15961 = 10'h79 == r_count_21_io_out ? io_r_121_b : _GEN_15960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15962 = 10'h7a == r_count_21_io_out ? io_r_122_b : _GEN_15961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15963 = 10'h7b == r_count_21_io_out ? io_r_123_b : _GEN_15962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15964 = 10'h7c == r_count_21_io_out ? io_r_124_b : _GEN_15963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15965 = 10'h7d == r_count_21_io_out ? io_r_125_b : _GEN_15964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15966 = 10'h7e == r_count_21_io_out ? io_r_126_b : _GEN_15965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15967 = 10'h7f == r_count_21_io_out ? io_r_127_b : _GEN_15966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15968 = 10'h80 == r_count_21_io_out ? io_r_128_b : _GEN_15967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15969 = 10'h81 == r_count_21_io_out ? io_r_129_b : _GEN_15968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15970 = 10'h82 == r_count_21_io_out ? io_r_130_b : _GEN_15969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15971 = 10'h83 == r_count_21_io_out ? io_r_131_b : _GEN_15970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15972 = 10'h84 == r_count_21_io_out ? io_r_132_b : _GEN_15971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15973 = 10'h85 == r_count_21_io_out ? io_r_133_b : _GEN_15972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15974 = 10'h86 == r_count_21_io_out ? io_r_134_b : _GEN_15973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15975 = 10'h87 == r_count_21_io_out ? io_r_135_b : _GEN_15974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15976 = 10'h88 == r_count_21_io_out ? io_r_136_b : _GEN_15975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15977 = 10'h89 == r_count_21_io_out ? io_r_137_b : _GEN_15976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15978 = 10'h8a == r_count_21_io_out ? io_r_138_b : _GEN_15977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15979 = 10'h8b == r_count_21_io_out ? io_r_139_b : _GEN_15978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15980 = 10'h8c == r_count_21_io_out ? io_r_140_b : _GEN_15979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15981 = 10'h8d == r_count_21_io_out ? io_r_141_b : _GEN_15980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15982 = 10'h8e == r_count_21_io_out ? io_r_142_b : _GEN_15981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15983 = 10'h8f == r_count_21_io_out ? io_r_143_b : _GEN_15982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15984 = 10'h90 == r_count_21_io_out ? io_r_144_b : _GEN_15983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15985 = 10'h91 == r_count_21_io_out ? io_r_145_b : _GEN_15984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15986 = 10'h92 == r_count_21_io_out ? io_r_146_b : _GEN_15985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15987 = 10'h93 == r_count_21_io_out ? io_r_147_b : _GEN_15986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15988 = 10'h94 == r_count_21_io_out ? io_r_148_b : _GEN_15987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15989 = 10'h95 == r_count_21_io_out ? io_r_149_b : _GEN_15988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15990 = 10'h96 == r_count_21_io_out ? io_r_150_b : _GEN_15989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15991 = 10'h97 == r_count_21_io_out ? io_r_151_b : _GEN_15990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15992 = 10'h98 == r_count_21_io_out ? io_r_152_b : _GEN_15991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15993 = 10'h99 == r_count_21_io_out ? io_r_153_b : _GEN_15992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15994 = 10'h9a == r_count_21_io_out ? io_r_154_b : _GEN_15993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15995 = 10'h9b == r_count_21_io_out ? io_r_155_b : _GEN_15994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15996 = 10'h9c == r_count_21_io_out ? io_r_156_b : _GEN_15995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15997 = 10'h9d == r_count_21_io_out ? io_r_157_b : _GEN_15996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15998 = 10'h9e == r_count_21_io_out ? io_r_158_b : _GEN_15997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15999 = 10'h9f == r_count_21_io_out ? io_r_159_b : _GEN_15998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16000 = 10'ha0 == r_count_21_io_out ? io_r_160_b : _GEN_15999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16001 = 10'ha1 == r_count_21_io_out ? io_r_161_b : _GEN_16000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16002 = 10'ha2 == r_count_21_io_out ? io_r_162_b : _GEN_16001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16003 = 10'ha3 == r_count_21_io_out ? io_r_163_b : _GEN_16002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16004 = 10'ha4 == r_count_21_io_out ? io_r_164_b : _GEN_16003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16005 = 10'ha5 == r_count_21_io_out ? io_r_165_b : _GEN_16004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16006 = 10'ha6 == r_count_21_io_out ? io_r_166_b : _GEN_16005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16007 = 10'ha7 == r_count_21_io_out ? io_r_167_b : _GEN_16006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16008 = 10'ha8 == r_count_21_io_out ? io_r_168_b : _GEN_16007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16009 = 10'ha9 == r_count_21_io_out ? io_r_169_b : _GEN_16008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16010 = 10'haa == r_count_21_io_out ? io_r_170_b : _GEN_16009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16011 = 10'hab == r_count_21_io_out ? io_r_171_b : _GEN_16010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16012 = 10'hac == r_count_21_io_out ? io_r_172_b : _GEN_16011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16013 = 10'had == r_count_21_io_out ? io_r_173_b : _GEN_16012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16014 = 10'hae == r_count_21_io_out ? io_r_174_b : _GEN_16013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16015 = 10'haf == r_count_21_io_out ? io_r_175_b : _GEN_16014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16016 = 10'hb0 == r_count_21_io_out ? io_r_176_b : _GEN_16015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16017 = 10'hb1 == r_count_21_io_out ? io_r_177_b : _GEN_16016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16018 = 10'hb2 == r_count_21_io_out ? io_r_178_b : _GEN_16017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16019 = 10'hb3 == r_count_21_io_out ? io_r_179_b : _GEN_16018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16020 = 10'hb4 == r_count_21_io_out ? io_r_180_b : _GEN_16019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16021 = 10'hb5 == r_count_21_io_out ? io_r_181_b : _GEN_16020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16022 = 10'hb6 == r_count_21_io_out ? io_r_182_b : _GEN_16021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16023 = 10'hb7 == r_count_21_io_out ? io_r_183_b : _GEN_16022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16024 = 10'hb8 == r_count_21_io_out ? io_r_184_b : _GEN_16023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16025 = 10'hb9 == r_count_21_io_out ? io_r_185_b : _GEN_16024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16026 = 10'hba == r_count_21_io_out ? io_r_186_b : _GEN_16025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16027 = 10'hbb == r_count_21_io_out ? io_r_187_b : _GEN_16026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16028 = 10'hbc == r_count_21_io_out ? io_r_188_b : _GEN_16027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16029 = 10'hbd == r_count_21_io_out ? io_r_189_b : _GEN_16028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16030 = 10'hbe == r_count_21_io_out ? io_r_190_b : _GEN_16029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16031 = 10'hbf == r_count_21_io_out ? io_r_191_b : _GEN_16030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16032 = 10'hc0 == r_count_21_io_out ? io_r_192_b : _GEN_16031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16033 = 10'hc1 == r_count_21_io_out ? io_r_193_b : _GEN_16032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16034 = 10'hc2 == r_count_21_io_out ? io_r_194_b : _GEN_16033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16035 = 10'hc3 == r_count_21_io_out ? io_r_195_b : _GEN_16034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16036 = 10'hc4 == r_count_21_io_out ? io_r_196_b : _GEN_16035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16037 = 10'hc5 == r_count_21_io_out ? io_r_197_b : _GEN_16036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16038 = 10'hc6 == r_count_21_io_out ? io_r_198_b : _GEN_16037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16039 = 10'hc7 == r_count_21_io_out ? io_r_199_b : _GEN_16038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16040 = 10'hc8 == r_count_21_io_out ? io_r_200_b : _GEN_16039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16041 = 10'hc9 == r_count_21_io_out ? io_r_201_b : _GEN_16040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16042 = 10'hca == r_count_21_io_out ? io_r_202_b : _GEN_16041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16043 = 10'hcb == r_count_21_io_out ? io_r_203_b : _GEN_16042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16044 = 10'hcc == r_count_21_io_out ? io_r_204_b : _GEN_16043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16045 = 10'hcd == r_count_21_io_out ? io_r_205_b : _GEN_16044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16046 = 10'hce == r_count_21_io_out ? io_r_206_b : _GEN_16045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16047 = 10'hcf == r_count_21_io_out ? io_r_207_b : _GEN_16046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16048 = 10'hd0 == r_count_21_io_out ? io_r_208_b : _GEN_16047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16049 = 10'hd1 == r_count_21_io_out ? io_r_209_b : _GEN_16048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16050 = 10'hd2 == r_count_21_io_out ? io_r_210_b : _GEN_16049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16051 = 10'hd3 == r_count_21_io_out ? io_r_211_b : _GEN_16050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16052 = 10'hd4 == r_count_21_io_out ? io_r_212_b : _GEN_16051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16053 = 10'hd5 == r_count_21_io_out ? io_r_213_b : _GEN_16052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16054 = 10'hd6 == r_count_21_io_out ? io_r_214_b : _GEN_16053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16055 = 10'hd7 == r_count_21_io_out ? io_r_215_b : _GEN_16054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16056 = 10'hd8 == r_count_21_io_out ? io_r_216_b : _GEN_16055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16057 = 10'hd9 == r_count_21_io_out ? io_r_217_b : _GEN_16056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16058 = 10'hda == r_count_21_io_out ? io_r_218_b : _GEN_16057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16059 = 10'hdb == r_count_21_io_out ? io_r_219_b : _GEN_16058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16060 = 10'hdc == r_count_21_io_out ? io_r_220_b : _GEN_16059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16061 = 10'hdd == r_count_21_io_out ? io_r_221_b : _GEN_16060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16062 = 10'hde == r_count_21_io_out ? io_r_222_b : _GEN_16061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16063 = 10'hdf == r_count_21_io_out ? io_r_223_b : _GEN_16062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16064 = 10'he0 == r_count_21_io_out ? io_r_224_b : _GEN_16063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16065 = 10'he1 == r_count_21_io_out ? io_r_225_b : _GEN_16064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16066 = 10'he2 == r_count_21_io_out ? io_r_226_b : _GEN_16065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16067 = 10'he3 == r_count_21_io_out ? io_r_227_b : _GEN_16066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16068 = 10'he4 == r_count_21_io_out ? io_r_228_b : _GEN_16067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16069 = 10'he5 == r_count_21_io_out ? io_r_229_b : _GEN_16068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16070 = 10'he6 == r_count_21_io_out ? io_r_230_b : _GEN_16069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16071 = 10'he7 == r_count_21_io_out ? io_r_231_b : _GEN_16070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16072 = 10'he8 == r_count_21_io_out ? io_r_232_b : _GEN_16071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16073 = 10'he9 == r_count_21_io_out ? io_r_233_b : _GEN_16072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16074 = 10'hea == r_count_21_io_out ? io_r_234_b : _GEN_16073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16075 = 10'heb == r_count_21_io_out ? io_r_235_b : _GEN_16074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16076 = 10'hec == r_count_21_io_out ? io_r_236_b : _GEN_16075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16077 = 10'hed == r_count_21_io_out ? io_r_237_b : _GEN_16076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16078 = 10'hee == r_count_21_io_out ? io_r_238_b : _GEN_16077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16079 = 10'hef == r_count_21_io_out ? io_r_239_b : _GEN_16078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16080 = 10'hf0 == r_count_21_io_out ? io_r_240_b : _GEN_16079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16081 = 10'hf1 == r_count_21_io_out ? io_r_241_b : _GEN_16080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16082 = 10'hf2 == r_count_21_io_out ? io_r_242_b : _GEN_16081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16083 = 10'hf3 == r_count_21_io_out ? io_r_243_b : _GEN_16082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16084 = 10'hf4 == r_count_21_io_out ? io_r_244_b : _GEN_16083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16085 = 10'hf5 == r_count_21_io_out ? io_r_245_b : _GEN_16084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16086 = 10'hf6 == r_count_21_io_out ? io_r_246_b : _GEN_16085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16087 = 10'hf7 == r_count_21_io_out ? io_r_247_b : _GEN_16086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16088 = 10'hf8 == r_count_21_io_out ? io_r_248_b : _GEN_16087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16089 = 10'hf9 == r_count_21_io_out ? io_r_249_b : _GEN_16088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16090 = 10'hfa == r_count_21_io_out ? io_r_250_b : _GEN_16089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16091 = 10'hfb == r_count_21_io_out ? io_r_251_b : _GEN_16090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16092 = 10'hfc == r_count_21_io_out ? io_r_252_b : _GEN_16091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16093 = 10'hfd == r_count_21_io_out ? io_r_253_b : _GEN_16092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16094 = 10'hfe == r_count_21_io_out ? io_r_254_b : _GEN_16093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16095 = 10'hff == r_count_21_io_out ? io_r_255_b : _GEN_16094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16096 = 10'h100 == r_count_21_io_out ? io_r_256_b : _GEN_16095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16097 = 10'h101 == r_count_21_io_out ? io_r_257_b : _GEN_16096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16098 = 10'h102 == r_count_21_io_out ? io_r_258_b : _GEN_16097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16099 = 10'h103 == r_count_21_io_out ? io_r_259_b : _GEN_16098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16100 = 10'h104 == r_count_21_io_out ? io_r_260_b : _GEN_16099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16101 = 10'h105 == r_count_21_io_out ? io_r_261_b : _GEN_16100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16102 = 10'h106 == r_count_21_io_out ? io_r_262_b : _GEN_16101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16103 = 10'h107 == r_count_21_io_out ? io_r_263_b : _GEN_16102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16104 = 10'h108 == r_count_21_io_out ? io_r_264_b : _GEN_16103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16105 = 10'h109 == r_count_21_io_out ? io_r_265_b : _GEN_16104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16106 = 10'h10a == r_count_21_io_out ? io_r_266_b : _GEN_16105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16107 = 10'h10b == r_count_21_io_out ? io_r_267_b : _GEN_16106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16108 = 10'h10c == r_count_21_io_out ? io_r_268_b : _GEN_16107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16109 = 10'h10d == r_count_21_io_out ? io_r_269_b : _GEN_16108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16110 = 10'h10e == r_count_21_io_out ? io_r_270_b : _GEN_16109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16111 = 10'h10f == r_count_21_io_out ? io_r_271_b : _GEN_16110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16112 = 10'h110 == r_count_21_io_out ? io_r_272_b : _GEN_16111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16113 = 10'h111 == r_count_21_io_out ? io_r_273_b : _GEN_16112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16114 = 10'h112 == r_count_21_io_out ? io_r_274_b : _GEN_16113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16115 = 10'h113 == r_count_21_io_out ? io_r_275_b : _GEN_16114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16116 = 10'h114 == r_count_21_io_out ? io_r_276_b : _GEN_16115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16117 = 10'h115 == r_count_21_io_out ? io_r_277_b : _GEN_16116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16118 = 10'h116 == r_count_21_io_out ? io_r_278_b : _GEN_16117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16119 = 10'h117 == r_count_21_io_out ? io_r_279_b : _GEN_16118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16120 = 10'h118 == r_count_21_io_out ? io_r_280_b : _GEN_16119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16121 = 10'h119 == r_count_21_io_out ? io_r_281_b : _GEN_16120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16122 = 10'h11a == r_count_21_io_out ? io_r_282_b : _GEN_16121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16123 = 10'h11b == r_count_21_io_out ? io_r_283_b : _GEN_16122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16124 = 10'h11c == r_count_21_io_out ? io_r_284_b : _GEN_16123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16125 = 10'h11d == r_count_21_io_out ? io_r_285_b : _GEN_16124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16126 = 10'h11e == r_count_21_io_out ? io_r_286_b : _GEN_16125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16127 = 10'h11f == r_count_21_io_out ? io_r_287_b : _GEN_16126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16128 = 10'h120 == r_count_21_io_out ? io_r_288_b : _GEN_16127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16129 = 10'h121 == r_count_21_io_out ? io_r_289_b : _GEN_16128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16130 = 10'h122 == r_count_21_io_out ? io_r_290_b : _GEN_16129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16131 = 10'h123 == r_count_21_io_out ? io_r_291_b : _GEN_16130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16132 = 10'h124 == r_count_21_io_out ? io_r_292_b : _GEN_16131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16133 = 10'h125 == r_count_21_io_out ? io_r_293_b : _GEN_16132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16134 = 10'h126 == r_count_21_io_out ? io_r_294_b : _GEN_16133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16135 = 10'h127 == r_count_21_io_out ? io_r_295_b : _GEN_16134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16136 = 10'h128 == r_count_21_io_out ? io_r_296_b : _GEN_16135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16137 = 10'h129 == r_count_21_io_out ? io_r_297_b : _GEN_16136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16138 = 10'h12a == r_count_21_io_out ? io_r_298_b : _GEN_16137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16139 = 10'h12b == r_count_21_io_out ? io_r_299_b : _GEN_16138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16140 = 10'h12c == r_count_21_io_out ? io_r_300_b : _GEN_16139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16141 = 10'h12d == r_count_21_io_out ? io_r_301_b : _GEN_16140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16142 = 10'h12e == r_count_21_io_out ? io_r_302_b : _GEN_16141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16143 = 10'h12f == r_count_21_io_out ? io_r_303_b : _GEN_16142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16144 = 10'h130 == r_count_21_io_out ? io_r_304_b : _GEN_16143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16145 = 10'h131 == r_count_21_io_out ? io_r_305_b : _GEN_16144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16146 = 10'h132 == r_count_21_io_out ? io_r_306_b : _GEN_16145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16147 = 10'h133 == r_count_21_io_out ? io_r_307_b : _GEN_16146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16148 = 10'h134 == r_count_21_io_out ? io_r_308_b : _GEN_16147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16149 = 10'h135 == r_count_21_io_out ? io_r_309_b : _GEN_16148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16150 = 10'h136 == r_count_21_io_out ? io_r_310_b : _GEN_16149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16151 = 10'h137 == r_count_21_io_out ? io_r_311_b : _GEN_16150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16152 = 10'h138 == r_count_21_io_out ? io_r_312_b : _GEN_16151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16153 = 10'h139 == r_count_21_io_out ? io_r_313_b : _GEN_16152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16154 = 10'h13a == r_count_21_io_out ? io_r_314_b : _GEN_16153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16155 = 10'h13b == r_count_21_io_out ? io_r_315_b : _GEN_16154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16156 = 10'h13c == r_count_21_io_out ? io_r_316_b : _GEN_16155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16157 = 10'h13d == r_count_21_io_out ? io_r_317_b : _GEN_16156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16158 = 10'h13e == r_count_21_io_out ? io_r_318_b : _GEN_16157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16159 = 10'h13f == r_count_21_io_out ? io_r_319_b : _GEN_16158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16160 = 10'h140 == r_count_21_io_out ? io_r_320_b : _GEN_16159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16161 = 10'h141 == r_count_21_io_out ? io_r_321_b : _GEN_16160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16162 = 10'h142 == r_count_21_io_out ? io_r_322_b : _GEN_16161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16163 = 10'h143 == r_count_21_io_out ? io_r_323_b : _GEN_16162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16164 = 10'h144 == r_count_21_io_out ? io_r_324_b : _GEN_16163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16165 = 10'h145 == r_count_21_io_out ? io_r_325_b : _GEN_16164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16166 = 10'h146 == r_count_21_io_out ? io_r_326_b : _GEN_16165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16167 = 10'h147 == r_count_21_io_out ? io_r_327_b : _GEN_16166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16168 = 10'h148 == r_count_21_io_out ? io_r_328_b : _GEN_16167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16169 = 10'h149 == r_count_21_io_out ? io_r_329_b : _GEN_16168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16170 = 10'h14a == r_count_21_io_out ? io_r_330_b : _GEN_16169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16171 = 10'h14b == r_count_21_io_out ? io_r_331_b : _GEN_16170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16172 = 10'h14c == r_count_21_io_out ? io_r_332_b : _GEN_16171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16173 = 10'h14d == r_count_21_io_out ? io_r_333_b : _GEN_16172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16174 = 10'h14e == r_count_21_io_out ? io_r_334_b : _GEN_16173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16175 = 10'h14f == r_count_21_io_out ? io_r_335_b : _GEN_16174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16176 = 10'h150 == r_count_21_io_out ? io_r_336_b : _GEN_16175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16177 = 10'h151 == r_count_21_io_out ? io_r_337_b : _GEN_16176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16178 = 10'h152 == r_count_21_io_out ? io_r_338_b : _GEN_16177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16179 = 10'h153 == r_count_21_io_out ? io_r_339_b : _GEN_16178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16180 = 10'h154 == r_count_21_io_out ? io_r_340_b : _GEN_16179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16181 = 10'h155 == r_count_21_io_out ? io_r_341_b : _GEN_16180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16182 = 10'h156 == r_count_21_io_out ? io_r_342_b : _GEN_16181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16183 = 10'h157 == r_count_21_io_out ? io_r_343_b : _GEN_16182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16184 = 10'h158 == r_count_21_io_out ? io_r_344_b : _GEN_16183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16185 = 10'h159 == r_count_21_io_out ? io_r_345_b : _GEN_16184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16186 = 10'h15a == r_count_21_io_out ? io_r_346_b : _GEN_16185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16187 = 10'h15b == r_count_21_io_out ? io_r_347_b : _GEN_16186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16188 = 10'h15c == r_count_21_io_out ? io_r_348_b : _GEN_16187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16189 = 10'h15d == r_count_21_io_out ? io_r_349_b : _GEN_16188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16190 = 10'h15e == r_count_21_io_out ? io_r_350_b : _GEN_16189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16191 = 10'h15f == r_count_21_io_out ? io_r_351_b : _GEN_16190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16192 = 10'h160 == r_count_21_io_out ? io_r_352_b : _GEN_16191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16193 = 10'h161 == r_count_21_io_out ? io_r_353_b : _GEN_16192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16194 = 10'h162 == r_count_21_io_out ? io_r_354_b : _GEN_16193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16195 = 10'h163 == r_count_21_io_out ? io_r_355_b : _GEN_16194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16196 = 10'h164 == r_count_21_io_out ? io_r_356_b : _GEN_16195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16197 = 10'h165 == r_count_21_io_out ? io_r_357_b : _GEN_16196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16198 = 10'h166 == r_count_21_io_out ? io_r_358_b : _GEN_16197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16199 = 10'h167 == r_count_21_io_out ? io_r_359_b : _GEN_16198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16200 = 10'h168 == r_count_21_io_out ? io_r_360_b : _GEN_16199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16201 = 10'h169 == r_count_21_io_out ? io_r_361_b : _GEN_16200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16202 = 10'h16a == r_count_21_io_out ? io_r_362_b : _GEN_16201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16203 = 10'h16b == r_count_21_io_out ? io_r_363_b : _GEN_16202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16204 = 10'h16c == r_count_21_io_out ? io_r_364_b : _GEN_16203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16205 = 10'h16d == r_count_21_io_out ? io_r_365_b : _GEN_16204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16206 = 10'h16e == r_count_21_io_out ? io_r_366_b : _GEN_16205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16207 = 10'h16f == r_count_21_io_out ? io_r_367_b : _GEN_16206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16208 = 10'h170 == r_count_21_io_out ? io_r_368_b : _GEN_16207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16209 = 10'h171 == r_count_21_io_out ? io_r_369_b : _GEN_16208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16210 = 10'h172 == r_count_21_io_out ? io_r_370_b : _GEN_16209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16211 = 10'h173 == r_count_21_io_out ? io_r_371_b : _GEN_16210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16212 = 10'h174 == r_count_21_io_out ? io_r_372_b : _GEN_16211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16213 = 10'h175 == r_count_21_io_out ? io_r_373_b : _GEN_16212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16214 = 10'h176 == r_count_21_io_out ? io_r_374_b : _GEN_16213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16215 = 10'h177 == r_count_21_io_out ? io_r_375_b : _GEN_16214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16216 = 10'h178 == r_count_21_io_out ? io_r_376_b : _GEN_16215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16217 = 10'h179 == r_count_21_io_out ? io_r_377_b : _GEN_16216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16218 = 10'h17a == r_count_21_io_out ? io_r_378_b : _GEN_16217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16219 = 10'h17b == r_count_21_io_out ? io_r_379_b : _GEN_16218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16220 = 10'h17c == r_count_21_io_out ? io_r_380_b : _GEN_16219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16221 = 10'h17d == r_count_21_io_out ? io_r_381_b : _GEN_16220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16222 = 10'h17e == r_count_21_io_out ? io_r_382_b : _GEN_16221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16223 = 10'h17f == r_count_21_io_out ? io_r_383_b : _GEN_16222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16224 = 10'h180 == r_count_21_io_out ? io_r_384_b : _GEN_16223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16225 = 10'h181 == r_count_21_io_out ? io_r_385_b : _GEN_16224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16226 = 10'h182 == r_count_21_io_out ? io_r_386_b : _GEN_16225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16227 = 10'h183 == r_count_21_io_out ? io_r_387_b : _GEN_16226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16228 = 10'h184 == r_count_21_io_out ? io_r_388_b : _GEN_16227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16229 = 10'h185 == r_count_21_io_out ? io_r_389_b : _GEN_16228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16230 = 10'h186 == r_count_21_io_out ? io_r_390_b : _GEN_16229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16231 = 10'h187 == r_count_21_io_out ? io_r_391_b : _GEN_16230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16232 = 10'h188 == r_count_21_io_out ? io_r_392_b : _GEN_16231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16233 = 10'h189 == r_count_21_io_out ? io_r_393_b : _GEN_16232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16234 = 10'h18a == r_count_21_io_out ? io_r_394_b : _GEN_16233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16235 = 10'h18b == r_count_21_io_out ? io_r_395_b : _GEN_16234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16236 = 10'h18c == r_count_21_io_out ? io_r_396_b : _GEN_16235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16237 = 10'h18d == r_count_21_io_out ? io_r_397_b : _GEN_16236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16238 = 10'h18e == r_count_21_io_out ? io_r_398_b : _GEN_16237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16239 = 10'h18f == r_count_21_io_out ? io_r_399_b : _GEN_16238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16240 = 10'h190 == r_count_21_io_out ? io_r_400_b : _GEN_16239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16241 = 10'h191 == r_count_21_io_out ? io_r_401_b : _GEN_16240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16242 = 10'h192 == r_count_21_io_out ? io_r_402_b : _GEN_16241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16243 = 10'h193 == r_count_21_io_out ? io_r_403_b : _GEN_16242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16244 = 10'h194 == r_count_21_io_out ? io_r_404_b : _GEN_16243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16245 = 10'h195 == r_count_21_io_out ? io_r_405_b : _GEN_16244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16246 = 10'h196 == r_count_21_io_out ? io_r_406_b : _GEN_16245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16247 = 10'h197 == r_count_21_io_out ? io_r_407_b : _GEN_16246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16248 = 10'h198 == r_count_21_io_out ? io_r_408_b : _GEN_16247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16249 = 10'h199 == r_count_21_io_out ? io_r_409_b : _GEN_16248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16250 = 10'h19a == r_count_21_io_out ? io_r_410_b : _GEN_16249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16251 = 10'h19b == r_count_21_io_out ? io_r_411_b : _GEN_16250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16252 = 10'h19c == r_count_21_io_out ? io_r_412_b : _GEN_16251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16253 = 10'h19d == r_count_21_io_out ? io_r_413_b : _GEN_16252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16254 = 10'h19e == r_count_21_io_out ? io_r_414_b : _GEN_16253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16255 = 10'h19f == r_count_21_io_out ? io_r_415_b : _GEN_16254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16256 = 10'h1a0 == r_count_21_io_out ? io_r_416_b : _GEN_16255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16257 = 10'h1a1 == r_count_21_io_out ? io_r_417_b : _GEN_16256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16258 = 10'h1a2 == r_count_21_io_out ? io_r_418_b : _GEN_16257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16259 = 10'h1a3 == r_count_21_io_out ? io_r_419_b : _GEN_16258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16260 = 10'h1a4 == r_count_21_io_out ? io_r_420_b : _GEN_16259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16261 = 10'h1a5 == r_count_21_io_out ? io_r_421_b : _GEN_16260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16262 = 10'h1a6 == r_count_21_io_out ? io_r_422_b : _GEN_16261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16263 = 10'h1a7 == r_count_21_io_out ? io_r_423_b : _GEN_16262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16264 = 10'h1a8 == r_count_21_io_out ? io_r_424_b : _GEN_16263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16265 = 10'h1a9 == r_count_21_io_out ? io_r_425_b : _GEN_16264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16266 = 10'h1aa == r_count_21_io_out ? io_r_426_b : _GEN_16265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16267 = 10'h1ab == r_count_21_io_out ? io_r_427_b : _GEN_16266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16268 = 10'h1ac == r_count_21_io_out ? io_r_428_b : _GEN_16267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16269 = 10'h1ad == r_count_21_io_out ? io_r_429_b : _GEN_16268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16270 = 10'h1ae == r_count_21_io_out ? io_r_430_b : _GEN_16269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16271 = 10'h1af == r_count_21_io_out ? io_r_431_b : _GEN_16270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16272 = 10'h1b0 == r_count_21_io_out ? io_r_432_b : _GEN_16271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16273 = 10'h1b1 == r_count_21_io_out ? io_r_433_b : _GEN_16272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16274 = 10'h1b2 == r_count_21_io_out ? io_r_434_b : _GEN_16273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16275 = 10'h1b3 == r_count_21_io_out ? io_r_435_b : _GEN_16274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16276 = 10'h1b4 == r_count_21_io_out ? io_r_436_b : _GEN_16275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16277 = 10'h1b5 == r_count_21_io_out ? io_r_437_b : _GEN_16276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16278 = 10'h1b6 == r_count_21_io_out ? io_r_438_b : _GEN_16277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16279 = 10'h1b7 == r_count_21_io_out ? io_r_439_b : _GEN_16278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16280 = 10'h1b8 == r_count_21_io_out ? io_r_440_b : _GEN_16279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16281 = 10'h1b9 == r_count_21_io_out ? io_r_441_b : _GEN_16280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16282 = 10'h1ba == r_count_21_io_out ? io_r_442_b : _GEN_16281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16283 = 10'h1bb == r_count_21_io_out ? io_r_443_b : _GEN_16282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16284 = 10'h1bc == r_count_21_io_out ? io_r_444_b : _GEN_16283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16285 = 10'h1bd == r_count_21_io_out ? io_r_445_b : _GEN_16284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16286 = 10'h1be == r_count_21_io_out ? io_r_446_b : _GEN_16285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16287 = 10'h1bf == r_count_21_io_out ? io_r_447_b : _GEN_16286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16288 = 10'h1c0 == r_count_21_io_out ? io_r_448_b : _GEN_16287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16289 = 10'h1c1 == r_count_21_io_out ? io_r_449_b : _GEN_16288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16290 = 10'h1c2 == r_count_21_io_out ? io_r_450_b : _GEN_16289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16291 = 10'h1c3 == r_count_21_io_out ? io_r_451_b : _GEN_16290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16292 = 10'h1c4 == r_count_21_io_out ? io_r_452_b : _GEN_16291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16293 = 10'h1c5 == r_count_21_io_out ? io_r_453_b : _GEN_16292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16294 = 10'h1c6 == r_count_21_io_out ? io_r_454_b : _GEN_16293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16295 = 10'h1c7 == r_count_21_io_out ? io_r_455_b : _GEN_16294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16296 = 10'h1c8 == r_count_21_io_out ? io_r_456_b : _GEN_16295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16297 = 10'h1c9 == r_count_21_io_out ? io_r_457_b : _GEN_16296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16298 = 10'h1ca == r_count_21_io_out ? io_r_458_b : _GEN_16297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16299 = 10'h1cb == r_count_21_io_out ? io_r_459_b : _GEN_16298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16300 = 10'h1cc == r_count_21_io_out ? io_r_460_b : _GEN_16299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16301 = 10'h1cd == r_count_21_io_out ? io_r_461_b : _GEN_16300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16302 = 10'h1ce == r_count_21_io_out ? io_r_462_b : _GEN_16301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16303 = 10'h1cf == r_count_21_io_out ? io_r_463_b : _GEN_16302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16304 = 10'h1d0 == r_count_21_io_out ? io_r_464_b : _GEN_16303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16305 = 10'h1d1 == r_count_21_io_out ? io_r_465_b : _GEN_16304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16306 = 10'h1d2 == r_count_21_io_out ? io_r_466_b : _GEN_16305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16307 = 10'h1d3 == r_count_21_io_out ? io_r_467_b : _GEN_16306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16308 = 10'h1d4 == r_count_21_io_out ? io_r_468_b : _GEN_16307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16309 = 10'h1d5 == r_count_21_io_out ? io_r_469_b : _GEN_16308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16310 = 10'h1d6 == r_count_21_io_out ? io_r_470_b : _GEN_16309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16311 = 10'h1d7 == r_count_21_io_out ? io_r_471_b : _GEN_16310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16312 = 10'h1d8 == r_count_21_io_out ? io_r_472_b : _GEN_16311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16313 = 10'h1d9 == r_count_21_io_out ? io_r_473_b : _GEN_16312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16314 = 10'h1da == r_count_21_io_out ? io_r_474_b : _GEN_16313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16315 = 10'h1db == r_count_21_io_out ? io_r_475_b : _GEN_16314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16316 = 10'h1dc == r_count_21_io_out ? io_r_476_b : _GEN_16315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16317 = 10'h1dd == r_count_21_io_out ? io_r_477_b : _GEN_16316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16318 = 10'h1de == r_count_21_io_out ? io_r_478_b : _GEN_16317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16319 = 10'h1df == r_count_21_io_out ? io_r_479_b : _GEN_16318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16320 = 10'h1e0 == r_count_21_io_out ? io_r_480_b : _GEN_16319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16321 = 10'h1e1 == r_count_21_io_out ? io_r_481_b : _GEN_16320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16322 = 10'h1e2 == r_count_21_io_out ? io_r_482_b : _GEN_16321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16323 = 10'h1e3 == r_count_21_io_out ? io_r_483_b : _GEN_16322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16324 = 10'h1e4 == r_count_21_io_out ? io_r_484_b : _GEN_16323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16325 = 10'h1e5 == r_count_21_io_out ? io_r_485_b : _GEN_16324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16326 = 10'h1e6 == r_count_21_io_out ? io_r_486_b : _GEN_16325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16327 = 10'h1e7 == r_count_21_io_out ? io_r_487_b : _GEN_16326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16328 = 10'h1e8 == r_count_21_io_out ? io_r_488_b : _GEN_16327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16329 = 10'h1e9 == r_count_21_io_out ? io_r_489_b : _GEN_16328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16330 = 10'h1ea == r_count_21_io_out ? io_r_490_b : _GEN_16329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16331 = 10'h1eb == r_count_21_io_out ? io_r_491_b : _GEN_16330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16332 = 10'h1ec == r_count_21_io_out ? io_r_492_b : _GEN_16331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16333 = 10'h1ed == r_count_21_io_out ? io_r_493_b : _GEN_16332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16334 = 10'h1ee == r_count_21_io_out ? io_r_494_b : _GEN_16333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16335 = 10'h1ef == r_count_21_io_out ? io_r_495_b : _GEN_16334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16336 = 10'h1f0 == r_count_21_io_out ? io_r_496_b : _GEN_16335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16337 = 10'h1f1 == r_count_21_io_out ? io_r_497_b : _GEN_16336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16338 = 10'h1f2 == r_count_21_io_out ? io_r_498_b : _GEN_16337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16339 = 10'h1f3 == r_count_21_io_out ? io_r_499_b : _GEN_16338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16340 = 10'h1f4 == r_count_21_io_out ? io_r_500_b : _GEN_16339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16341 = 10'h1f5 == r_count_21_io_out ? io_r_501_b : _GEN_16340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16342 = 10'h1f6 == r_count_21_io_out ? io_r_502_b : _GEN_16341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16343 = 10'h1f7 == r_count_21_io_out ? io_r_503_b : _GEN_16342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16344 = 10'h1f8 == r_count_21_io_out ? io_r_504_b : _GEN_16343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16345 = 10'h1f9 == r_count_21_io_out ? io_r_505_b : _GEN_16344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16346 = 10'h1fa == r_count_21_io_out ? io_r_506_b : _GEN_16345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16347 = 10'h1fb == r_count_21_io_out ? io_r_507_b : _GEN_16346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16348 = 10'h1fc == r_count_21_io_out ? io_r_508_b : _GEN_16347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16349 = 10'h1fd == r_count_21_io_out ? io_r_509_b : _GEN_16348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16350 = 10'h1fe == r_count_21_io_out ? io_r_510_b : _GEN_16349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16351 = 10'h1ff == r_count_21_io_out ? io_r_511_b : _GEN_16350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16352 = 10'h200 == r_count_21_io_out ? io_r_512_b : _GEN_16351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16353 = 10'h201 == r_count_21_io_out ? io_r_513_b : _GEN_16352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16354 = 10'h202 == r_count_21_io_out ? io_r_514_b : _GEN_16353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16355 = 10'h203 == r_count_21_io_out ? io_r_515_b : _GEN_16354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16356 = 10'h204 == r_count_21_io_out ? io_r_516_b : _GEN_16355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16357 = 10'h205 == r_count_21_io_out ? io_r_517_b : _GEN_16356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16358 = 10'h206 == r_count_21_io_out ? io_r_518_b : _GEN_16357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16359 = 10'h207 == r_count_21_io_out ? io_r_519_b : _GEN_16358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16360 = 10'h208 == r_count_21_io_out ? io_r_520_b : _GEN_16359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16361 = 10'h209 == r_count_21_io_out ? io_r_521_b : _GEN_16360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16362 = 10'h20a == r_count_21_io_out ? io_r_522_b : _GEN_16361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16363 = 10'h20b == r_count_21_io_out ? io_r_523_b : _GEN_16362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16364 = 10'h20c == r_count_21_io_out ? io_r_524_b : _GEN_16363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16365 = 10'h20d == r_count_21_io_out ? io_r_525_b : _GEN_16364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16366 = 10'h20e == r_count_21_io_out ? io_r_526_b : _GEN_16365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16367 = 10'h20f == r_count_21_io_out ? io_r_527_b : _GEN_16366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16368 = 10'h210 == r_count_21_io_out ? io_r_528_b : _GEN_16367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16369 = 10'h211 == r_count_21_io_out ? io_r_529_b : _GEN_16368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16370 = 10'h212 == r_count_21_io_out ? io_r_530_b : _GEN_16369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16371 = 10'h213 == r_count_21_io_out ? io_r_531_b : _GEN_16370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16372 = 10'h214 == r_count_21_io_out ? io_r_532_b : _GEN_16371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16373 = 10'h215 == r_count_21_io_out ? io_r_533_b : _GEN_16372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16374 = 10'h216 == r_count_21_io_out ? io_r_534_b : _GEN_16373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16375 = 10'h217 == r_count_21_io_out ? io_r_535_b : _GEN_16374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16376 = 10'h218 == r_count_21_io_out ? io_r_536_b : _GEN_16375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16377 = 10'h219 == r_count_21_io_out ? io_r_537_b : _GEN_16376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16378 = 10'h21a == r_count_21_io_out ? io_r_538_b : _GEN_16377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16379 = 10'h21b == r_count_21_io_out ? io_r_539_b : _GEN_16378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16380 = 10'h21c == r_count_21_io_out ? io_r_540_b : _GEN_16379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16381 = 10'h21d == r_count_21_io_out ? io_r_541_b : _GEN_16380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16382 = 10'h21e == r_count_21_io_out ? io_r_542_b : _GEN_16381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16383 = 10'h21f == r_count_21_io_out ? io_r_543_b : _GEN_16382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16384 = 10'h220 == r_count_21_io_out ? io_r_544_b : _GEN_16383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16385 = 10'h221 == r_count_21_io_out ? io_r_545_b : _GEN_16384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16386 = 10'h222 == r_count_21_io_out ? io_r_546_b : _GEN_16385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16387 = 10'h223 == r_count_21_io_out ? io_r_547_b : _GEN_16386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16388 = 10'h224 == r_count_21_io_out ? io_r_548_b : _GEN_16387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16389 = 10'h225 == r_count_21_io_out ? io_r_549_b : _GEN_16388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16390 = 10'h226 == r_count_21_io_out ? io_r_550_b : _GEN_16389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16391 = 10'h227 == r_count_21_io_out ? io_r_551_b : _GEN_16390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16392 = 10'h228 == r_count_21_io_out ? io_r_552_b : _GEN_16391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16393 = 10'h229 == r_count_21_io_out ? io_r_553_b : _GEN_16392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16394 = 10'h22a == r_count_21_io_out ? io_r_554_b : _GEN_16393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16395 = 10'h22b == r_count_21_io_out ? io_r_555_b : _GEN_16394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16396 = 10'h22c == r_count_21_io_out ? io_r_556_b : _GEN_16395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16397 = 10'h22d == r_count_21_io_out ? io_r_557_b : _GEN_16396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16398 = 10'h22e == r_count_21_io_out ? io_r_558_b : _GEN_16397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16399 = 10'h22f == r_count_21_io_out ? io_r_559_b : _GEN_16398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16400 = 10'h230 == r_count_21_io_out ? io_r_560_b : _GEN_16399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16401 = 10'h231 == r_count_21_io_out ? io_r_561_b : _GEN_16400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16402 = 10'h232 == r_count_21_io_out ? io_r_562_b : _GEN_16401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16403 = 10'h233 == r_count_21_io_out ? io_r_563_b : _GEN_16402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16404 = 10'h234 == r_count_21_io_out ? io_r_564_b : _GEN_16403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16405 = 10'h235 == r_count_21_io_out ? io_r_565_b : _GEN_16404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16406 = 10'h236 == r_count_21_io_out ? io_r_566_b : _GEN_16405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16407 = 10'h237 == r_count_21_io_out ? io_r_567_b : _GEN_16406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16408 = 10'h238 == r_count_21_io_out ? io_r_568_b : _GEN_16407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16409 = 10'h239 == r_count_21_io_out ? io_r_569_b : _GEN_16408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16410 = 10'h23a == r_count_21_io_out ? io_r_570_b : _GEN_16409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16411 = 10'h23b == r_count_21_io_out ? io_r_571_b : _GEN_16410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16412 = 10'h23c == r_count_21_io_out ? io_r_572_b : _GEN_16411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16413 = 10'h23d == r_count_21_io_out ? io_r_573_b : _GEN_16412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16414 = 10'h23e == r_count_21_io_out ? io_r_574_b : _GEN_16413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16415 = 10'h23f == r_count_21_io_out ? io_r_575_b : _GEN_16414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16416 = 10'h240 == r_count_21_io_out ? io_r_576_b : _GEN_16415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16417 = 10'h241 == r_count_21_io_out ? io_r_577_b : _GEN_16416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16418 = 10'h242 == r_count_21_io_out ? io_r_578_b : _GEN_16417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16419 = 10'h243 == r_count_21_io_out ? io_r_579_b : _GEN_16418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16420 = 10'h244 == r_count_21_io_out ? io_r_580_b : _GEN_16419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16421 = 10'h245 == r_count_21_io_out ? io_r_581_b : _GEN_16420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16422 = 10'h246 == r_count_21_io_out ? io_r_582_b : _GEN_16421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16423 = 10'h247 == r_count_21_io_out ? io_r_583_b : _GEN_16422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16424 = 10'h248 == r_count_21_io_out ? io_r_584_b : _GEN_16423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16425 = 10'h249 == r_count_21_io_out ? io_r_585_b : _GEN_16424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16426 = 10'h24a == r_count_21_io_out ? io_r_586_b : _GEN_16425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16427 = 10'h24b == r_count_21_io_out ? io_r_587_b : _GEN_16426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16428 = 10'h24c == r_count_21_io_out ? io_r_588_b : _GEN_16427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16429 = 10'h24d == r_count_21_io_out ? io_r_589_b : _GEN_16428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16430 = 10'h24e == r_count_21_io_out ? io_r_590_b : _GEN_16429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16431 = 10'h24f == r_count_21_io_out ? io_r_591_b : _GEN_16430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16432 = 10'h250 == r_count_21_io_out ? io_r_592_b : _GEN_16431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16433 = 10'h251 == r_count_21_io_out ? io_r_593_b : _GEN_16432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16434 = 10'h252 == r_count_21_io_out ? io_r_594_b : _GEN_16433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16435 = 10'h253 == r_count_21_io_out ? io_r_595_b : _GEN_16434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16436 = 10'h254 == r_count_21_io_out ? io_r_596_b : _GEN_16435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16437 = 10'h255 == r_count_21_io_out ? io_r_597_b : _GEN_16436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16438 = 10'h256 == r_count_21_io_out ? io_r_598_b : _GEN_16437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16439 = 10'h257 == r_count_21_io_out ? io_r_599_b : _GEN_16438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16440 = 10'h258 == r_count_21_io_out ? io_r_600_b : _GEN_16439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16441 = 10'h259 == r_count_21_io_out ? io_r_601_b : _GEN_16440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16442 = 10'h25a == r_count_21_io_out ? io_r_602_b : _GEN_16441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16443 = 10'h25b == r_count_21_io_out ? io_r_603_b : _GEN_16442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16444 = 10'h25c == r_count_21_io_out ? io_r_604_b : _GEN_16443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16445 = 10'h25d == r_count_21_io_out ? io_r_605_b : _GEN_16444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16446 = 10'h25e == r_count_21_io_out ? io_r_606_b : _GEN_16445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16447 = 10'h25f == r_count_21_io_out ? io_r_607_b : _GEN_16446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16448 = 10'h260 == r_count_21_io_out ? io_r_608_b : _GEN_16447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16449 = 10'h261 == r_count_21_io_out ? io_r_609_b : _GEN_16448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16450 = 10'h262 == r_count_21_io_out ? io_r_610_b : _GEN_16449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16451 = 10'h263 == r_count_21_io_out ? io_r_611_b : _GEN_16450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16452 = 10'h264 == r_count_21_io_out ? io_r_612_b : _GEN_16451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16453 = 10'h265 == r_count_21_io_out ? io_r_613_b : _GEN_16452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16454 = 10'h266 == r_count_21_io_out ? io_r_614_b : _GEN_16453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16455 = 10'h267 == r_count_21_io_out ? io_r_615_b : _GEN_16454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16456 = 10'h268 == r_count_21_io_out ? io_r_616_b : _GEN_16455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16457 = 10'h269 == r_count_21_io_out ? io_r_617_b : _GEN_16456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16458 = 10'h26a == r_count_21_io_out ? io_r_618_b : _GEN_16457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16459 = 10'h26b == r_count_21_io_out ? io_r_619_b : _GEN_16458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16460 = 10'h26c == r_count_21_io_out ? io_r_620_b : _GEN_16459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16461 = 10'h26d == r_count_21_io_out ? io_r_621_b : _GEN_16460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16462 = 10'h26e == r_count_21_io_out ? io_r_622_b : _GEN_16461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16463 = 10'h26f == r_count_21_io_out ? io_r_623_b : _GEN_16462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16464 = 10'h270 == r_count_21_io_out ? io_r_624_b : _GEN_16463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16465 = 10'h271 == r_count_21_io_out ? io_r_625_b : _GEN_16464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16466 = 10'h272 == r_count_21_io_out ? io_r_626_b : _GEN_16465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16467 = 10'h273 == r_count_21_io_out ? io_r_627_b : _GEN_16466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16468 = 10'h274 == r_count_21_io_out ? io_r_628_b : _GEN_16467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16469 = 10'h275 == r_count_21_io_out ? io_r_629_b : _GEN_16468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16470 = 10'h276 == r_count_21_io_out ? io_r_630_b : _GEN_16469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16471 = 10'h277 == r_count_21_io_out ? io_r_631_b : _GEN_16470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16472 = 10'h278 == r_count_21_io_out ? io_r_632_b : _GEN_16471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16473 = 10'h279 == r_count_21_io_out ? io_r_633_b : _GEN_16472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16474 = 10'h27a == r_count_21_io_out ? io_r_634_b : _GEN_16473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16475 = 10'h27b == r_count_21_io_out ? io_r_635_b : _GEN_16474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16476 = 10'h27c == r_count_21_io_out ? io_r_636_b : _GEN_16475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16477 = 10'h27d == r_count_21_io_out ? io_r_637_b : _GEN_16476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16478 = 10'h27e == r_count_21_io_out ? io_r_638_b : _GEN_16477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16479 = 10'h27f == r_count_21_io_out ? io_r_639_b : _GEN_16478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16480 = 10'h280 == r_count_21_io_out ? io_r_640_b : _GEN_16479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16481 = 10'h281 == r_count_21_io_out ? io_r_641_b : _GEN_16480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16482 = 10'h282 == r_count_21_io_out ? io_r_642_b : _GEN_16481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16483 = 10'h283 == r_count_21_io_out ? io_r_643_b : _GEN_16482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16484 = 10'h284 == r_count_21_io_out ? io_r_644_b : _GEN_16483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16485 = 10'h285 == r_count_21_io_out ? io_r_645_b : _GEN_16484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16486 = 10'h286 == r_count_21_io_out ? io_r_646_b : _GEN_16485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16487 = 10'h287 == r_count_21_io_out ? io_r_647_b : _GEN_16486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16488 = 10'h288 == r_count_21_io_out ? io_r_648_b : _GEN_16487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16489 = 10'h289 == r_count_21_io_out ? io_r_649_b : _GEN_16488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16490 = 10'h28a == r_count_21_io_out ? io_r_650_b : _GEN_16489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16491 = 10'h28b == r_count_21_io_out ? io_r_651_b : _GEN_16490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16492 = 10'h28c == r_count_21_io_out ? io_r_652_b : _GEN_16491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16493 = 10'h28d == r_count_21_io_out ? io_r_653_b : _GEN_16492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16494 = 10'h28e == r_count_21_io_out ? io_r_654_b : _GEN_16493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16495 = 10'h28f == r_count_21_io_out ? io_r_655_b : _GEN_16494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16496 = 10'h290 == r_count_21_io_out ? io_r_656_b : _GEN_16495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16497 = 10'h291 == r_count_21_io_out ? io_r_657_b : _GEN_16496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16498 = 10'h292 == r_count_21_io_out ? io_r_658_b : _GEN_16497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16499 = 10'h293 == r_count_21_io_out ? io_r_659_b : _GEN_16498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16500 = 10'h294 == r_count_21_io_out ? io_r_660_b : _GEN_16499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16501 = 10'h295 == r_count_21_io_out ? io_r_661_b : _GEN_16500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16502 = 10'h296 == r_count_21_io_out ? io_r_662_b : _GEN_16501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16503 = 10'h297 == r_count_21_io_out ? io_r_663_b : _GEN_16502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16504 = 10'h298 == r_count_21_io_out ? io_r_664_b : _GEN_16503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16505 = 10'h299 == r_count_21_io_out ? io_r_665_b : _GEN_16504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16506 = 10'h29a == r_count_21_io_out ? io_r_666_b : _GEN_16505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16507 = 10'h29b == r_count_21_io_out ? io_r_667_b : _GEN_16506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16508 = 10'h29c == r_count_21_io_out ? io_r_668_b : _GEN_16507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16509 = 10'h29d == r_count_21_io_out ? io_r_669_b : _GEN_16508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16510 = 10'h29e == r_count_21_io_out ? io_r_670_b : _GEN_16509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16511 = 10'h29f == r_count_21_io_out ? io_r_671_b : _GEN_16510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16512 = 10'h2a0 == r_count_21_io_out ? io_r_672_b : _GEN_16511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16513 = 10'h2a1 == r_count_21_io_out ? io_r_673_b : _GEN_16512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16514 = 10'h2a2 == r_count_21_io_out ? io_r_674_b : _GEN_16513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16515 = 10'h2a3 == r_count_21_io_out ? io_r_675_b : _GEN_16514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16516 = 10'h2a4 == r_count_21_io_out ? io_r_676_b : _GEN_16515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16517 = 10'h2a5 == r_count_21_io_out ? io_r_677_b : _GEN_16516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16518 = 10'h2a6 == r_count_21_io_out ? io_r_678_b : _GEN_16517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16519 = 10'h2a7 == r_count_21_io_out ? io_r_679_b : _GEN_16518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16520 = 10'h2a8 == r_count_21_io_out ? io_r_680_b : _GEN_16519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16521 = 10'h2a9 == r_count_21_io_out ? io_r_681_b : _GEN_16520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16522 = 10'h2aa == r_count_21_io_out ? io_r_682_b : _GEN_16521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16523 = 10'h2ab == r_count_21_io_out ? io_r_683_b : _GEN_16522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16524 = 10'h2ac == r_count_21_io_out ? io_r_684_b : _GEN_16523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16525 = 10'h2ad == r_count_21_io_out ? io_r_685_b : _GEN_16524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16526 = 10'h2ae == r_count_21_io_out ? io_r_686_b : _GEN_16525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16527 = 10'h2af == r_count_21_io_out ? io_r_687_b : _GEN_16526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16528 = 10'h2b0 == r_count_21_io_out ? io_r_688_b : _GEN_16527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16529 = 10'h2b1 == r_count_21_io_out ? io_r_689_b : _GEN_16528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16530 = 10'h2b2 == r_count_21_io_out ? io_r_690_b : _GEN_16529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16531 = 10'h2b3 == r_count_21_io_out ? io_r_691_b : _GEN_16530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16532 = 10'h2b4 == r_count_21_io_out ? io_r_692_b : _GEN_16531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16533 = 10'h2b5 == r_count_21_io_out ? io_r_693_b : _GEN_16532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16534 = 10'h2b6 == r_count_21_io_out ? io_r_694_b : _GEN_16533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16535 = 10'h2b7 == r_count_21_io_out ? io_r_695_b : _GEN_16534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16536 = 10'h2b8 == r_count_21_io_out ? io_r_696_b : _GEN_16535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16537 = 10'h2b9 == r_count_21_io_out ? io_r_697_b : _GEN_16536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16538 = 10'h2ba == r_count_21_io_out ? io_r_698_b : _GEN_16537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16539 = 10'h2bb == r_count_21_io_out ? io_r_699_b : _GEN_16538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16540 = 10'h2bc == r_count_21_io_out ? io_r_700_b : _GEN_16539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16541 = 10'h2bd == r_count_21_io_out ? io_r_701_b : _GEN_16540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16542 = 10'h2be == r_count_21_io_out ? io_r_702_b : _GEN_16541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16543 = 10'h2bf == r_count_21_io_out ? io_r_703_b : _GEN_16542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16544 = 10'h2c0 == r_count_21_io_out ? io_r_704_b : _GEN_16543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16545 = 10'h2c1 == r_count_21_io_out ? io_r_705_b : _GEN_16544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16546 = 10'h2c2 == r_count_21_io_out ? io_r_706_b : _GEN_16545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16547 = 10'h2c3 == r_count_21_io_out ? io_r_707_b : _GEN_16546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16548 = 10'h2c4 == r_count_21_io_out ? io_r_708_b : _GEN_16547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16549 = 10'h2c5 == r_count_21_io_out ? io_r_709_b : _GEN_16548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16550 = 10'h2c6 == r_count_21_io_out ? io_r_710_b : _GEN_16549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16551 = 10'h2c7 == r_count_21_io_out ? io_r_711_b : _GEN_16550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16552 = 10'h2c8 == r_count_21_io_out ? io_r_712_b : _GEN_16551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16553 = 10'h2c9 == r_count_21_io_out ? io_r_713_b : _GEN_16552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16554 = 10'h2ca == r_count_21_io_out ? io_r_714_b : _GEN_16553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16555 = 10'h2cb == r_count_21_io_out ? io_r_715_b : _GEN_16554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16556 = 10'h2cc == r_count_21_io_out ? io_r_716_b : _GEN_16555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16557 = 10'h2cd == r_count_21_io_out ? io_r_717_b : _GEN_16556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16558 = 10'h2ce == r_count_21_io_out ? io_r_718_b : _GEN_16557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16559 = 10'h2cf == r_count_21_io_out ? io_r_719_b : _GEN_16558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16560 = 10'h2d0 == r_count_21_io_out ? io_r_720_b : _GEN_16559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16561 = 10'h2d1 == r_count_21_io_out ? io_r_721_b : _GEN_16560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16562 = 10'h2d2 == r_count_21_io_out ? io_r_722_b : _GEN_16561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16563 = 10'h2d3 == r_count_21_io_out ? io_r_723_b : _GEN_16562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16564 = 10'h2d4 == r_count_21_io_out ? io_r_724_b : _GEN_16563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16565 = 10'h2d5 == r_count_21_io_out ? io_r_725_b : _GEN_16564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16566 = 10'h2d6 == r_count_21_io_out ? io_r_726_b : _GEN_16565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16567 = 10'h2d7 == r_count_21_io_out ? io_r_727_b : _GEN_16566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16568 = 10'h2d8 == r_count_21_io_out ? io_r_728_b : _GEN_16567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16569 = 10'h2d9 == r_count_21_io_out ? io_r_729_b : _GEN_16568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16570 = 10'h2da == r_count_21_io_out ? io_r_730_b : _GEN_16569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16571 = 10'h2db == r_count_21_io_out ? io_r_731_b : _GEN_16570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16572 = 10'h2dc == r_count_21_io_out ? io_r_732_b : _GEN_16571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16573 = 10'h2dd == r_count_21_io_out ? io_r_733_b : _GEN_16572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16574 = 10'h2de == r_count_21_io_out ? io_r_734_b : _GEN_16573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16575 = 10'h2df == r_count_21_io_out ? io_r_735_b : _GEN_16574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16576 = 10'h2e0 == r_count_21_io_out ? io_r_736_b : _GEN_16575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16577 = 10'h2e1 == r_count_21_io_out ? io_r_737_b : _GEN_16576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16578 = 10'h2e2 == r_count_21_io_out ? io_r_738_b : _GEN_16577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16579 = 10'h2e3 == r_count_21_io_out ? io_r_739_b : _GEN_16578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16580 = 10'h2e4 == r_count_21_io_out ? io_r_740_b : _GEN_16579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16581 = 10'h2e5 == r_count_21_io_out ? io_r_741_b : _GEN_16580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16582 = 10'h2e6 == r_count_21_io_out ? io_r_742_b : _GEN_16581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16583 = 10'h2e7 == r_count_21_io_out ? io_r_743_b : _GEN_16582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16584 = 10'h2e8 == r_count_21_io_out ? io_r_744_b : _GEN_16583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16585 = 10'h2e9 == r_count_21_io_out ? io_r_745_b : _GEN_16584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16586 = 10'h2ea == r_count_21_io_out ? io_r_746_b : _GEN_16585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16587 = 10'h2eb == r_count_21_io_out ? io_r_747_b : _GEN_16586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16588 = 10'h2ec == r_count_21_io_out ? io_r_748_b : _GEN_16587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16591 = 10'h1 == r_count_22_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16592 = 10'h2 == r_count_22_io_out ? io_r_2_b : _GEN_16591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16593 = 10'h3 == r_count_22_io_out ? io_r_3_b : _GEN_16592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16594 = 10'h4 == r_count_22_io_out ? io_r_4_b : _GEN_16593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16595 = 10'h5 == r_count_22_io_out ? io_r_5_b : _GEN_16594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16596 = 10'h6 == r_count_22_io_out ? io_r_6_b : _GEN_16595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16597 = 10'h7 == r_count_22_io_out ? io_r_7_b : _GEN_16596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16598 = 10'h8 == r_count_22_io_out ? io_r_8_b : _GEN_16597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16599 = 10'h9 == r_count_22_io_out ? io_r_9_b : _GEN_16598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16600 = 10'ha == r_count_22_io_out ? io_r_10_b : _GEN_16599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16601 = 10'hb == r_count_22_io_out ? io_r_11_b : _GEN_16600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16602 = 10'hc == r_count_22_io_out ? io_r_12_b : _GEN_16601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16603 = 10'hd == r_count_22_io_out ? io_r_13_b : _GEN_16602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16604 = 10'he == r_count_22_io_out ? io_r_14_b : _GEN_16603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16605 = 10'hf == r_count_22_io_out ? io_r_15_b : _GEN_16604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16606 = 10'h10 == r_count_22_io_out ? io_r_16_b : _GEN_16605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16607 = 10'h11 == r_count_22_io_out ? io_r_17_b : _GEN_16606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16608 = 10'h12 == r_count_22_io_out ? io_r_18_b : _GEN_16607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16609 = 10'h13 == r_count_22_io_out ? io_r_19_b : _GEN_16608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16610 = 10'h14 == r_count_22_io_out ? io_r_20_b : _GEN_16609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16611 = 10'h15 == r_count_22_io_out ? io_r_21_b : _GEN_16610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16612 = 10'h16 == r_count_22_io_out ? io_r_22_b : _GEN_16611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16613 = 10'h17 == r_count_22_io_out ? io_r_23_b : _GEN_16612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16614 = 10'h18 == r_count_22_io_out ? io_r_24_b : _GEN_16613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16615 = 10'h19 == r_count_22_io_out ? io_r_25_b : _GEN_16614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16616 = 10'h1a == r_count_22_io_out ? io_r_26_b : _GEN_16615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16617 = 10'h1b == r_count_22_io_out ? io_r_27_b : _GEN_16616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16618 = 10'h1c == r_count_22_io_out ? io_r_28_b : _GEN_16617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16619 = 10'h1d == r_count_22_io_out ? io_r_29_b : _GEN_16618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16620 = 10'h1e == r_count_22_io_out ? io_r_30_b : _GEN_16619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16621 = 10'h1f == r_count_22_io_out ? io_r_31_b : _GEN_16620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16622 = 10'h20 == r_count_22_io_out ? io_r_32_b : _GEN_16621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16623 = 10'h21 == r_count_22_io_out ? io_r_33_b : _GEN_16622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16624 = 10'h22 == r_count_22_io_out ? io_r_34_b : _GEN_16623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16625 = 10'h23 == r_count_22_io_out ? io_r_35_b : _GEN_16624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16626 = 10'h24 == r_count_22_io_out ? io_r_36_b : _GEN_16625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16627 = 10'h25 == r_count_22_io_out ? io_r_37_b : _GEN_16626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16628 = 10'h26 == r_count_22_io_out ? io_r_38_b : _GEN_16627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16629 = 10'h27 == r_count_22_io_out ? io_r_39_b : _GEN_16628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16630 = 10'h28 == r_count_22_io_out ? io_r_40_b : _GEN_16629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16631 = 10'h29 == r_count_22_io_out ? io_r_41_b : _GEN_16630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16632 = 10'h2a == r_count_22_io_out ? io_r_42_b : _GEN_16631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16633 = 10'h2b == r_count_22_io_out ? io_r_43_b : _GEN_16632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16634 = 10'h2c == r_count_22_io_out ? io_r_44_b : _GEN_16633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16635 = 10'h2d == r_count_22_io_out ? io_r_45_b : _GEN_16634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16636 = 10'h2e == r_count_22_io_out ? io_r_46_b : _GEN_16635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16637 = 10'h2f == r_count_22_io_out ? io_r_47_b : _GEN_16636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16638 = 10'h30 == r_count_22_io_out ? io_r_48_b : _GEN_16637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16639 = 10'h31 == r_count_22_io_out ? io_r_49_b : _GEN_16638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16640 = 10'h32 == r_count_22_io_out ? io_r_50_b : _GEN_16639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16641 = 10'h33 == r_count_22_io_out ? io_r_51_b : _GEN_16640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16642 = 10'h34 == r_count_22_io_out ? io_r_52_b : _GEN_16641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16643 = 10'h35 == r_count_22_io_out ? io_r_53_b : _GEN_16642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16644 = 10'h36 == r_count_22_io_out ? io_r_54_b : _GEN_16643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16645 = 10'h37 == r_count_22_io_out ? io_r_55_b : _GEN_16644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16646 = 10'h38 == r_count_22_io_out ? io_r_56_b : _GEN_16645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16647 = 10'h39 == r_count_22_io_out ? io_r_57_b : _GEN_16646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16648 = 10'h3a == r_count_22_io_out ? io_r_58_b : _GEN_16647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16649 = 10'h3b == r_count_22_io_out ? io_r_59_b : _GEN_16648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16650 = 10'h3c == r_count_22_io_out ? io_r_60_b : _GEN_16649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16651 = 10'h3d == r_count_22_io_out ? io_r_61_b : _GEN_16650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16652 = 10'h3e == r_count_22_io_out ? io_r_62_b : _GEN_16651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16653 = 10'h3f == r_count_22_io_out ? io_r_63_b : _GEN_16652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16654 = 10'h40 == r_count_22_io_out ? io_r_64_b : _GEN_16653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16655 = 10'h41 == r_count_22_io_out ? io_r_65_b : _GEN_16654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16656 = 10'h42 == r_count_22_io_out ? io_r_66_b : _GEN_16655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16657 = 10'h43 == r_count_22_io_out ? io_r_67_b : _GEN_16656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16658 = 10'h44 == r_count_22_io_out ? io_r_68_b : _GEN_16657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16659 = 10'h45 == r_count_22_io_out ? io_r_69_b : _GEN_16658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16660 = 10'h46 == r_count_22_io_out ? io_r_70_b : _GEN_16659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16661 = 10'h47 == r_count_22_io_out ? io_r_71_b : _GEN_16660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16662 = 10'h48 == r_count_22_io_out ? io_r_72_b : _GEN_16661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16663 = 10'h49 == r_count_22_io_out ? io_r_73_b : _GEN_16662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16664 = 10'h4a == r_count_22_io_out ? io_r_74_b : _GEN_16663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16665 = 10'h4b == r_count_22_io_out ? io_r_75_b : _GEN_16664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16666 = 10'h4c == r_count_22_io_out ? io_r_76_b : _GEN_16665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16667 = 10'h4d == r_count_22_io_out ? io_r_77_b : _GEN_16666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16668 = 10'h4e == r_count_22_io_out ? io_r_78_b : _GEN_16667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16669 = 10'h4f == r_count_22_io_out ? io_r_79_b : _GEN_16668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16670 = 10'h50 == r_count_22_io_out ? io_r_80_b : _GEN_16669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16671 = 10'h51 == r_count_22_io_out ? io_r_81_b : _GEN_16670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16672 = 10'h52 == r_count_22_io_out ? io_r_82_b : _GEN_16671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16673 = 10'h53 == r_count_22_io_out ? io_r_83_b : _GEN_16672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16674 = 10'h54 == r_count_22_io_out ? io_r_84_b : _GEN_16673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16675 = 10'h55 == r_count_22_io_out ? io_r_85_b : _GEN_16674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16676 = 10'h56 == r_count_22_io_out ? io_r_86_b : _GEN_16675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16677 = 10'h57 == r_count_22_io_out ? io_r_87_b : _GEN_16676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16678 = 10'h58 == r_count_22_io_out ? io_r_88_b : _GEN_16677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16679 = 10'h59 == r_count_22_io_out ? io_r_89_b : _GEN_16678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16680 = 10'h5a == r_count_22_io_out ? io_r_90_b : _GEN_16679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16681 = 10'h5b == r_count_22_io_out ? io_r_91_b : _GEN_16680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16682 = 10'h5c == r_count_22_io_out ? io_r_92_b : _GEN_16681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16683 = 10'h5d == r_count_22_io_out ? io_r_93_b : _GEN_16682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16684 = 10'h5e == r_count_22_io_out ? io_r_94_b : _GEN_16683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16685 = 10'h5f == r_count_22_io_out ? io_r_95_b : _GEN_16684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16686 = 10'h60 == r_count_22_io_out ? io_r_96_b : _GEN_16685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16687 = 10'h61 == r_count_22_io_out ? io_r_97_b : _GEN_16686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16688 = 10'h62 == r_count_22_io_out ? io_r_98_b : _GEN_16687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16689 = 10'h63 == r_count_22_io_out ? io_r_99_b : _GEN_16688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16690 = 10'h64 == r_count_22_io_out ? io_r_100_b : _GEN_16689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16691 = 10'h65 == r_count_22_io_out ? io_r_101_b : _GEN_16690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16692 = 10'h66 == r_count_22_io_out ? io_r_102_b : _GEN_16691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16693 = 10'h67 == r_count_22_io_out ? io_r_103_b : _GEN_16692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16694 = 10'h68 == r_count_22_io_out ? io_r_104_b : _GEN_16693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16695 = 10'h69 == r_count_22_io_out ? io_r_105_b : _GEN_16694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16696 = 10'h6a == r_count_22_io_out ? io_r_106_b : _GEN_16695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16697 = 10'h6b == r_count_22_io_out ? io_r_107_b : _GEN_16696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16698 = 10'h6c == r_count_22_io_out ? io_r_108_b : _GEN_16697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16699 = 10'h6d == r_count_22_io_out ? io_r_109_b : _GEN_16698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16700 = 10'h6e == r_count_22_io_out ? io_r_110_b : _GEN_16699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16701 = 10'h6f == r_count_22_io_out ? io_r_111_b : _GEN_16700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16702 = 10'h70 == r_count_22_io_out ? io_r_112_b : _GEN_16701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16703 = 10'h71 == r_count_22_io_out ? io_r_113_b : _GEN_16702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16704 = 10'h72 == r_count_22_io_out ? io_r_114_b : _GEN_16703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16705 = 10'h73 == r_count_22_io_out ? io_r_115_b : _GEN_16704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16706 = 10'h74 == r_count_22_io_out ? io_r_116_b : _GEN_16705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16707 = 10'h75 == r_count_22_io_out ? io_r_117_b : _GEN_16706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16708 = 10'h76 == r_count_22_io_out ? io_r_118_b : _GEN_16707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16709 = 10'h77 == r_count_22_io_out ? io_r_119_b : _GEN_16708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16710 = 10'h78 == r_count_22_io_out ? io_r_120_b : _GEN_16709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16711 = 10'h79 == r_count_22_io_out ? io_r_121_b : _GEN_16710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16712 = 10'h7a == r_count_22_io_out ? io_r_122_b : _GEN_16711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16713 = 10'h7b == r_count_22_io_out ? io_r_123_b : _GEN_16712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16714 = 10'h7c == r_count_22_io_out ? io_r_124_b : _GEN_16713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16715 = 10'h7d == r_count_22_io_out ? io_r_125_b : _GEN_16714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16716 = 10'h7e == r_count_22_io_out ? io_r_126_b : _GEN_16715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16717 = 10'h7f == r_count_22_io_out ? io_r_127_b : _GEN_16716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16718 = 10'h80 == r_count_22_io_out ? io_r_128_b : _GEN_16717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16719 = 10'h81 == r_count_22_io_out ? io_r_129_b : _GEN_16718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16720 = 10'h82 == r_count_22_io_out ? io_r_130_b : _GEN_16719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16721 = 10'h83 == r_count_22_io_out ? io_r_131_b : _GEN_16720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16722 = 10'h84 == r_count_22_io_out ? io_r_132_b : _GEN_16721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16723 = 10'h85 == r_count_22_io_out ? io_r_133_b : _GEN_16722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16724 = 10'h86 == r_count_22_io_out ? io_r_134_b : _GEN_16723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16725 = 10'h87 == r_count_22_io_out ? io_r_135_b : _GEN_16724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16726 = 10'h88 == r_count_22_io_out ? io_r_136_b : _GEN_16725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16727 = 10'h89 == r_count_22_io_out ? io_r_137_b : _GEN_16726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16728 = 10'h8a == r_count_22_io_out ? io_r_138_b : _GEN_16727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16729 = 10'h8b == r_count_22_io_out ? io_r_139_b : _GEN_16728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16730 = 10'h8c == r_count_22_io_out ? io_r_140_b : _GEN_16729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16731 = 10'h8d == r_count_22_io_out ? io_r_141_b : _GEN_16730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16732 = 10'h8e == r_count_22_io_out ? io_r_142_b : _GEN_16731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16733 = 10'h8f == r_count_22_io_out ? io_r_143_b : _GEN_16732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16734 = 10'h90 == r_count_22_io_out ? io_r_144_b : _GEN_16733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16735 = 10'h91 == r_count_22_io_out ? io_r_145_b : _GEN_16734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16736 = 10'h92 == r_count_22_io_out ? io_r_146_b : _GEN_16735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16737 = 10'h93 == r_count_22_io_out ? io_r_147_b : _GEN_16736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16738 = 10'h94 == r_count_22_io_out ? io_r_148_b : _GEN_16737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16739 = 10'h95 == r_count_22_io_out ? io_r_149_b : _GEN_16738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16740 = 10'h96 == r_count_22_io_out ? io_r_150_b : _GEN_16739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16741 = 10'h97 == r_count_22_io_out ? io_r_151_b : _GEN_16740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16742 = 10'h98 == r_count_22_io_out ? io_r_152_b : _GEN_16741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16743 = 10'h99 == r_count_22_io_out ? io_r_153_b : _GEN_16742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16744 = 10'h9a == r_count_22_io_out ? io_r_154_b : _GEN_16743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16745 = 10'h9b == r_count_22_io_out ? io_r_155_b : _GEN_16744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16746 = 10'h9c == r_count_22_io_out ? io_r_156_b : _GEN_16745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16747 = 10'h9d == r_count_22_io_out ? io_r_157_b : _GEN_16746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16748 = 10'h9e == r_count_22_io_out ? io_r_158_b : _GEN_16747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16749 = 10'h9f == r_count_22_io_out ? io_r_159_b : _GEN_16748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16750 = 10'ha0 == r_count_22_io_out ? io_r_160_b : _GEN_16749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16751 = 10'ha1 == r_count_22_io_out ? io_r_161_b : _GEN_16750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16752 = 10'ha2 == r_count_22_io_out ? io_r_162_b : _GEN_16751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16753 = 10'ha3 == r_count_22_io_out ? io_r_163_b : _GEN_16752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16754 = 10'ha4 == r_count_22_io_out ? io_r_164_b : _GEN_16753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16755 = 10'ha5 == r_count_22_io_out ? io_r_165_b : _GEN_16754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16756 = 10'ha6 == r_count_22_io_out ? io_r_166_b : _GEN_16755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16757 = 10'ha7 == r_count_22_io_out ? io_r_167_b : _GEN_16756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16758 = 10'ha8 == r_count_22_io_out ? io_r_168_b : _GEN_16757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16759 = 10'ha9 == r_count_22_io_out ? io_r_169_b : _GEN_16758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16760 = 10'haa == r_count_22_io_out ? io_r_170_b : _GEN_16759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16761 = 10'hab == r_count_22_io_out ? io_r_171_b : _GEN_16760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16762 = 10'hac == r_count_22_io_out ? io_r_172_b : _GEN_16761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16763 = 10'had == r_count_22_io_out ? io_r_173_b : _GEN_16762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16764 = 10'hae == r_count_22_io_out ? io_r_174_b : _GEN_16763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16765 = 10'haf == r_count_22_io_out ? io_r_175_b : _GEN_16764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16766 = 10'hb0 == r_count_22_io_out ? io_r_176_b : _GEN_16765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16767 = 10'hb1 == r_count_22_io_out ? io_r_177_b : _GEN_16766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16768 = 10'hb2 == r_count_22_io_out ? io_r_178_b : _GEN_16767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16769 = 10'hb3 == r_count_22_io_out ? io_r_179_b : _GEN_16768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16770 = 10'hb4 == r_count_22_io_out ? io_r_180_b : _GEN_16769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16771 = 10'hb5 == r_count_22_io_out ? io_r_181_b : _GEN_16770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16772 = 10'hb6 == r_count_22_io_out ? io_r_182_b : _GEN_16771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16773 = 10'hb7 == r_count_22_io_out ? io_r_183_b : _GEN_16772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16774 = 10'hb8 == r_count_22_io_out ? io_r_184_b : _GEN_16773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16775 = 10'hb9 == r_count_22_io_out ? io_r_185_b : _GEN_16774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16776 = 10'hba == r_count_22_io_out ? io_r_186_b : _GEN_16775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16777 = 10'hbb == r_count_22_io_out ? io_r_187_b : _GEN_16776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16778 = 10'hbc == r_count_22_io_out ? io_r_188_b : _GEN_16777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16779 = 10'hbd == r_count_22_io_out ? io_r_189_b : _GEN_16778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16780 = 10'hbe == r_count_22_io_out ? io_r_190_b : _GEN_16779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16781 = 10'hbf == r_count_22_io_out ? io_r_191_b : _GEN_16780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16782 = 10'hc0 == r_count_22_io_out ? io_r_192_b : _GEN_16781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16783 = 10'hc1 == r_count_22_io_out ? io_r_193_b : _GEN_16782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16784 = 10'hc2 == r_count_22_io_out ? io_r_194_b : _GEN_16783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16785 = 10'hc3 == r_count_22_io_out ? io_r_195_b : _GEN_16784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16786 = 10'hc4 == r_count_22_io_out ? io_r_196_b : _GEN_16785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16787 = 10'hc5 == r_count_22_io_out ? io_r_197_b : _GEN_16786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16788 = 10'hc6 == r_count_22_io_out ? io_r_198_b : _GEN_16787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16789 = 10'hc7 == r_count_22_io_out ? io_r_199_b : _GEN_16788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16790 = 10'hc8 == r_count_22_io_out ? io_r_200_b : _GEN_16789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16791 = 10'hc9 == r_count_22_io_out ? io_r_201_b : _GEN_16790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16792 = 10'hca == r_count_22_io_out ? io_r_202_b : _GEN_16791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16793 = 10'hcb == r_count_22_io_out ? io_r_203_b : _GEN_16792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16794 = 10'hcc == r_count_22_io_out ? io_r_204_b : _GEN_16793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16795 = 10'hcd == r_count_22_io_out ? io_r_205_b : _GEN_16794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16796 = 10'hce == r_count_22_io_out ? io_r_206_b : _GEN_16795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16797 = 10'hcf == r_count_22_io_out ? io_r_207_b : _GEN_16796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16798 = 10'hd0 == r_count_22_io_out ? io_r_208_b : _GEN_16797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16799 = 10'hd1 == r_count_22_io_out ? io_r_209_b : _GEN_16798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16800 = 10'hd2 == r_count_22_io_out ? io_r_210_b : _GEN_16799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16801 = 10'hd3 == r_count_22_io_out ? io_r_211_b : _GEN_16800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16802 = 10'hd4 == r_count_22_io_out ? io_r_212_b : _GEN_16801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16803 = 10'hd5 == r_count_22_io_out ? io_r_213_b : _GEN_16802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16804 = 10'hd6 == r_count_22_io_out ? io_r_214_b : _GEN_16803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16805 = 10'hd7 == r_count_22_io_out ? io_r_215_b : _GEN_16804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16806 = 10'hd8 == r_count_22_io_out ? io_r_216_b : _GEN_16805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16807 = 10'hd9 == r_count_22_io_out ? io_r_217_b : _GEN_16806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16808 = 10'hda == r_count_22_io_out ? io_r_218_b : _GEN_16807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16809 = 10'hdb == r_count_22_io_out ? io_r_219_b : _GEN_16808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16810 = 10'hdc == r_count_22_io_out ? io_r_220_b : _GEN_16809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16811 = 10'hdd == r_count_22_io_out ? io_r_221_b : _GEN_16810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16812 = 10'hde == r_count_22_io_out ? io_r_222_b : _GEN_16811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16813 = 10'hdf == r_count_22_io_out ? io_r_223_b : _GEN_16812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16814 = 10'he0 == r_count_22_io_out ? io_r_224_b : _GEN_16813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16815 = 10'he1 == r_count_22_io_out ? io_r_225_b : _GEN_16814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16816 = 10'he2 == r_count_22_io_out ? io_r_226_b : _GEN_16815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16817 = 10'he3 == r_count_22_io_out ? io_r_227_b : _GEN_16816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16818 = 10'he4 == r_count_22_io_out ? io_r_228_b : _GEN_16817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16819 = 10'he5 == r_count_22_io_out ? io_r_229_b : _GEN_16818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16820 = 10'he6 == r_count_22_io_out ? io_r_230_b : _GEN_16819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16821 = 10'he7 == r_count_22_io_out ? io_r_231_b : _GEN_16820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16822 = 10'he8 == r_count_22_io_out ? io_r_232_b : _GEN_16821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16823 = 10'he9 == r_count_22_io_out ? io_r_233_b : _GEN_16822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16824 = 10'hea == r_count_22_io_out ? io_r_234_b : _GEN_16823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16825 = 10'heb == r_count_22_io_out ? io_r_235_b : _GEN_16824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16826 = 10'hec == r_count_22_io_out ? io_r_236_b : _GEN_16825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16827 = 10'hed == r_count_22_io_out ? io_r_237_b : _GEN_16826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16828 = 10'hee == r_count_22_io_out ? io_r_238_b : _GEN_16827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16829 = 10'hef == r_count_22_io_out ? io_r_239_b : _GEN_16828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16830 = 10'hf0 == r_count_22_io_out ? io_r_240_b : _GEN_16829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16831 = 10'hf1 == r_count_22_io_out ? io_r_241_b : _GEN_16830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16832 = 10'hf2 == r_count_22_io_out ? io_r_242_b : _GEN_16831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16833 = 10'hf3 == r_count_22_io_out ? io_r_243_b : _GEN_16832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16834 = 10'hf4 == r_count_22_io_out ? io_r_244_b : _GEN_16833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16835 = 10'hf5 == r_count_22_io_out ? io_r_245_b : _GEN_16834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16836 = 10'hf6 == r_count_22_io_out ? io_r_246_b : _GEN_16835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16837 = 10'hf7 == r_count_22_io_out ? io_r_247_b : _GEN_16836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16838 = 10'hf8 == r_count_22_io_out ? io_r_248_b : _GEN_16837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16839 = 10'hf9 == r_count_22_io_out ? io_r_249_b : _GEN_16838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16840 = 10'hfa == r_count_22_io_out ? io_r_250_b : _GEN_16839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16841 = 10'hfb == r_count_22_io_out ? io_r_251_b : _GEN_16840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16842 = 10'hfc == r_count_22_io_out ? io_r_252_b : _GEN_16841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16843 = 10'hfd == r_count_22_io_out ? io_r_253_b : _GEN_16842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16844 = 10'hfe == r_count_22_io_out ? io_r_254_b : _GEN_16843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16845 = 10'hff == r_count_22_io_out ? io_r_255_b : _GEN_16844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16846 = 10'h100 == r_count_22_io_out ? io_r_256_b : _GEN_16845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16847 = 10'h101 == r_count_22_io_out ? io_r_257_b : _GEN_16846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16848 = 10'h102 == r_count_22_io_out ? io_r_258_b : _GEN_16847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16849 = 10'h103 == r_count_22_io_out ? io_r_259_b : _GEN_16848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16850 = 10'h104 == r_count_22_io_out ? io_r_260_b : _GEN_16849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16851 = 10'h105 == r_count_22_io_out ? io_r_261_b : _GEN_16850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16852 = 10'h106 == r_count_22_io_out ? io_r_262_b : _GEN_16851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16853 = 10'h107 == r_count_22_io_out ? io_r_263_b : _GEN_16852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16854 = 10'h108 == r_count_22_io_out ? io_r_264_b : _GEN_16853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16855 = 10'h109 == r_count_22_io_out ? io_r_265_b : _GEN_16854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16856 = 10'h10a == r_count_22_io_out ? io_r_266_b : _GEN_16855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16857 = 10'h10b == r_count_22_io_out ? io_r_267_b : _GEN_16856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16858 = 10'h10c == r_count_22_io_out ? io_r_268_b : _GEN_16857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16859 = 10'h10d == r_count_22_io_out ? io_r_269_b : _GEN_16858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16860 = 10'h10e == r_count_22_io_out ? io_r_270_b : _GEN_16859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16861 = 10'h10f == r_count_22_io_out ? io_r_271_b : _GEN_16860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16862 = 10'h110 == r_count_22_io_out ? io_r_272_b : _GEN_16861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16863 = 10'h111 == r_count_22_io_out ? io_r_273_b : _GEN_16862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16864 = 10'h112 == r_count_22_io_out ? io_r_274_b : _GEN_16863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16865 = 10'h113 == r_count_22_io_out ? io_r_275_b : _GEN_16864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16866 = 10'h114 == r_count_22_io_out ? io_r_276_b : _GEN_16865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16867 = 10'h115 == r_count_22_io_out ? io_r_277_b : _GEN_16866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16868 = 10'h116 == r_count_22_io_out ? io_r_278_b : _GEN_16867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16869 = 10'h117 == r_count_22_io_out ? io_r_279_b : _GEN_16868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16870 = 10'h118 == r_count_22_io_out ? io_r_280_b : _GEN_16869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16871 = 10'h119 == r_count_22_io_out ? io_r_281_b : _GEN_16870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16872 = 10'h11a == r_count_22_io_out ? io_r_282_b : _GEN_16871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16873 = 10'h11b == r_count_22_io_out ? io_r_283_b : _GEN_16872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16874 = 10'h11c == r_count_22_io_out ? io_r_284_b : _GEN_16873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16875 = 10'h11d == r_count_22_io_out ? io_r_285_b : _GEN_16874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16876 = 10'h11e == r_count_22_io_out ? io_r_286_b : _GEN_16875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16877 = 10'h11f == r_count_22_io_out ? io_r_287_b : _GEN_16876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16878 = 10'h120 == r_count_22_io_out ? io_r_288_b : _GEN_16877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16879 = 10'h121 == r_count_22_io_out ? io_r_289_b : _GEN_16878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16880 = 10'h122 == r_count_22_io_out ? io_r_290_b : _GEN_16879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16881 = 10'h123 == r_count_22_io_out ? io_r_291_b : _GEN_16880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16882 = 10'h124 == r_count_22_io_out ? io_r_292_b : _GEN_16881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16883 = 10'h125 == r_count_22_io_out ? io_r_293_b : _GEN_16882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16884 = 10'h126 == r_count_22_io_out ? io_r_294_b : _GEN_16883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16885 = 10'h127 == r_count_22_io_out ? io_r_295_b : _GEN_16884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16886 = 10'h128 == r_count_22_io_out ? io_r_296_b : _GEN_16885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16887 = 10'h129 == r_count_22_io_out ? io_r_297_b : _GEN_16886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16888 = 10'h12a == r_count_22_io_out ? io_r_298_b : _GEN_16887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16889 = 10'h12b == r_count_22_io_out ? io_r_299_b : _GEN_16888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16890 = 10'h12c == r_count_22_io_out ? io_r_300_b : _GEN_16889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16891 = 10'h12d == r_count_22_io_out ? io_r_301_b : _GEN_16890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16892 = 10'h12e == r_count_22_io_out ? io_r_302_b : _GEN_16891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16893 = 10'h12f == r_count_22_io_out ? io_r_303_b : _GEN_16892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16894 = 10'h130 == r_count_22_io_out ? io_r_304_b : _GEN_16893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16895 = 10'h131 == r_count_22_io_out ? io_r_305_b : _GEN_16894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16896 = 10'h132 == r_count_22_io_out ? io_r_306_b : _GEN_16895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16897 = 10'h133 == r_count_22_io_out ? io_r_307_b : _GEN_16896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16898 = 10'h134 == r_count_22_io_out ? io_r_308_b : _GEN_16897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16899 = 10'h135 == r_count_22_io_out ? io_r_309_b : _GEN_16898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16900 = 10'h136 == r_count_22_io_out ? io_r_310_b : _GEN_16899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16901 = 10'h137 == r_count_22_io_out ? io_r_311_b : _GEN_16900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16902 = 10'h138 == r_count_22_io_out ? io_r_312_b : _GEN_16901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16903 = 10'h139 == r_count_22_io_out ? io_r_313_b : _GEN_16902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16904 = 10'h13a == r_count_22_io_out ? io_r_314_b : _GEN_16903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16905 = 10'h13b == r_count_22_io_out ? io_r_315_b : _GEN_16904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16906 = 10'h13c == r_count_22_io_out ? io_r_316_b : _GEN_16905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16907 = 10'h13d == r_count_22_io_out ? io_r_317_b : _GEN_16906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16908 = 10'h13e == r_count_22_io_out ? io_r_318_b : _GEN_16907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16909 = 10'h13f == r_count_22_io_out ? io_r_319_b : _GEN_16908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16910 = 10'h140 == r_count_22_io_out ? io_r_320_b : _GEN_16909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16911 = 10'h141 == r_count_22_io_out ? io_r_321_b : _GEN_16910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16912 = 10'h142 == r_count_22_io_out ? io_r_322_b : _GEN_16911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16913 = 10'h143 == r_count_22_io_out ? io_r_323_b : _GEN_16912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16914 = 10'h144 == r_count_22_io_out ? io_r_324_b : _GEN_16913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16915 = 10'h145 == r_count_22_io_out ? io_r_325_b : _GEN_16914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16916 = 10'h146 == r_count_22_io_out ? io_r_326_b : _GEN_16915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16917 = 10'h147 == r_count_22_io_out ? io_r_327_b : _GEN_16916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16918 = 10'h148 == r_count_22_io_out ? io_r_328_b : _GEN_16917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16919 = 10'h149 == r_count_22_io_out ? io_r_329_b : _GEN_16918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16920 = 10'h14a == r_count_22_io_out ? io_r_330_b : _GEN_16919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16921 = 10'h14b == r_count_22_io_out ? io_r_331_b : _GEN_16920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16922 = 10'h14c == r_count_22_io_out ? io_r_332_b : _GEN_16921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16923 = 10'h14d == r_count_22_io_out ? io_r_333_b : _GEN_16922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16924 = 10'h14e == r_count_22_io_out ? io_r_334_b : _GEN_16923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16925 = 10'h14f == r_count_22_io_out ? io_r_335_b : _GEN_16924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16926 = 10'h150 == r_count_22_io_out ? io_r_336_b : _GEN_16925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16927 = 10'h151 == r_count_22_io_out ? io_r_337_b : _GEN_16926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16928 = 10'h152 == r_count_22_io_out ? io_r_338_b : _GEN_16927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16929 = 10'h153 == r_count_22_io_out ? io_r_339_b : _GEN_16928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16930 = 10'h154 == r_count_22_io_out ? io_r_340_b : _GEN_16929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16931 = 10'h155 == r_count_22_io_out ? io_r_341_b : _GEN_16930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16932 = 10'h156 == r_count_22_io_out ? io_r_342_b : _GEN_16931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16933 = 10'h157 == r_count_22_io_out ? io_r_343_b : _GEN_16932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16934 = 10'h158 == r_count_22_io_out ? io_r_344_b : _GEN_16933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16935 = 10'h159 == r_count_22_io_out ? io_r_345_b : _GEN_16934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16936 = 10'h15a == r_count_22_io_out ? io_r_346_b : _GEN_16935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16937 = 10'h15b == r_count_22_io_out ? io_r_347_b : _GEN_16936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16938 = 10'h15c == r_count_22_io_out ? io_r_348_b : _GEN_16937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16939 = 10'h15d == r_count_22_io_out ? io_r_349_b : _GEN_16938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16940 = 10'h15e == r_count_22_io_out ? io_r_350_b : _GEN_16939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16941 = 10'h15f == r_count_22_io_out ? io_r_351_b : _GEN_16940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16942 = 10'h160 == r_count_22_io_out ? io_r_352_b : _GEN_16941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16943 = 10'h161 == r_count_22_io_out ? io_r_353_b : _GEN_16942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16944 = 10'h162 == r_count_22_io_out ? io_r_354_b : _GEN_16943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16945 = 10'h163 == r_count_22_io_out ? io_r_355_b : _GEN_16944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16946 = 10'h164 == r_count_22_io_out ? io_r_356_b : _GEN_16945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16947 = 10'h165 == r_count_22_io_out ? io_r_357_b : _GEN_16946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16948 = 10'h166 == r_count_22_io_out ? io_r_358_b : _GEN_16947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16949 = 10'h167 == r_count_22_io_out ? io_r_359_b : _GEN_16948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16950 = 10'h168 == r_count_22_io_out ? io_r_360_b : _GEN_16949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16951 = 10'h169 == r_count_22_io_out ? io_r_361_b : _GEN_16950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16952 = 10'h16a == r_count_22_io_out ? io_r_362_b : _GEN_16951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16953 = 10'h16b == r_count_22_io_out ? io_r_363_b : _GEN_16952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16954 = 10'h16c == r_count_22_io_out ? io_r_364_b : _GEN_16953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16955 = 10'h16d == r_count_22_io_out ? io_r_365_b : _GEN_16954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16956 = 10'h16e == r_count_22_io_out ? io_r_366_b : _GEN_16955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16957 = 10'h16f == r_count_22_io_out ? io_r_367_b : _GEN_16956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16958 = 10'h170 == r_count_22_io_out ? io_r_368_b : _GEN_16957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16959 = 10'h171 == r_count_22_io_out ? io_r_369_b : _GEN_16958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16960 = 10'h172 == r_count_22_io_out ? io_r_370_b : _GEN_16959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16961 = 10'h173 == r_count_22_io_out ? io_r_371_b : _GEN_16960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16962 = 10'h174 == r_count_22_io_out ? io_r_372_b : _GEN_16961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16963 = 10'h175 == r_count_22_io_out ? io_r_373_b : _GEN_16962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16964 = 10'h176 == r_count_22_io_out ? io_r_374_b : _GEN_16963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16965 = 10'h177 == r_count_22_io_out ? io_r_375_b : _GEN_16964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16966 = 10'h178 == r_count_22_io_out ? io_r_376_b : _GEN_16965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16967 = 10'h179 == r_count_22_io_out ? io_r_377_b : _GEN_16966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16968 = 10'h17a == r_count_22_io_out ? io_r_378_b : _GEN_16967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16969 = 10'h17b == r_count_22_io_out ? io_r_379_b : _GEN_16968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16970 = 10'h17c == r_count_22_io_out ? io_r_380_b : _GEN_16969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16971 = 10'h17d == r_count_22_io_out ? io_r_381_b : _GEN_16970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16972 = 10'h17e == r_count_22_io_out ? io_r_382_b : _GEN_16971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16973 = 10'h17f == r_count_22_io_out ? io_r_383_b : _GEN_16972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16974 = 10'h180 == r_count_22_io_out ? io_r_384_b : _GEN_16973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16975 = 10'h181 == r_count_22_io_out ? io_r_385_b : _GEN_16974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16976 = 10'h182 == r_count_22_io_out ? io_r_386_b : _GEN_16975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16977 = 10'h183 == r_count_22_io_out ? io_r_387_b : _GEN_16976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16978 = 10'h184 == r_count_22_io_out ? io_r_388_b : _GEN_16977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16979 = 10'h185 == r_count_22_io_out ? io_r_389_b : _GEN_16978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16980 = 10'h186 == r_count_22_io_out ? io_r_390_b : _GEN_16979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16981 = 10'h187 == r_count_22_io_out ? io_r_391_b : _GEN_16980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16982 = 10'h188 == r_count_22_io_out ? io_r_392_b : _GEN_16981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16983 = 10'h189 == r_count_22_io_out ? io_r_393_b : _GEN_16982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16984 = 10'h18a == r_count_22_io_out ? io_r_394_b : _GEN_16983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16985 = 10'h18b == r_count_22_io_out ? io_r_395_b : _GEN_16984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16986 = 10'h18c == r_count_22_io_out ? io_r_396_b : _GEN_16985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16987 = 10'h18d == r_count_22_io_out ? io_r_397_b : _GEN_16986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16988 = 10'h18e == r_count_22_io_out ? io_r_398_b : _GEN_16987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16989 = 10'h18f == r_count_22_io_out ? io_r_399_b : _GEN_16988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16990 = 10'h190 == r_count_22_io_out ? io_r_400_b : _GEN_16989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16991 = 10'h191 == r_count_22_io_out ? io_r_401_b : _GEN_16990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16992 = 10'h192 == r_count_22_io_out ? io_r_402_b : _GEN_16991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16993 = 10'h193 == r_count_22_io_out ? io_r_403_b : _GEN_16992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16994 = 10'h194 == r_count_22_io_out ? io_r_404_b : _GEN_16993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16995 = 10'h195 == r_count_22_io_out ? io_r_405_b : _GEN_16994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16996 = 10'h196 == r_count_22_io_out ? io_r_406_b : _GEN_16995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16997 = 10'h197 == r_count_22_io_out ? io_r_407_b : _GEN_16996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16998 = 10'h198 == r_count_22_io_out ? io_r_408_b : _GEN_16997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16999 = 10'h199 == r_count_22_io_out ? io_r_409_b : _GEN_16998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17000 = 10'h19a == r_count_22_io_out ? io_r_410_b : _GEN_16999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17001 = 10'h19b == r_count_22_io_out ? io_r_411_b : _GEN_17000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17002 = 10'h19c == r_count_22_io_out ? io_r_412_b : _GEN_17001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17003 = 10'h19d == r_count_22_io_out ? io_r_413_b : _GEN_17002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17004 = 10'h19e == r_count_22_io_out ? io_r_414_b : _GEN_17003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17005 = 10'h19f == r_count_22_io_out ? io_r_415_b : _GEN_17004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17006 = 10'h1a0 == r_count_22_io_out ? io_r_416_b : _GEN_17005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17007 = 10'h1a1 == r_count_22_io_out ? io_r_417_b : _GEN_17006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17008 = 10'h1a2 == r_count_22_io_out ? io_r_418_b : _GEN_17007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17009 = 10'h1a3 == r_count_22_io_out ? io_r_419_b : _GEN_17008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17010 = 10'h1a4 == r_count_22_io_out ? io_r_420_b : _GEN_17009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17011 = 10'h1a5 == r_count_22_io_out ? io_r_421_b : _GEN_17010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17012 = 10'h1a6 == r_count_22_io_out ? io_r_422_b : _GEN_17011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17013 = 10'h1a7 == r_count_22_io_out ? io_r_423_b : _GEN_17012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17014 = 10'h1a8 == r_count_22_io_out ? io_r_424_b : _GEN_17013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17015 = 10'h1a9 == r_count_22_io_out ? io_r_425_b : _GEN_17014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17016 = 10'h1aa == r_count_22_io_out ? io_r_426_b : _GEN_17015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17017 = 10'h1ab == r_count_22_io_out ? io_r_427_b : _GEN_17016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17018 = 10'h1ac == r_count_22_io_out ? io_r_428_b : _GEN_17017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17019 = 10'h1ad == r_count_22_io_out ? io_r_429_b : _GEN_17018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17020 = 10'h1ae == r_count_22_io_out ? io_r_430_b : _GEN_17019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17021 = 10'h1af == r_count_22_io_out ? io_r_431_b : _GEN_17020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17022 = 10'h1b0 == r_count_22_io_out ? io_r_432_b : _GEN_17021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17023 = 10'h1b1 == r_count_22_io_out ? io_r_433_b : _GEN_17022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17024 = 10'h1b2 == r_count_22_io_out ? io_r_434_b : _GEN_17023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17025 = 10'h1b3 == r_count_22_io_out ? io_r_435_b : _GEN_17024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17026 = 10'h1b4 == r_count_22_io_out ? io_r_436_b : _GEN_17025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17027 = 10'h1b5 == r_count_22_io_out ? io_r_437_b : _GEN_17026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17028 = 10'h1b6 == r_count_22_io_out ? io_r_438_b : _GEN_17027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17029 = 10'h1b7 == r_count_22_io_out ? io_r_439_b : _GEN_17028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17030 = 10'h1b8 == r_count_22_io_out ? io_r_440_b : _GEN_17029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17031 = 10'h1b9 == r_count_22_io_out ? io_r_441_b : _GEN_17030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17032 = 10'h1ba == r_count_22_io_out ? io_r_442_b : _GEN_17031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17033 = 10'h1bb == r_count_22_io_out ? io_r_443_b : _GEN_17032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17034 = 10'h1bc == r_count_22_io_out ? io_r_444_b : _GEN_17033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17035 = 10'h1bd == r_count_22_io_out ? io_r_445_b : _GEN_17034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17036 = 10'h1be == r_count_22_io_out ? io_r_446_b : _GEN_17035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17037 = 10'h1bf == r_count_22_io_out ? io_r_447_b : _GEN_17036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17038 = 10'h1c0 == r_count_22_io_out ? io_r_448_b : _GEN_17037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17039 = 10'h1c1 == r_count_22_io_out ? io_r_449_b : _GEN_17038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17040 = 10'h1c2 == r_count_22_io_out ? io_r_450_b : _GEN_17039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17041 = 10'h1c3 == r_count_22_io_out ? io_r_451_b : _GEN_17040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17042 = 10'h1c4 == r_count_22_io_out ? io_r_452_b : _GEN_17041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17043 = 10'h1c5 == r_count_22_io_out ? io_r_453_b : _GEN_17042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17044 = 10'h1c6 == r_count_22_io_out ? io_r_454_b : _GEN_17043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17045 = 10'h1c7 == r_count_22_io_out ? io_r_455_b : _GEN_17044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17046 = 10'h1c8 == r_count_22_io_out ? io_r_456_b : _GEN_17045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17047 = 10'h1c9 == r_count_22_io_out ? io_r_457_b : _GEN_17046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17048 = 10'h1ca == r_count_22_io_out ? io_r_458_b : _GEN_17047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17049 = 10'h1cb == r_count_22_io_out ? io_r_459_b : _GEN_17048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17050 = 10'h1cc == r_count_22_io_out ? io_r_460_b : _GEN_17049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17051 = 10'h1cd == r_count_22_io_out ? io_r_461_b : _GEN_17050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17052 = 10'h1ce == r_count_22_io_out ? io_r_462_b : _GEN_17051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17053 = 10'h1cf == r_count_22_io_out ? io_r_463_b : _GEN_17052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17054 = 10'h1d0 == r_count_22_io_out ? io_r_464_b : _GEN_17053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17055 = 10'h1d1 == r_count_22_io_out ? io_r_465_b : _GEN_17054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17056 = 10'h1d2 == r_count_22_io_out ? io_r_466_b : _GEN_17055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17057 = 10'h1d3 == r_count_22_io_out ? io_r_467_b : _GEN_17056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17058 = 10'h1d4 == r_count_22_io_out ? io_r_468_b : _GEN_17057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17059 = 10'h1d5 == r_count_22_io_out ? io_r_469_b : _GEN_17058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17060 = 10'h1d6 == r_count_22_io_out ? io_r_470_b : _GEN_17059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17061 = 10'h1d7 == r_count_22_io_out ? io_r_471_b : _GEN_17060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17062 = 10'h1d8 == r_count_22_io_out ? io_r_472_b : _GEN_17061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17063 = 10'h1d9 == r_count_22_io_out ? io_r_473_b : _GEN_17062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17064 = 10'h1da == r_count_22_io_out ? io_r_474_b : _GEN_17063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17065 = 10'h1db == r_count_22_io_out ? io_r_475_b : _GEN_17064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17066 = 10'h1dc == r_count_22_io_out ? io_r_476_b : _GEN_17065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17067 = 10'h1dd == r_count_22_io_out ? io_r_477_b : _GEN_17066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17068 = 10'h1de == r_count_22_io_out ? io_r_478_b : _GEN_17067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17069 = 10'h1df == r_count_22_io_out ? io_r_479_b : _GEN_17068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17070 = 10'h1e0 == r_count_22_io_out ? io_r_480_b : _GEN_17069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17071 = 10'h1e1 == r_count_22_io_out ? io_r_481_b : _GEN_17070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17072 = 10'h1e2 == r_count_22_io_out ? io_r_482_b : _GEN_17071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17073 = 10'h1e3 == r_count_22_io_out ? io_r_483_b : _GEN_17072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17074 = 10'h1e4 == r_count_22_io_out ? io_r_484_b : _GEN_17073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17075 = 10'h1e5 == r_count_22_io_out ? io_r_485_b : _GEN_17074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17076 = 10'h1e6 == r_count_22_io_out ? io_r_486_b : _GEN_17075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17077 = 10'h1e7 == r_count_22_io_out ? io_r_487_b : _GEN_17076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17078 = 10'h1e8 == r_count_22_io_out ? io_r_488_b : _GEN_17077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17079 = 10'h1e9 == r_count_22_io_out ? io_r_489_b : _GEN_17078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17080 = 10'h1ea == r_count_22_io_out ? io_r_490_b : _GEN_17079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17081 = 10'h1eb == r_count_22_io_out ? io_r_491_b : _GEN_17080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17082 = 10'h1ec == r_count_22_io_out ? io_r_492_b : _GEN_17081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17083 = 10'h1ed == r_count_22_io_out ? io_r_493_b : _GEN_17082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17084 = 10'h1ee == r_count_22_io_out ? io_r_494_b : _GEN_17083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17085 = 10'h1ef == r_count_22_io_out ? io_r_495_b : _GEN_17084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17086 = 10'h1f0 == r_count_22_io_out ? io_r_496_b : _GEN_17085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17087 = 10'h1f1 == r_count_22_io_out ? io_r_497_b : _GEN_17086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17088 = 10'h1f2 == r_count_22_io_out ? io_r_498_b : _GEN_17087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17089 = 10'h1f3 == r_count_22_io_out ? io_r_499_b : _GEN_17088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17090 = 10'h1f4 == r_count_22_io_out ? io_r_500_b : _GEN_17089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17091 = 10'h1f5 == r_count_22_io_out ? io_r_501_b : _GEN_17090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17092 = 10'h1f6 == r_count_22_io_out ? io_r_502_b : _GEN_17091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17093 = 10'h1f7 == r_count_22_io_out ? io_r_503_b : _GEN_17092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17094 = 10'h1f8 == r_count_22_io_out ? io_r_504_b : _GEN_17093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17095 = 10'h1f9 == r_count_22_io_out ? io_r_505_b : _GEN_17094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17096 = 10'h1fa == r_count_22_io_out ? io_r_506_b : _GEN_17095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17097 = 10'h1fb == r_count_22_io_out ? io_r_507_b : _GEN_17096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17098 = 10'h1fc == r_count_22_io_out ? io_r_508_b : _GEN_17097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17099 = 10'h1fd == r_count_22_io_out ? io_r_509_b : _GEN_17098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17100 = 10'h1fe == r_count_22_io_out ? io_r_510_b : _GEN_17099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17101 = 10'h1ff == r_count_22_io_out ? io_r_511_b : _GEN_17100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17102 = 10'h200 == r_count_22_io_out ? io_r_512_b : _GEN_17101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17103 = 10'h201 == r_count_22_io_out ? io_r_513_b : _GEN_17102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17104 = 10'h202 == r_count_22_io_out ? io_r_514_b : _GEN_17103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17105 = 10'h203 == r_count_22_io_out ? io_r_515_b : _GEN_17104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17106 = 10'h204 == r_count_22_io_out ? io_r_516_b : _GEN_17105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17107 = 10'h205 == r_count_22_io_out ? io_r_517_b : _GEN_17106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17108 = 10'h206 == r_count_22_io_out ? io_r_518_b : _GEN_17107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17109 = 10'h207 == r_count_22_io_out ? io_r_519_b : _GEN_17108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17110 = 10'h208 == r_count_22_io_out ? io_r_520_b : _GEN_17109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17111 = 10'h209 == r_count_22_io_out ? io_r_521_b : _GEN_17110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17112 = 10'h20a == r_count_22_io_out ? io_r_522_b : _GEN_17111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17113 = 10'h20b == r_count_22_io_out ? io_r_523_b : _GEN_17112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17114 = 10'h20c == r_count_22_io_out ? io_r_524_b : _GEN_17113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17115 = 10'h20d == r_count_22_io_out ? io_r_525_b : _GEN_17114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17116 = 10'h20e == r_count_22_io_out ? io_r_526_b : _GEN_17115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17117 = 10'h20f == r_count_22_io_out ? io_r_527_b : _GEN_17116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17118 = 10'h210 == r_count_22_io_out ? io_r_528_b : _GEN_17117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17119 = 10'h211 == r_count_22_io_out ? io_r_529_b : _GEN_17118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17120 = 10'h212 == r_count_22_io_out ? io_r_530_b : _GEN_17119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17121 = 10'h213 == r_count_22_io_out ? io_r_531_b : _GEN_17120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17122 = 10'h214 == r_count_22_io_out ? io_r_532_b : _GEN_17121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17123 = 10'h215 == r_count_22_io_out ? io_r_533_b : _GEN_17122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17124 = 10'h216 == r_count_22_io_out ? io_r_534_b : _GEN_17123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17125 = 10'h217 == r_count_22_io_out ? io_r_535_b : _GEN_17124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17126 = 10'h218 == r_count_22_io_out ? io_r_536_b : _GEN_17125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17127 = 10'h219 == r_count_22_io_out ? io_r_537_b : _GEN_17126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17128 = 10'h21a == r_count_22_io_out ? io_r_538_b : _GEN_17127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17129 = 10'h21b == r_count_22_io_out ? io_r_539_b : _GEN_17128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17130 = 10'h21c == r_count_22_io_out ? io_r_540_b : _GEN_17129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17131 = 10'h21d == r_count_22_io_out ? io_r_541_b : _GEN_17130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17132 = 10'h21e == r_count_22_io_out ? io_r_542_b : _GEN_17131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17133 = 10'h21f == r_count_22_io_out ? io_r_543_b : _GEN_17132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17134 = 10'h220 == r_count_22_io_out ? io_r_544_b : _GEN_17133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17135 = 10'h221 == r_count_22_io_out ? io_r_545_b : _GEN_17134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17136 = 10'h222 == r_count_22_io_out ? io_r_546_b : _GEN_17135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17137 = 10'h223 == r_count_22_io_out ? io_r_547_b : _GEN_17136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17138 = 10'h224 == r_count_22_io_out ? io_r_548_b : _GEN_17137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17139 = 10'h225 == r_count_22_io_out ? io_r_549_b : _GEN_17138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17140 = 10'h226 == r_count_22_io_out ? io_r_550_b : _GEN_17139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17141 = 10'h227 == r_count_22_io_out ? io_r_551_b : _GEN_17140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17142 = 10'h228 == r_count_22_io_out ? io_r_552_b : _GEN_17141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17143 = 10'h229 == r_count_22_io_out ? io_r_553_b : _GEN_17142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17144 = 10'h22a == r_count_22_io_out ? io_r_554_b : _GEN_17143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17145 = 10'h22b == r_count_22_io_out ? io_r_555_b : _GEN_17144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17146 = 10'h22c == r_count_22_io_out ? io_r_556_b : _GEN_17145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17147 = 10'h22d == r_count_22_io_out ? io_r_557_b : _GEN_17146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17148 = 10'h22e == r_count_22_io_out ? io_r_558_b : _GEN_17147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17149 = 10'h22f == r_count_22_io_out ? io_r_559_b : _GEN_17148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17150 = 10'h230 == r_count_22_io_out ? io_r_560_b : _GEN_17149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17151 = 10'h231 == r_count_22_io_out ? io_r_561_b : _GEN_17150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17152 = 10'h232 == r_count_22_io_out ? io_r_562_b : _GEN_17151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17153 = 10'h233 == r_count_22_io_out ? io_r_563_b : _GEN_17152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17154 = 10'h234 == r_count_22_io_out ? io_r_564_b : _GEN_17153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17155 = 10'h235 == r_count_22_io_out ? io_r_565_b : _GEN_17154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17156 = 10'h236 == r_count_22_io_out ? io_r_566_b : _GEN_17155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17157 = 10'h237 == r_count_22_io_out ? io_r_567_b : _GEN_17156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17158 = 10'h238 == r_count_22_io_out ? io_r_568_b : _GEN_17157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17159 = 10'h239 == r_count_22_io_out ? io_r_569_b : _GEN_17158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17160 = 10'h23a == r_count_22_io_out ? io_r_570_b : _GEN_17159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17161 = 10'h23b == r_count_22_io_out ? io_r_571_b : _GEN_17160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17162 = 10'h23c == r_count_22_io_out ? io_r_572_b : _GEN_17161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17163 = 10'h23d == r_count_22_io_out ? io_r_573_b : _GEN_17162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17164 = 10'h23e == r_count_22_io_out ? io_r_574_b : _GEN_17163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17165 = 10'h23f == r_count_22_io_out ? io_r_575_b : _GEN_17164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17166 = 10'h240 == r_count_22_io_out ? io_r_576_b : _GEN_17165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17167 = 10'h241 == r_count_22_io_out ? io_r_577_b : _GEN_17166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17168 = 10'h242 == r_count_22_io_out ? io_r_578_b : _GEN_17167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17169 = 10'h243 == r_count_22_io_out ? io_r_579_b : _GEN_17168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17170 = 10'h244 == r_count_22_io_out ? io_r_580_b : _GEN_17169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17171 = 10'h245 == r_count_22_io_out ? io_r_581_b : _GEN_17170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17172 = 10'h246 == r_count_22_io_out ? io_r_582_b : _GEN_17171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17173 = 10'h247 == r_count_22_io_out ? io_r_583_b : _GEN_17172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17174 = 10'h248 == r_count_22_io_out ? io_r_584_b : _GEN_17173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17175 = 10'h249 == r_count_22_io_out ? io_r_585_b : _GEN_17174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17176 = 10'h24a == r_count_22_io_out ? io_r_586_b : _GEN_17175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17177 = 10'h24b == r_count_22_io_out ? io_r_587_b : _GEN_17176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17178 = 10'h24c == r_count_22_io_out ? io_r_588_b : _GEN_17177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17179 = 10'h24d == r_count_22_io_out ? io_r_589_b : _GEN_17178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17180 = 10'h24e == r_count_22_io_out ? io_r_590_b : _GEN_17179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17181 = 10'h24f == r_count_22_io_out ? io_r_591_b : _GEN_17180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17182 = 10'h250 == r_count_22_io_out ? io_r_592_b : _GEN_17181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17183 = 10'h251 == r_count_22_io_out ? io_r_593_b : _GEN_17182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17184 = 10'h252 == r_count_22_io_out ? io_r_594_b : _GEN_17183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17185 = 10'h253 == r_count_22_io_out ? io_r_595_b : _GEN_17184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17186 = 10'h254 == r_count_22_io_out ? io_r_596_b : _GEN_17185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17187 = 10'h255 == r_count_22_io_out ? io_r_597_b : _GEN_17186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17188 = 10'h256 == r_count_22_io_out ? io_r_598_b : _GEN_17187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17189 = 10'h257 == r_count_22_io_out ? io_r_599_b : _GEN_17188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17190 = 10'h258 == r_count_22_io_out ? io_r_600_b : _GEN_17189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17191 = 10'h259 == r_count_22_io_out ? io_r_601_b : _GEN_17190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17192 = 10'h25a == r_count_22_io_out ? io_r_602_b : _GEN_17191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17193 = 10'h25b == r_count_22_io_out ? io_r_603_b : _GEN_17192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17194 = 10'h25c == r_count_22_io_out ? io_r_604_b : _GEN_17193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17195 = 10'h25d == r_count_22_io_out ? io_r_605_b : _GEN_17194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17196 = 10'h25e == r_count_22_io_out ? io_r_606_b : _GEN_17195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17197 = 10'h25f == r_count_22_io_out ? io_r_607_b : _GEN_17196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17198 = 10'h260 == r_count_22_io_out ? io_r_608_b : _GEN_17197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17199 = 10'h261 == r_count_22_io_out ? io_r_609_b : _GEN_17198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17200 = 10'h262 == r_count_22_io_out ? io_r_610_b : _GEN_17199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17201 = 10'h263 == r_count_22_io_out ? io_r_611_b : _GEN_17200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17202 = 10'h264 == r_count_22_io_out ? io_r_612_b : _GEN_17201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17203 = 10'h265 == r_count_22_io_out ? io_r_613_b : _GEN_17202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17204 = 10'h266 == r_count_22_io_out ? io_r_614_b : _GEN_17203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17205 = 10'h267 == r_count_22_io_out ? io_r_615_b : _GEN_17204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17206 = 10'h268 == r_count_22_io_out ? io_r_616_b : _GEN_17205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17207 = 10'h269 == r_count_22_io_out ? io_r_617_b : _GEN_17206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17208 = 10'h26a == r_count_22_io_out ? io_r_618_b : _GEN_17207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17209 = 10'h26b == r_count_22_io_out ? io_r_619_b : _GEN_17208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17210 = 10'h26c == r_count_22_io_out ? io_r_620_b : _GEN_17209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17211 = 10'h26d == r_count_22_io_out ? io_r_621_b : _GEN_17210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17212 = 10'h26e == r_count_22_io_out ? io_r_622_b : _GEN_17211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17213 = 10'h26f == r_count_22_io_out ? io_r_623_b : _GEN_17212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17214 = 10'h270 == r_count_22_io_out ? io_r_624_b : _GEN_17213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17215 = 10'h271 == r_count_22_io_out ? io_r_625_b : _GEN_17214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17216 = 10'h272 == r_count_22_io_out ? io_r_626_b : _GEN_17215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17217 = 10'h273 == r_count_22_io_out ? io_r_627_b : _GEN_17216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17218 = 10'h274 == r_count_22_io_out ? io_r_628_b : _GEN_17217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17219 = 10'h275 == r_count_22_io_out ? io_r_629_b : _GEN_17218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17220 = 10'h276 == r_count_22_io_out ? io_r_630_b : _GEN_17219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17221 = 10'h277 == r_count_22_io_out ? io_r_631_b : _GEN_17220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17222 = 10'h278 == r_count_22_io_out ? io_r_632_b : _GEN_17221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17223 = 10'h279 == r_count_22_io_out ? io_r_633_b : _GEN_17222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17224 = 10'h27a == r_count_22_io_out ? io_r_634_b : _GEN_17223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17225 = 10'h27b == r_count_22_io_out ? io_r_635_b : _GEN_17224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17226 = 10'h27c == r_count_22_io_out ? io_r_636_b : _GEN_17225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17227 = 10'h27d == r_count_22_io_out ? io_r_637_b : _GEN_17226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17228 = 10'h27e == r_count_22_io_out ? io_r_638_b : _GEN_17227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17229 = 10'h27f == r_count_22_io_out ? io_r_639_b : _GEN_17228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17230 = 10'h280 == r_count_22_io_out ? io_r_640_b : _GEN_17229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17231 = 10'h281 == r_count_22_io_out ? io_r_641_b : _GEN_17230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17232 = 10'h282 == r_count_22_io_out ? io_r_642_b : _GEN_17231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17233 = 10'h283 == r_count_22_io_out ? io_r_643_b : _GEN_17232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17234 = 10'h284 == r_count_22_io_out ? io_r_644_b : _GEN_17233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17235 = 10'h285 == r_count_22_io_out ? io_r_645_b : _GEN_17234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17236 = 10'h286 == r_count_22_io_out ? io_r_646_b : _GEN_17235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17237 = 10'h287 == r_count_22_io_out ? io_r_647_b : _GEN_17236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17238 = 10'h288 == r_count_22_io_out ? io_r_648_b : _GEN_17237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17239 = 10'h289 == r_count_22_io_out ? io_r_649_b : _GEN_17238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17240 = 10'h28a == r_count_22_io_out ? io_r_650_b : _GEN_17239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17241 = 10'h28b == r_count_22_io_out ? io_r_651_b : _GEN_17240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17242 = 10'h28c == r_count_22_io_out ? io_r_652_b : _GEN_17241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17243 = 10'h28d == r_count_22_io_out ? io_r_653_b : _GEN_17242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17244 = 10'h28e == r_count_22_io_out ? io_r_654_b : _GEN_17243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17245 = 10'h28f == r_count_22_io_out ? io_r_655_b : _GEN_17244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17246 = 10'h290 == r_count_22_io_out ? io_r_656_b : _GEN_17245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17247 = 10'h291 == r_count_22_io_out ? io_r_657_b : _GEN_17246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17248 = 10'h292 == r_count_22_io_out ? io_r_658_b : _GEN_17247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17249 = 10'h293 == r_count_22_io_out ? io_r_659_b : _GEN_17248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17250 = 10'h294 == r_count_22_io_out ? io_r_660_b : _GEN_17249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17251 = 10'h295 == r_count_22_io_out ? io_r_661_b : _GEN_17250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17252 = 10'h296 == r_count_22_io_out ? io_r_662_b : _GEN_17251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17253 = 10'h297 == r_count_22_io_out ? io_r_663_b : _GEN_17252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17254 = 10'h298 == r_count_22_io_out ? io_r_664_b : _GEN_17253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17255 = 10'h299 == r_count_22_io_out ? io_r_665_b : _GEN_17254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17256 = 10'h29a == r_count_22_io_out ? io_r_666_b : _GEN_17255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17257 = 10'h29b == r_count_22_io_out ? io_r_667_b : _GEN_17256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17258 = 10'h29c == r_count_22_io_out ? io_r_668_b : _GEN_17257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17259 = 10'h29d == r_count_22_io_out ? io_r_669_b : _GEN_17258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17260 = 10'h29e == r_count_22_io_out ? io_r_670_b : _GEN_17259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17261 = 10'h29f == r_count_22_io_out ? io_r_671_b : _GEN_17260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17262 = 10'h2a0 == r_count_22_io_out ? io_r_672_b : _GEN_17261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17263 = 10'h2a1 == r_count_22_io_out ? io_r_673_b : _GEN_17262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17264 = 10'h2a2 == r_count_22_io_out ? io_r_674_b : _GEN_17263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17265 = 10'h2a3 == r_count_22_io_out ? io_r_675_b : _GEN_17264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17266 = 10'h2a4 == r_count_22_io_out ? io_r_676_b : _GEN_17265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17267 = 10'h2a5 == r_count_22_io_out ? io_r_677_b : _GEN_17266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17268 = 10'h2a6 == r_count_22_io_out ? io_r_678_b : _GEN_17267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17269 = 10'h2a7 == r_count_22_io_out ? io_r_679_b : _GEN_17268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17270 = 10'h2a8 == r_count_22_io_out ? io_r_680_b : _GEN_17269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17271 = 10'h2a9 == r_count_22_io_out ? io_r_681_b : _GEN_17270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17272 = 10'h2aa == r_count_22_io_out ? io_r_682_b : _GEN_17271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17273 = 10'h2ab == r_count_22_io_out ? io_r_683_b : _GEN_17272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17274 = 10'h2ac == r_count_22_io_out ? io_r_684_b : _GEN_17273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17275 = 10'h2ad == r_count_22_io_out ? io_r_685_b : _GEN_17274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17276 = 10'h2ae == r_count_22_io_out ? io_r_686_b : _GEN_17275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17277 = 10'h2af == r_count_22_io_out ? io_r_687_b : _GEN_17276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17278 = 10'h2b0 == r_count_22_io_out ? io_r_688_b : _GEN_17277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17279 = 10'h2b1 == r_count_22_io_out ? io_r_689_b : _GEN_17278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17280 = 10'h2b2 == r_count_22_io_out ? io_r_690_b : _GEN_17279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17281 = 10'h2b3 == r_count_22_io_out ? io_r_691_b : _GEN_17280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17282 = 10'h2b4 == r_count_22_io_out ? io_r_692_b : _GEN_17281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17283 = 10'h2b5 == r_count_22_io_out ? io_r_693_b : _GEN_17282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17284 = 10'h2b6 == r_count_22_io_out ? io_r_694_b : _GEN_17283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17285 = 10'h2b7 == r_count_22_io_out ? io_r_695_b : _GEN_17284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17286 = 10'h2b8 == r_count_22_io_out ? io_r_696_b : _GEN_17285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17287 = 10'h2b9 == r_count_22_io_out ? io_r_697_b : _GEN_17286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17288 = 10'h2ba == r_count_22_io_out ? io_r_698_b : _GEN_17287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17289 = 10'h2bb == r_count_22_io_out ? io_r_699_b : _GEN_17288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17290 = 10'h2bc == r_count_22_io_out ? io_r_700_b : _GEN_17289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17291 = 10'h2bd == r_count_22_io_out ? io_r_701_b : _GEN_17290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17292 = 10'h2be == r_count_22_io_out ? io_r_702_b : _GEN_17291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17293 = 10'h2bf == r_count_22_io_out ? io_r_703_b : _GEN_17292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17294 = 10'h2c0 == r_count_22_io_out ? io_r_704_b : _GEN_17293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17295 = 10'h2c1 == r_count_22_io_out ? io_r_705_b : _GEN_17294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17296 = 10'h2c2 == r_count_22_io_out ? io_r_706_b : _GEN_17295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17297 = 10'h2c3 == r_count_22_io_out ? io_r_707_b : _GEN_17296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17298 = 10'h2c4 == r_count_22_io_out ? io_r_708_b : _GEN_17297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17299 = 10'h2c5 == r_count_22_io_out ? io_r_709_b : _GEN_17298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17300 = 10'h2c6 == r_count_22_io_out ? io_r_710_b : _GEN_17299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17301 = 10'h2c7 == r_count_22_io_out ? io_r_711_b : _GEN_17300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17302 = 10'h2c8 == r_count_22_io_out ? io_r_712_b : _GEN_17301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17303 = 10'h2c9 == r_count_22_io_out ? io_r_713_b : _GEN_17302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17304 = 10'h2ca == r_count_22_io_out ? io_r_714_b : _GEN_17303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17305 = 10'h2cb == r_count_22_io_out ? io_r_715_b : _GEN_17304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17306 = 10'h2cc == r_count_22_io_out ? io_r_716_b : _GEN_17305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17307 = 10'h2cd == r_count_22_io_out ? io_r_717_b : _GEN_17306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17308 = 10'h2ce == r_count_22_io_out ? io_r_718_b : _GEN_17307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17309 = 10'h2cf == r_count_22_io_out ? io_r_719_b : _GEN_17308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17310 = 10'h2d0 == r_count_22_io_out ? io_r_720_b : _GEN_17309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17311 = 10'h2d1 == r_count_22_io_out ? io_r_721_b : _GEN_17310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17312 = 10'h2d2 == r_count_22_io_out ? io_r_722_b : _GEN_17311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17313 = 10'h2d3 == r_count_22_io_out ? io_r_723_b : _GEN_17312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17314 = 10'h2d4 == r_count_22_io_out ? io_r_724_b : _GEN_17313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17315 = 10'h2d5 == r_count_22_io_out ? io_r_725_b : _GEN_17314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17316 = 10'h2d6 == r_count_22_io_out ? io_r_726_b : _GEN_17315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17317 = 10'h2d7 == r_count_22_io_out ? io_r_727_b : _GEN_17316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17318 = 10'h2d8 == r_count_22_io_out ? io_r_728_b : _GEN_17317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17319 = 10'h2d9 == r_count_22_io_out ? io_r_729_b : _GEN_17318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17320 = 10'h2da == r_count_22_io_out ? io_r_730_b : _GEN_17319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17321 = 10'h2db == r_count_22_io_out ? io_r_731_b : _GEN_17320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17322 = 10'h2dc == r_count_22_io_out ? io_r_732_b : _GEN_17321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17323 = 10'h2dd == r_count_22_io_out ? io_r_733_b : _GEN_17322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17324 = 10'h2de == r_count_22_io_out ? io_r_734_b : _GEN_17323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17325 = 10'h2df == r_count_22_io_out ? io_r_735_b : _GEN_17324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17326 = 10'h2e0 == r_count_22_io_out ? io_r_736_b : _GEN_17325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17327 = 10'h2e1 == r_count_22_io_out ? io_r_737_b : _GEN_17326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17328 = 10'h2e2 == r_count_22_io_out ? io_r_738_b : _GEN_17327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17329 = 10'h2e3 == r_count_22_io_out ? io_r_739_b : _GEN_17328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17330 = 10'h2e4 == r_count_22_io_out ? io_r_740_b : _GEN_17329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17331 = 10'h2e5 == r_count_22_io_out ? io_r_741_b : _GEN_17330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17332 = 10'h2e6 == r_count_22_io_out ? io_r_742_b : _GEN_17331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17333 = 10'h2e7 == r_count_22_io_out ? io_r_743_b : _GEN_17332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17334 = 10'h2e8 == r_count_22_io_out ? io_r_744_b : _GEN_17333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17335 = 10'h2e9 == r_count_22_io_out ? io_r_745_b : _GEN_17334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17336 = 10'h2ea == r_count_22_io_out ? io_r_746_b : _GEN_17335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17337 = 10'h2eb == r_count_22_io_out ? io_r_747_b : _GEN_17336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17338 = 10'h2ec == r_count_22_io_out ? io_r_748_b : _GEN_17337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17341 = 10'h1 == r_count_23_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17342 = 10'h2 == r_count_23_io_out ? io_r_2_b : _GEN_17341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17343 = 10'h3 == r_count_23_io_out ? io_r_3_b : _GEN_17342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17344 = 10'h4 == r_count_23_io_out ? io_r_4_b : _GEN_17343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17345 = 10'h5 == r_count_23_io_out ? io_r_5_b : _GEN_17344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17346 = 10'h6 == r_count_23_io_out ? io_r_6_b : _GEN_17345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17347 = 10'h7 == r_count_23_io_out ? io_r_7_b : _GEN_17346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17348 = 10'h8 == r_count_23_io_out ? io_r_8_b : _GEN_17347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17349 = 10'h9 == r_count_23_io_out ? io_r_9_b : _GEN_17348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17350 = 10'ha == r_count_23_io_out ? io_r_10_b : _GEN_17349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17351 = 10'hb == r_count_23_io_out ? io_r_11_b : _GEN_17350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17352 = 10'hc == r_count_23_io_out ? io_r_12_b : _GEN_17351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17353 = 10'hd == r_count_23_io_out ? io_r_13_b : _GEN_17352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17354 = 10'he == r_count_23_io_out ? io_r_14_b : _GEN_17353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17355 = 10'hf == r_count_23_io_out ? io_r_15_b : _GEN_17354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17356 = 10'h10 == r_count_23_io_out ? io_r_16_b : _GEN_17355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17357 = 10'h11 == r_count_23_io_out ? io_r_17_b : _GEN_17356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17358 = 10'h12 == r_count_23_io_out ? io_r_18_b : _GEN_17357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17359 = 10'h13 == r_count_23_io_out ? io_r_19_b : _GEN_17358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17360 = 10'h14 == r_count_23_io_out ? io_r_20_b : _GEN_17359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17361 = 10'h15 == r_count_23_io_out ? io_r_21_b : _GEN_17360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17362 = 10'h16 == r_count_23_io_out ? io_r_22_b : _GEN_17361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17363 = 10'h17 == r_count_23_io_out ? io_r_23_b : _GEN_17362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17364 = 10'h18 == r_count_23_io_out ? io_r_24_b : _GEN_17363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17365 = 10'h19 == r_count_23_io_out ? io_r_25_b : _GEN_17364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17366 = 10'h1a == r_count_23_io_out ? io_r_26_b : _GEN_17365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17367 = 10'h1b == r_count_23_io_out ? io_r_27_b : _GEN_17366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17368 = 10'h1c == r_count_23_io_out ? io_r_28_b : _GEN_17367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17369 = 10'h1d == r_count_23_io_out ? io_r_29_b : _GEN_17368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17370 = 10'h1e == r_count_23_io_out ? io_r_30_b : _GEN_17369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17371 = 10'h1f == r_count_23_io_out ? io_r_31_b : _GEN_17370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17372 = 10'h20 == r_count_23_io_out ? io_r_32_b : _GEN_17371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17373 = 10'h21 == r_count_23_io_out ? io_r_33_b : _GEN_17372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17374 = 10'h22 == r_count_23_io_out ? io_r_34_b : _GEN_17373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17375 = 10'h23 == r_count_23_io_out ? io_r_35_b : _GEN_17374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17376 = 10'h24 == r_count_23_io_out ? io_r_36_b : _GEN_17375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17377 = 10'h25 == r_count_23_io_out ? io_r_37_b : _GEN_17376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17378 = 10'h26 == r_count_23_io_out ? io_r_38_b : _GEN_17377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17379 = 10'h27 == r_count_23_io_out ? io_r_39_b : _GEN_17378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17380 = 10'h28 == r_count_23_io_out ? io_r_40_b : _GEN_17379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17381 = 10'h29 == r_count_23_io_out ? io_r_41_b : _GEN_17380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17382 = 10'h2a == r_count_23_io_out ? io_r_42_b : _GEN_17381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17383 = 10'h2b == r_count_23_io_out ? io_r_43_b : _GEN_17382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17384 = 10'h2c == r_count_23_io_out ? io_r_44_b : _GEN_17383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17385 = 10'h2d == r_count_23_io_out ? io_r_45_b : _GEN_17384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17386 = 10'h2e == r_count_23_io_out ? io_r_46_b : _GEN_17385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17387 = 10'h2f == r_count_23_io_out ? io_r_47_b : _GEN_17386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17388 = 10'h30 == r_count_23_io_out ? io_r_48_b : _GEN_17387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17389 = 10'h31 == r_count_23_io_out ? io_r_49_b : _GEN_17388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17390 = 10'h32 == r_count_23_io_out ? io_r_50_b : _GEN_17389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17391 = 10'h33 == r_count_23_io_out ? io_r_51_b : _GEN_17390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17392 = 10'h34 == r_count_23_io_out ? io_r_52_b : _GEN_17391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17393 = 10'h35 == r_count_23_io_out ? io_r_53_b : _GEN_17392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17394 = 10'h36 == r_count_23_io_out ? io_r_54_b : _GEN_17393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17395 = 10'h37 == r_count_23_io_out ? io_r_55_b : _GEN_17394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17396 = 10'h38 == r_count_23_io_out ? io_r_56_b : _GEN_17395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17397 = 10'h39 == r_count_23_io_out ? io_r_57_b : _GEN_17396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17398 = 10'h3a == r_count_23_io_out ? io_r_58_b : _GEN_17397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17399 = 10'h3b == r_count_23_io_out ? io_r_59_b : _GEN_17398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17400 = 10'h3c == r_count_23_io_out ? io_r_60_b : _GEN_17399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17401 = 10'h3d == r_count_23_io_out ? io_r_61_b : _GEN_17400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17402 = 10'h3e == r_count_23_io_out ? io_r_62_b : _GEN_17401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17403 = 10'h3f == r_count_23_io_out ? io_r_63_b : _GEN_17402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17404 = 10'h40 == r_count_23_io_out ? io_r_64_b : _GEN_17403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17405 = 10'h41 == r_count_23_io_out ? io_r_65_b : _GEN_17404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17406 = 10'h42 == r_count_23_io_out ? io_r_66_b : _GEN_17405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17407 = 10'h43 == r_count_23_io_out ? io_r_67_b : _GEN_17406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17408 = 10'h44 == r_count_23_io_out ? io_r_68_b : _GEN_17407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17409 = 10'h45 == r_count_23_io_out ? io_r_69_b : _GEN_17408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17410 = 10'h46 == r_count_23_io_out ? io_r_70_b : _GEN_17409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17411 = 10'h47 == r_count_23_io_out ? io_r_71_b : _GEN_17410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17412 = 10'h48 == r_count_23_io_out ? io_r_72_b : _GEN_17411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17413 = 10'h49 == r_count_23_io_out ? io_r_73_b : _GEN_17412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17414 = 10'h4a == r_count_23_io_out ? io_r_74_b : _GEN_17413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17415 = 10'h4b == r_count_23_io_out ? io_r_75_b : _GEN_17414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17416 = 10'h4c == r_count_23_io_out ? io_r_76_b : _GEN_17415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17417 = 10'h4d == r_count_23_io_out ? io_r_77_b : _GEN_17416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17418 = 10'h4e == r_count_23_io_out ? io_r_78_b : _GEN_17417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17419 = 10'h4f == r_count_23_io_out ? io_r_79_b : _GEN_17418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17420 = 10'h50 == r_count_23_io_out ? io_r_80_b : _GEN_17419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17421 = 10'h51 == r_count_23_io_out ? io_r_81_b : _GEN_17420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17422 = 10'h52 == r_count_23_io_out ? io_r_82_b : _GEN_17421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17423 = 10'h53 == r_count_23_io_out ? io_r_83_b : _GEN_17422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17424 = 10'h54 == r_count_23_io_out ? io_r_84_b : _GEN_17423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17425 = 10'h55 == r_count_23_io_out ? io_r_85_b : _GEN_17424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17426 = 10'h56 == r_count_23_io_out ? io_r_86_b : _GEN_17425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17427 = 10'h57 == r_count_23_io_out ? io_r_87_b : _GEN_17426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17428 = 10'h58 == r_count_23_io_out ? io_r_88_b : _GEN_17427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17429 = 10'h59 == r_count_23_io_out ? io_r_89_b : _GEN_17428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17430 = 10'h5a == r_count_23_io_out ? io_r_90_b : _GEN_17429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17431 = 10'h5b == r_count_23_io_out ? io_r_91_b : _GEN_17430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17432 = 10'h5c == r_count_23_io_out ? io_r_92_b : _GEN_17431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17433 = 10'h5d == r_count_23_io_out ? io_r_93_b : _GEN_17432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17434 = 10'h5e == r_count_23_io_out ? io_r_94_b : _GEN_17433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17435 = 10'h5f == r_count_23_io_out ? io_r_95_b : _GEN_17434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17436 = 10'h60 == r_count_23_io_out ? io_r_96_b : _GEN_17435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17437 = 10'h61 == r_count_23_io_out ? io_r_97_b : _GEN_17436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17438 = 10'h62 == r_count_23_io_out ? io_r_98_b : _GEN_17437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17439 = 10'h63 == r_count_23_io_out ? io_r_99_b : _GEN_17438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17440 = 10'h64 == r_count_23_io_out ? io_r_100_b : _GEN_17439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17441 = 10'h65 == r_count_23_io_out ? io_r_101_b : _GEN_17440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17442 = 10'h66 == r_count_23_io_out ? io_r_102_b : _GEN_17441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17443 = 10'h67 == r_count_23_io_out ? io_r_103_b : _GEN_17442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17444 = 10'h68 == r_count_23_io_out ? io_r_104_b : _GEN_17443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17445 = 10'h69 == r_count_23_io_out ? io_r_105_b : _GEN_17444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17446 = 10'h6a == r_count_23_io_out ? io_r_106_b : _GEN_17445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17447 = 10'h6b == r_count_23_io_out ? io_r_107_b : _GEN_17446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17448 = 10'h6c == r_count_23_io_out ? io_r_108_b : _GEN_17447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17449 = 10'h6d == r_count_23_io_out ? io_r_109_b : _GEN_17448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17450 = 10'h6e == r_count_23_io_out ? io_r_110_b : _GEN_17449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17451 = 10'h6f == r_count_23_io_out ? io_r_111_b : _GEN_17450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17452 = 10'h70 == r_count_23_io_out ? io_r_112_b : _GEN_17451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17453 = 10'h71 == r_count_23_io_out ? io_r_113_b : _GEN_17452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17454 = 10'h72 == r_count_23_io_out ? io_r_114_b : _GEN_17453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17455 = 10'h73 == r_count_23_io_out ? io_r_115_b : _GEN_17454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17456 = 10'h74 == r_count_23_io_out ? io_r_116_b : _GEN_17455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17457 = 10'h75 == r_count_23_io_out ? io_r_117_b : _GEN_17456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17458 = 10'h76 == r_count_23_io_out ? io_r_118_b : _GEN_17457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17459 = 10'h77 == r_count_23_io_out ? io_r_119_b : _GEN_17458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17460 = 10'h78 == r_count_23_io_out ? io_r_120_b : _GEN_17459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17461 = 10'h79 == r_count_23_io_out ? io_r_121_b : _GEN_17460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17462 = 10'h7a == r_count_23_io_out ? io_r_122_b : _GEN_17461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17463 = 10'h7b == r_count_23_io_out ? io_r_123_b : _GEN_17462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17464 = 10'h7c == r_count_23_io_out ? io_r_124_b : _GEN_17463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17465 = 10'h7d == r_count_23_io_out ? io_r_125_b : _GEN_17464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17466 = 10'h7e == r_count_23_io_out ? io_r_126_b : _GEN_17465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17467 = 10'h7f == r_count_23_io_out ? io_r_127_b : _GEN_17466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17468 = 10'h80 == r_count_23_io_out ? io_r_128_b : _GEN_17467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17469 = 10'h81 == r_count_23_io_out ? io_r_129_b : _GEN_17468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17470 = 10'h82 == r_count_23_io_out ? io_r_130_b : _GEN_17469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17471 = 10'h83 == r_count_23_io_out ? io_r_131_b : _GEN_17470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17472 = 10'h84 == r_count_23_io_out ? io_r_132_b : _GEN_17471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17473 = 10'h85 == r_count_23_io_out ? io_r_133_b : _GEN_17472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17474 = 10'h86 == r_count_23_io_out ? io_r_134_b : _GEN_17473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17475 = 10'h87 == r_count_23_io_out ? io_r_135_b : _GEN_17474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17476 = 10'h88 == r_count_23_io_out ? io_r_136_b : _GEN_17475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17477 = 10'h89 == r_count_23_io_out ? io_r_137_b : _GEN_17476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17478 = 10'h8a == r_count_23_io_out ? io_r_138_b : _GEN_17477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17479 = 10'h8b == r_count_23_io_out ? io_r_139_b : _GEN_17478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17480 = 10'h8c == r_count_23_io_out ? io_r_140_b : _GEN_17479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17481 = 10'h8d == r_count_23_io_out ? io_r_141_b : _GEN_17480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17482 = 10'h8e == r_count_23_io_out ? io_r_142_b : _GEN_17481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17483 = 10'h8f == r_count_23_io_out ? io_r_143_b : _GEN_17482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17484 = 10'h90 == r_count_23_io_out ? io_r_144_b : _GEN_17483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17485 = 10'h91 == r_count_23_io_out ? io_r_145_b : _GEN_17484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17486 = 10'h92 == r_count_23_io_out ? io_r_146_b : _GEN_17485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17487 = 10'h93 == r_count_23_io_out ? io_r_147_b : _GEN_17486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17488 = 10'h94 == r_count_23_io_out ? io_r_148_b : _GEN_17487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17489 = 10'h95 == r_count_23_io_out ? io_r_149_b : _GEN_17488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17490 = 10'h96 == r_count_23_io_out ? io_r_150_b : _GEN_17489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17491 = 10'h97 == r_count_23_io_out ? io_r_151_b : _GEN_17490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17492 = 10'h98 == r_count_23_io_out ? io_r_152_b : _GEN_17491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17493 = 10'h99 == r_count_23_io_out ? io_r_153_b : _GEN_17492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17494 = 10'h9a == r_count_23_io_out ? io_r_154_b : _GEN_17493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17495 = 10'h9b == r_count_23_io_out ? io_r_155_b : _GEN_17494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17496 = 10'h9c == r_count_23_io_out ? io_r_156_b : _GEN_17495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17497 = 10'h9d == r_count_23_io_out ? io_r_157_b : _GEN_17496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17498 = 10'h9e == r_count_23_io_out ? io_r_158_b : _GEN_17497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17499 = 10'h9f == r_count_23_io_out ? io_r_159_b : _GEN_17498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17500 = 10'ha0 == r_count_23_io_out ? io_r_160_b : _GEN_17499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17501 = 10'ha1 == r_count_23_io_out ? io_r_161_b : _GEN_17500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17502 = 10'ha2 == r_count_23_io_out ? io_r_162_b : _GEN_17501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17503 = 10'ha3 == r_count_23_io_out ? io_r_163_b : _GEN_17502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17504 = 10'ha4 == r_count_23_io_out ? io_r_164_b : _GEN_17503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17505 = 10'ha5 == r_count_23_io_out ? io_r_165_b : _GEN_17504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17506 = 10'ha6 == r_count_23_io_out ? io_r_166_b : _GEN_17505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17507 = 10'ha7 == r_count_23_io_out ? io_r_167_b : _GEN_17506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17508 = 10'ha8 == r_count_23_io_out ? io_r_168_b : _GEN_17507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17509 = 10'ha9 == r_count_23_io_out ? io_r_169_b : _GEN_17508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17510 = 10'haa == r_count_23_io_out ? io_r_170_b : _GEN_17509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17511 = 10'hab == r_count_23_io_out ? io_r_171_b : _GEN_17510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17512 = 10'hac == r_count_23_io_out ? io_r_172_b : _GEN_17511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17513 = 10'had == r_count_23_io_out ? io_r_173_b : _GEN_17512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17514 = 10'hae == r_count_23_io_out ? io_r_174_b : _GEN_17513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17515 = 10'haf == r_count_23_io_out ? io_r_175_b : _GEN_17514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17516 = 10'hb0 == r_count_23_io_out ? io_r_176_b : _GEN_17515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17517 = 10'hb1 == r_count_23_io_out ? io_r_177_b : _GEN_17516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17518 = 10'hb2 == r_count_23_io_out ? io_r_178_b : _GEN_17517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17519 = 10'hb3 == r_count_23_io_out ? io_r_179_b : _GEN_17518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17520 = 10'hb4 == r_count_23_io_out ? io_r_180_b : _GEN_17519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17521 = 10'hb5 == r_count_23_io_out ? io_r_181_b : _GEN_17520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17522 = 10'hb6 == r_count_23_io_out ? io_r_182_b : _GEN_17521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17523 = 10'hb7 == r_count_23_io_out ? io_r_183_b : _GEN_17522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17524 = 10'hb8 == r_count_23_io_out ? io_r_184_b : _GEN_17523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17525 = 10'hb9 == r_count_23_io_out ? io_r_185_b : _GEN_17524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17526 = 10'hba == r_count_23_io_out ? io_r_186_b : _GEN_17525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17527 = 10'hbb == r_count_23_io_out ? io_r_187_b : _GEN_17526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17528 = 10'hbc == r_count_23_io_out ? io_r_188_b : _GEN_17527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17529 = 10'hbd == r_count_23_io_out ? io_r_189_b : _GEN_17528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17530 = 10'hbe == r_count_23_io_out ? io_r_190_b : _GEN_17529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17531 = 10'hbf == r_count_23_io_out ? io_r_191_b : _GEN_17530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17532 = 10'hc0 == r_count_23_io_out ? io_r_192_b : _GEN_17531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17533 = 10'hc1 == r_count_23_io_out ? io_r_193_b : _GEN_17532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17534 = 10'hc2 == r_count_23_io_out ? io_r_194_b : _GEN_17533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17535 = 10'hc3 == r_count_23_io_out ? io_r_195_b : _GEN_17534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17536 = 10'hc4 == r_count_23_io_out ? io_r_196_b : _GEN_17535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17537 = 10'hc5 == r_count_23_io_out ? io_r_197_b : _GEN_17536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17538 = 10'hc6 == r_count_23_io_out ? io_r_198_b : _GEN_17537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17539 = 10'hc7 == r_count_23_io_out ? io_r_199_b : _GEN_17538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17540 = 10'hc8 == r_count_23_io_out ? io_r_200_b : _GEN_17539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17541 = 10'hc9 == r_count_23_io_out ? io_r_201_b : _GEN_17540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17542 = 10'hca == r_count_23_io_out ? io_r_202_b : _GEN_17541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17543 = 10'hcb == r_count_23_io_out ? io_r_203_b : _GEN_17542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17544 = 10'hcc == r_count_23_io_out ? io_r_204_b : _GEN_17543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17545 = 10'hcd == r_count_23_io_out ? io_r_205_b : _GEN_17544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17546 = 10'hce == r_count_23_io_out ? io_r_206_b : _GEN_17545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17547 = 10'hcf == r_count_23_io_out ? io_r_207_b : _GEN_17546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17548 = 10'hd0 == r_count_23_io_out ? io_r_208_b : _GEN_17547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17549 = 10'hd1 == r_count_23_io_out ? io_r_209_b : _GEN_17548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17550 = 10'hd2 == r_count_23_io_out ? io_r_210_b : _GEN_17549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17551 = 10'hd3 == r_count_23_io_out ? io_r_211_b : _GEN_17550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17552 = 10'hd4 == r_count_23_io_out ? io_r_212_b : _GEN_17551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17553 = 10'hd5 == r_count_23_io_out ? io_r_213_b : _GEN_17552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17554 = 10'hd6 == r_count_23_io_out ? io_r_214_b : _GEN_17553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17555 = 10'hd7 == r_count_23_io_out ? io_r_215_b : _GEN_17554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17556 = 10'hd8 == r_count_23_io_out ? io_r_216_b : _GEN_17555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17557 = 10'hd9 == r_count_23_io_out ? io_r_217_b : _GEN_17556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17558 = 10'hda == r_count_23_io_out ? io_r_218_b : _GEN_17557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17559 = 10'hdb == r_count_23_io_out ? io_r_219_b : _GEN_17558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17560 = 10'hdc == r_count_23_io_out ? io_r_220_b : _GEN_17559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17561 = 10'hdd == r_count_23_io_out ? io_r_221_b : _GEN_17560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17562 = 10'hde == r_count_23_io_out ? io_r_222_b : _GEN_17561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17563 = 10'hdf == r_count_23_io_out ? io_r_223_b : _GEN_17562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17564 = 10'he0 == r_count_23_io_out ? io_r_224_b : _GEN_17563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17565 = 10'he1 == r_count_23_io_out ? io_r_225_b : _GEN_17564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17566 = 10'he2 == r_count_23_io_out ? io_r_226_b : _GEN_17565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17567 = 10'he3 == r_count_23_io_out ? io_r_227_b : _GEN_17566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17568 = 10'he4 == r_count_23_io_out ? io_r_228_b : _GEN_17567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17569 = 10'he5 == r_count_23_io_out ? io_r_229_b : _GEN_17568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17570 = 10'he6 == r_count_23_io_out ? io_r_230_b : _GEN_17569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17571 = 10'he7 == r_count_23_io_out ? io_r_231_b : _GEN_17570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17572 = 10'he8 == r_count_23_io_out ? io_r_232_b : _GEN_17571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17573 = 10'he9 == r_count_23_io_out ? io_r_233_b : _GEN_17572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17574 = 10'hea == r_count_23_io_out ? io_r_234_b : _GEN_17573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17575 = 10'heb == r_count_23_io_out ? io_r_235_b : _GEN_17574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17576 = 10'hec == r_count_23_io_out ? io_r_236_b : _GEN_17575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17577 = 10'hed == r_count_23_io_out ? io_r_237_b : _GEN_17576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17578 = 10'hee == r_count_23_io_out ? io_r_238_b : _GEN_17577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17579 = 10'hef == r_count_23_io_out ? io_r_239_b : _GEN_17578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17580 = 10'hf0 == r_count_23_io_out ? io_r_240_b : _GEN_17579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17581 = 10'hf1 == r_count_23_io_out ? io_r_241_b : _GEN_17580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17582 = 10'hf2 == r_count_23_io_out ? io_r_242_b : _GEN_17581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17583 = 10'hf3 == r_count_23_io_out ? io_r_243_b : _GEN_17582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17584 = 10'hf4 == r_count_23_io_out ? io_r_244_b : _GEN_17583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17585 = 10'hf5 == r_count_23_io_out ? io_r_245_b : _GEN_17584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17586 = 10'hf6 == r_count_23_io_out ? io_r_246_b : _GEN_17585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17587 = 10'hf7 == r_count_23_io_out ? io_r_247_b : _GEN_17586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17588 = 10'hf8 == r_count_23_io_out ? io_r_248_b : _GEN_17587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17589 = 10'hf9 == r_count_23_io_out ? io_r_249_b : _GEN_17588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17590 = 10'hfa == r_count_23_io_out ? io_r_250_b : _GEN_17589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17591 = 10'hfb == r_count_23_io_out ? io_r_251_b : _GEN_17590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17592 = 10'hfc == r_count_23_io_out ? io_r_252_b : _GEN_17591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17593 = 10'hfd == r_count_23_io_out ? io_r_253_b : _GEN_17592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17594 = 10'hfe == r_count_23_io_out ? io_r_254_b : _GEN_17593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17595 = 10'hff == r_count_23_io_out ? io_r_255_b : _GEN_17594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17596 = 10'h100 == r_count_23_io_out ? io_r_256_b : _GEN_17595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17597 = 10'h101 == r_count_23_io_out ? io_r_257_b : _GEN_17596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17598 = 10'h102 == r_count_23_io_out ? io_r_258_b : _GEN_17597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17599 = 10'h103 == r_count_23_io_out ? io_r_259_b : _GEN_17598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17600 = 10'h104 == r_count_23_io_out ? io_r_260_b : _GEN_17599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17601 = 10'h105 == r_count_23_io_out ? io_r_261_b : _GEN_17600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17602 = 10'h106 == r_count_23_io_out ? io_r_262_b : _GEN_17601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17603 = 10'h107 == r_count_23_io_out ? io_r_263_b : _GEN_17602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17604 = 10'h108 == r_count_23_io_out ? io_r_264_b : _GEN_17603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17605 = 10'h109 == r_count_23_io_out ? io_r_265_b : _GEN_17604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17606 = 10'h10a == r_count_23_io_out ? io_r_266_b : _GEN_17605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17607 = 10'h10b == r_count_23_io_out ? io_r_267_b : _GEN_17606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17608 = 10'h10c == r_count_23_io_out ? io_r_268_b : _GEN_17607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17609 = 10'h10d == r_count_23_io_out ? io_r_269_b : _GEN_17608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17610 = 10'h10e == r_count_23_io_out ? io_r_270_b : _GEN_17609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17611 = 10'h10f == r_count_23_io_out ? io_r_271_b : _GEN_17610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17612 = 10'h110 == r_count_23_io_out ? io_r_272_b : _GEN_17611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17613 = 10'h111 == r_count_23_io_out ? io_r_273_b : _GEN_17612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17614 = 10'h112 == r_count_23_io_out ? io_r_274_b : _GEN_17613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17615 = 10'h113 == r_count_23_io_out ? io_r_275_b : _GEN_17614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17616 = 10'h114 == r_count_23_io_out ? io_r_276_b : _GEN_17615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17617 = 10'h115 == r_count_23_io_out ? io_r_277_b : _GEN_17616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17618 = 10'h116 == r_count_23_io_out ? io_r_278_b : _GEN_17617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17619 = 10'h117 == r_count_23_io_out ? io_r_279_b : _GEN_17618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17620 = 10'h118 == r_count_23_io_out ? io_r_280_b : _GEN_17619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17621 = 10'h119 == r_count_23_io_out ? io_r_281_b : _GEN_17620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17622 = 10'h11a == r_count_23_io_out ? io_r_282_b : _GEN_17621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17623 = 10'h11b == r_count_23_io_out ? io_r_283_b : _GEN_17622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17624 = 10'h11c == r_count_23_io_out ? io_r_284_b : _GEN_17623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17625 = 10'h11d == r_count_23_io_out ? io_r_285_b : _GEN_17624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17626 = 10'h11e == r_count_23_io_out ? io_r_286_b : _GEN_17625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17627 = 10'h11f == r_count_23_io_out ? io_r_287_b : _GEN_17626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17628 = 10'h120 == r_count_23_io_out ? io_r_288_b : _GEN_17627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17629 = 10'h121 == r_count_23_io_out ? io_r_289_b : _GEN_17628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17630 = 10'h122 == r_count_23_io_out ? io_r_290_b : _GEN_17629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17631 = 10'h123 == r_count_23_io_out ? io_r_291_b : _GEN_17630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17632 = 10'h124 == r_count_23_io_out ? io_r_292_b : _GEN_17631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17633 = 10'h125 == r_count_23_io_out ? io_r_293_b : _GEN_17632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17634 = 10'h126 == r_count_23_io_out ? io_r_294_b : _GEN_17633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17635 = 10'h127 == r_count_23_io_out ? io_r_295_b : _GEN_17634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17636 = 10'h128 == r_count_23_io_out ? io_r_296_b : _GEN_17635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17637 = 10'h129 == r_count_23_io_out ? io_r_297_b : _GEN_17636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17638 = 10'h12a == r_count_23_io_out ? io_r_298_b : _GEN_17637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17639 = 10'h12b == r_count_23_io_out ? io_r_299_b : _GEN_17638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17640 = 10'h12c == r_count_23_io_out ? io_r_300_b : _GEN_17639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17641 = 10'h12d == r_count_23_io_out ? io_r_301_b : _GEN_17640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17642 = 10'h12e == r_count_23_io_out ? io_r_302_b : _GEN_17641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17643 = 10'h12f == r_count_23_io_out ? io_r_303_b : _GEN_17642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17644 = 10'h130 == r_count_23_io_out ? io_r_304_b : _GEN_17643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17645 = 10'h131 == r_count_23_io_out ? io_r_305_b : _GEN_17644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17646 = 10'h132 == r_count_23_io_out ? io_r_306_b : _GEN_17645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17647 = 10'h133 == r_count_23_io_out ? io_r_307_b : _GEN_17646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17648 = 10'h134 == r_count_23_io_out ? io_r_308_b : _GEN_17647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17649 = 10'h135 == r_count_23_io_out ? io_r_309_b : _GEN_17648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17650 = 10'h136 == r_count_23_io_out ? io_r_310_b : _GEN_17649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17651 = 10'h137 == r_count_23_io_out ? io_r_311_b : _GEN_17650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17652 = 10'h138 == r_count_23_io_out ? io_r_312_b : _GEN_17651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17653 = 10'h139 == r_count_23_io_out ? io_r_313_b : _GEN_17652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17654 = 10'h13a == r_count_23_io_out ? io_r_314_b : _GEN_17653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17655 = 10'h13b == r_count_23_io_out ? io_r_315_b : _GEN_17654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17656 = 10'h13c == r_count_23_io_out ? io_r_316_b : _GEN_17655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17657 = 10'h13d == r_count_23_io_out ? io_r_317_b : _GEN_17656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17658 = 10'h13e == r_count_23_io_out ? io_r_318_b : _GEN_17657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17659 = 10'h13f == r_count_23_io_out ? io_r_319_b : _GEN_17658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17660 = 10'h140 == r_count_23_io_out ? io_r_320_b : _GEN_17659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17661 = 10'h141 == r_count_23_io_out ? io_r_321_b : _GEN_17660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17662 = 10'h142 == r_count_23_io_out ? io_r_322_b : _GEN_17661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17663 = 10'h143 == r_count_23_io_out ? io_r_323_b : _GEN_17662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17664 = 10'h144 == r_count_23_io_out ? io_r_324_b : _GEN_17663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17665 = 10'h145 == r_count_23_io_out ? io_r_325_b : _GEN_17664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17666 = 10'h146 == r_count_23_io_out ? io_r_326_b : _GEN_17665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17667 = 10'h147 == r_count_23_io_out ? io_r_327_b : _GEN_17666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17668 = 10'h148 == r_count_23_io_out ? io_r_328_b : _GEN_17667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17669 = 10'h149 == r_count_23_io_out ? io_r_329_b : _GEN_17668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17670 = 10'h14a == r_count_23_io_out ? io_r_330_b : _GEN_17669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17671 = 10'h14b == r_count_23_io_out ? io_r_331_b : _GEN_17670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17672 = 10'h14c == r_count_23_io_out ? io_r_332_b : _GEN_17671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17673 = 10'h14d == r_count_23_io_out ? io_r_333_b : _GEN_17672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17674 = 10'h14e == r_count_23_io_out ? io_r_334_b : _GEN_17673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17675 = 10'h14f == r_count_23_io_out ? io_r_335_b : _GEN_17674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17676 = 10'h150 == r_count_23_io_out ? io_r_336_b : _GEN_17675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17677 = 10'h151 == r_count_23_io_out ? io_r_337_b : _GEN_17676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17678 = 10'h152 == r_count_23_io_out ? io_r_338_b : _GEN_17677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17679 = 10'h153 == r_count_23_io_out ? io_r_339_b : _GEN_17678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17680 = 10'h154 == r_count_23_io_out ? io_r_340_b : _GEN_17679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17681 = 10'h155 == r_count_23_io_out ? io_r_341_b : _GEN_17680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17682 = 10'h156 == r_count_23_io_out ? io_r_342_b : _GEN_17681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17683 = 10'h157 == r_count_23_io_out ? io_r_343_b : _GEN_17682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17684 = 10'h158 == r_count_23_io_out ? io_r_344_b : _GEN_17683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17685 = 10'h159 == r_count_23_io_out ? io_r_345_b : _GEN_17684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17686 = 10'h15a == r_count_23_io_out ? io_r_346_b : _GEN_17685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17687 = 10'h15b == r_count_23_io_out ? io_r_347_b : _GEN_17686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17688 = 10'h15c == r_count_23_io_out ? io_r_348_b : _GEN_17687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17689 = 10'h15d == r_count_23_io_out ? io_r_349_b : _GEN_17688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17690 = 10'h15e == r_count_23_io_out ? io_r_350_b : _GEN_17689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17691 = 10'h15f == r_count_23_io_out ? io_r_351_b : _GEN_17690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17692 = 10'h160 == r_count_23_io_out ? io_r_352_b : _GEN_17691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17693 = 10'h161 == r_count_23_io_out ? io_r_353_b : _GEN_17692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17694 = 10'h162 == r_count_23_io_out ? io_r_354_b : _GEN_17693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17695 = 10'h163 == r_count_23_io_out ? io_r_355_b : _GEN_17694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17696 = 10'h164 == r_count_23_io_out ? io_r_356_b : _GEN_17695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17697 = 10'h165 == r_count_23_io_out ? io_r_357_b : _GEN_17696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17698 = 10'h166 == r_count_23_io_out ? io_r_358_b : _GEN_17697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17699 = 10'h167 == r_count_23_io_out ? io_r_359_b : _GEN_17698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17700 = 10'h168 == r_count_23_io_out ? io_r_360_b : _GEN_17699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17701 = 10'h169 == r_count_23_io_out ? io_r_361_b : _GEN_17700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17702 = 10'h16a == r_count_23_io_out ? io_r_362_b : _GEN_17701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17703 = 10'h16b == r_count_23_io_out ? io_r_363_b : _GEN_17702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17704 = 10'h16c == r_count_23_io_out ? io_r_364_b : _GEN_17703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17705 = 10'h16d == r_count_23_io_out ? io_r_365_b : _GEN_17704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17706 = 10'h16e == r_count_23_io_out ? io_r_366_b : _GEN_17705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17707 = 10'h16f == r_count_23_io_out ? io_r_367_b : _GEN_17706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17708 = 10'h170 == r_count_23_io_out ? io_r_368_b : _GEN_17707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17709 = 10'h171 == r_count_23_io_out ? io_r_369_b : _GEN_17708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17710 = 10'h172 == r_count_23_io_out ? io_r_370_b : _GEN_17709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17711 = 10'h173 == r_count_23_io_out ? io_r_371_b : _GEN_17710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17712 = 10'h174 == r_count_23_io_out ? io_r_372_b : _GEN_17711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17713 = 10'h175 == r_count_23_io_out ? io_r_373_b : _GEN_17712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17714 = 10'h176 == r_count_23_io_out ? io_r_374_b : _GEN_17713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17715 = 10'h177 == r_count_23_io_out ? io_r_375_b : _GEN_17714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17716 = 10'h178 == r_count_23_io_out ? io_r_376_b : _GEN_17715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17717 = 10'h179 == r_count_23_io_out ? io_r_377_b : _GEN_17716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17718 = 10'h17a == r_count_23_io_out ? io_r_378_b : _GEN_17717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17719 = 10'h17b == r_count_23_io_out ? io_r_379_b : _GEN_17718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17720 = 10'h17c == r_count_23_io_out ? io_r_380_b : _GEN_17719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17721 = 10'h17d == r_count_23_io_out ? io_r_381_b : _GEN_17720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17722 = 10'h17e == r_count_23_io_out ? io_r_382_b : _GEN_17721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17723 = 10'h17f == r_count_23_io_out ? io_r_383_b : _GEN_17722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17724 = 10'h180 == r_count_23_io_out ? io_r_384_b : _GEN_17723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17725 = 10'h181 == r_count_23_io_out ? io_r_385_b : _GEN_17724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17726 = 10'h182 == r_count_23_io_out ? io_r_386_b : _GEN_17725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17727 = 10'h183 == r_count_23_io_out ? io_r_387_b : _GEN_17726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17728 = 10'h184 == r_count_23_io_out ? io_r_388_b : _GEN_17727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17729 = 10'h185 == r_count_23_io_out ? io_r_389_b : _GEN_17728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17730 = 10'h186 == r_count_23_io_out ? io_r_390_b : _GEN_17729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17731 = 10'h187 == r_count_23_io_out ? io_r_391_b : _GEN_17730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17732 = 10'h188 == r_count_23_io_out ? io_r_392_b : _GEN_17731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17733 = 10'h189 == r_count_23_io_out ? io_r_393_b : _GEN_17732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17734 = 10'h18a == r_count_23_io_out ? io_r_394_b : _GEN_17733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17735 = 10'h18b == r_count_23_io_out ? io_r_395_b : _GEN_17734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17736 = 10'h18c == r_count_23_io_out ? io_r_396_b : _GEN_17735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17737 = 10'h18d == r_count_23_io_out ? io_r_397_b : _GEN_17736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17738 = 10'h18e == r_count_23_io_out ? io_r_398_b : _GEN_17737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17739 = 10'h18f == r_count_23_io_out ? io_r_399_b : _GEN_17738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17740 = 10'h190 == r_count_23_io_out ? io_r_400_b : _GEN_17739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17741 = 10'h191 == r_count_23_io_out ? io_r_401_b : _GEN_17740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17742 = 10'h192 == r_count_23_io_out ? io_r_402_b : _GEN_17741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17743 = 10'h193 == r_count_23_io_out ? io_r_403_b : _GEN_17742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17744 = 10'h194 == r_count_23_io_out ? io_r_404_b : _GEN_17743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17745 = 10'h195 == r_count_23_io_out ? io_r_405_b : _GEN_17744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17746 = 10'h196 == r_count_23_io_out ? io_r_406_b : _GEN_17745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17747 = 10'h197 == r_count_23_io_out ? io_r_407_b : _GEN_17746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17748 = 10'h198 == r_count_23_io_out ? io_r_408_b : _GEN_17747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17749 = 10'h199 == r_count_23_io_out ? io_r_409_b : _GEN_17748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17750 = 10'h19a == r_count_23_io_out ? io_r_410_b : _GEN_17749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17751 = 10'h19b == r_count_23_io_out ? io_r_411_b : _GEN_17750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17752 = 10'h19c == r_count_23_io_out ? io_r_412_b : _GEN_17751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17753 = 10'h19d == r_count_23_io_out ? io_r_413_b : _GEN_17752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17754 = 10'h19e == r_count_23_io_out ? io_r_414_b : _GEN_17753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17755 = 10'h19f == r_count_23_io_out ? io_r_415_b : _GEN_17754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17756 = 10'h1a0 == r_count_23_io_out ? io_r_416_b : _GEN_17755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17757 = 10'h1a1 == r_count_23_io_out ? io_r_417_b : _GEN_17756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17758 = 10'h1a2 == r_count_23_io_out ? io_r_418_b : _GEN_17757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17759 = 10'h1a3 == r_count_23_io_out ? io_r_419_b : _GEN_17758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17760 = 10'h1a4 == r_count_23_io_out ? io_r_420_b : _GEN_17759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17761 = 10'h1a5 == r_count_23_io_out ? io_r_421_b : _GEN_17760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17762 = 10'h1a6 == r_count_23_io_out ? io_r_422_b : _GEN_17761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17763 = 10'h1a7 == r_count_23_io_out ? io_r_423_b : _GEN_17762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17764 = 10'h1a8 == r_count_23_io_out ? io_r_424_b : _GEN_17763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17765 = 10'h1a9 == r_count_23_io_out ? io_r_425_b : _GEN_17764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17766 = 10'h1aa == r_count_23_io_out ? io_r_426_b : _GEN_17765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17767 = 10'h1ab == r_count_23_io_out ? io_r_427_b : _GEN_17766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17768 = 10'h1ac == r_count_23_io_out ? io_r_428_b : _GEN_17767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17769 = 10'h1ad == r_count_23_io_out ? io_r_429_b : _GEN_17768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17770 = 10'h1ae == r_count_23_io_out ? io_r_430_b : _GEN_17769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17771 = 10'h1af == r_count_23_io_out ? io_r_431_b : _GEN_17770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17772 = 10'h1b0 == r_count_23_io_out ? io_r_432_b : _GEN_17771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17773 = 10'h1b1 == r_count_23_io_out ? io_r_433_b : _GEN_17772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17774 = 10'h1b2 == r_count_23_io_out ? io_r_434_b : _GEN_17773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17775 = 10'h1b3 == r_count_23_io_out ? io_r_435_b : _GEN_17774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17776 = 10'h1b4 == r_count_23_io_out ? io_r_436_b : _GEN_17775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17777 = 10'h1b5 == r_count_23_io_out ? io_r_437_b : _GEN_17776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17778 = 10'h1b6 == r_count_23_io_out ? io_r_438_b : _GEN_17777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17779 = 10'h1b7 == r_count_23_io_out ? io_r_439_b : _GEN_17778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17780 = 10'h1b8 == r_count_23_io_out ? io_r_440_b : _GEN_17779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17781 = 10'h1b9 == r_count_23_io_out ? io_r_441_b : _GEN_17780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17782 = 10'h1ba == r_count_23_io_out ? io_r_442_b : _GEN_17781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17783 = 10'h1bb == r_count_23_io_out ? io_r_443_b : _GEN_17782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17784 = 10'h1bc == r_count_23_io_out ? io_r_444_b : _GEN_17783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17785 = 10'h1bd == r_count_23_io_out ? io_r_445_b : _GEN_17784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17786 = 10'h1be == r_count_23_io_out ? io_r_446_b : _GEN_17785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17787 = 10'h1bf == r_count_23_io_out ? io_r_447_b : _GEN_17786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17788 = 10'h1c0 == r_count_23_io_out ? io_r_448_b : _GEN_17787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17789 = 10'h1c1 == r_count_23_io_out ? io_r_449_b : _GEN_17788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17790 = 10'h1c2 == r_count_23_io_out ? io_r_450_b : _GEN_17789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17791 = 10'h1c3 == r_count_23_io_out ? io_r_451_b : _GEN_17790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17792 = 10'h1c4 == r_count_23_io_out ? io_r_452_b : _GEN_17791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17793 = 10'h1c5 == r_count_23_io_out ? io_r_453_b : _GEN_17792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17794 = 10'h1c6 == r_count_23_io_out ? io_r_454_b : _GEN_17793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17795 = 10'h1c7 == r_count_23_io_out ? io_r_455_b : _GEN_17794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17796 = 10'h1c8 == r_count_23_io_out ? io_r_456_b : _GEN_17795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17797 = 10'h1c9 == r_count_23_io_out ? io_r_457_b : _GEN_17796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17798 = 10'h1ca == r_count_23_io_out ? io_r_458_b : _GEN_17797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17799 = 10'h1cb == r_count_23_io_out ? io_r_459_b : _GEN_17798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17800 = 10'h1cc == r_count_23_io_out ? io_r_460_b : _GEN_17799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17801 = 10'h1cd == r_count_23_io_out ? io_r_461_b : _GEN_17800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17802 = 10'h1ce == r_count_23_io_out ? io_r_462_b : _GEN_17801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17803 = 10'h1cf == r_count_23_io_out ? io_r_463_b : _GEN_17802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17804 = 10'h1d0 == r_count_23_io_out ? io_r_464_b : _GEN_17803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17805 = 10'h1d1 == r_count_23_io_out ? io_r_465_b : _GEN_17804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17806 = 10'h1d2 == r_count_23_io_out ? io_r_466_b : _GEN_17805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17807 = 10'h1d3 == r_count_23_io_out ? io_r_467_b : _GEN_17806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17808 = 10'h1d4 == r_count_23_io_out ? io_r_468_b : _GEN_17807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17809 = 10'h1d5 == r_count_23_io_out ? io_r_469_b : _GEN_17808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17810 = 10'h1d6 == r_count_23_io_out ? io_r_470_b : _GEN_17809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17811 = 10'h1d7 == r_count_23_io_out ? io_r_471_b : _GEN_17810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17812 = 10'h1d8 == r_count_23_io_out ? io_r_472_b : _GEN_17811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17813 = 10'h1d9 == r_count_23_io_out ? io_r_473_b : _GEN_17812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17814 = 10'h1da == r_count_23_io_out ? io_r_474_b : _GEN_17813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17815 = 10'h1db == r_count_23_io_out ? io_r_475_b : _GEN_17814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17816 = 10'h1dc == r_count_23_io_out ? io_r_476_b : _GEN_17815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17817 = 10'h1dd == r_count_23_io_out ? io_r_477_b : _GEN_17816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17818 = 10'h1de == r_count_23_io_out ? io_r_478_b : _GEN_17817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17819 = 10'h1df == r_count_23_io_out ? io_r_479_b : _GEN_17818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17820 = 10'h1e0 == r_count_23_io_out ? io_r_480_b : _GEN_17819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17821 = 10'h1e1 == r_count_23_io_out ? io_r_481_b : _GEN_17820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17822 = 10'h1e2 == r_count_23_io_out ? io_r_482_b : _GEN_17821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17823 = 10'h1e3 == r_count_23_io_out ? io_r_483_b : _GEN_17822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17824 = 10'h1e4 == r_count_23_io_out ? io_r_484_b : _GEN_17823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17825 = 10'h1e5 == r_count_23_io_out ? io_r_485_b : _GEN_17824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17826 = 10'h1e6 == r_count_23_io_out ? io_r_486_b : _GEN_17825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17827 = 10'h1e7 == r_count_23_io_out ? io_r_487_b : _GEN_17826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17828 = 10'h1e8 == r_count_23_io_out ? io_r_488_b : _GEN_17827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17829 = 10'h1e9 == r_count_23_io_out ? io_r_489_b : _GEN_17828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17830 = 10'h1ea == r_count_23_io_out ? io_r_490_b : _GEN_17829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17831 = 10'h1eb == r_count_23_io_out ? io_r_491_b : _GEN_17830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17832 = 10'h1ec == r_count_23_io_out ? io_r_492_b : _GEN_17831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17833 = 10'h1ed == r_count_23_io_out ? io_r_493_b : _GEN_17832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17834 = 10'h1ee == r_count_23_io_out ? io_r_494_b : _GEN_17833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17835 = 10'h1ef == r_count_23_io_out ? io_r_495_b : _GEN_17834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17836 = 10'h1f0 == r_count_23_io_out ? io_r_496_b : _GEN_17835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17837 = 10'h1f1 == r_count_23_io_out ? io_r_497_b : _GEN_17836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17838 = 10'h1f2 == r_count_23_io_out ? io_r_498_b : _GEN_17837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17839 = 10'h1f3 == r_count_23_io_out ? io_r_499_b : _GEN_17838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17840 = 10'h1f4 == r_count_23_io_out ? io_r_500_b : _GEN_17839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17841 = 10'h1f5 == r_count_23_io_out ? io_r_501_b : _GEN_17840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17842 = 10'h1f6 == r_count_23_io_out ? io_r_502_b : _GEN_17841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17843 = 10'h1f7 == r_count_23_io_out ? io_r_503_b : _GEN_17842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17844 = 10'h1f8 == r_count_23_io_out ? io_r_504_b : _GEN_17843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17845 = 10'h1f9 == r_count_23_io_out ? io_r_505_b : _GEN_17844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17846 = 10'h1fa == r_count_23_io_out ? io_r_506_b : _GEN_17845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17847 = 10'h1fb == r_count_23_io_out ? io_r_507_b : _GEN_17846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17848 = 10'h1fc == r_count_23_io_out ? io_r_508_b : _GEN_17847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17849 = 10'h1fd == r_count_23_io_out ? io_r_509_b : _GEN_17848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17850 = 10'h1fe == r_count_23_io_out ? io_r_510_b : _GEN_17849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17851 = 10'h1ff == r_count_23_io_out ? io_r_511_b : _GEN_17850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17852 = 10'h200 == r_count_23_io_out ? io_r_512_b : _GEN_17851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17853 = 10'h201 == r_count_23_io_out ? io_r_513_b : _GEN_17852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17854 = 10'h202 == r_count_23_io_out ? io_r_514_b : _GEN_17853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17855 = 10'h203 == r_count_23_io_out ? io_r_515_b : _GEN_17854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17856 = 10'h204 == r_count_23_io_out ? io_r_516_b : _GEN_17855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17857 = 10'h205 == r_count_23_io_out ? io_r_517_b : _GEN_17856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17858 = 10'h206 == r_count_23_io_out ? io_r_518_b : _GEN_17857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17859 = 10'h207 == r_count_23_io_out ? io_r_519_b : _GEN_17858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17860 = 10'h208 == r_count_23_io_out ? io_r_520_b : _GEN_17859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17861 = 10'h209 == r_count_23_io_out ? io_r_521_b : _GEN_17860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17862 = 10'h20a == r_count_23_io_out ? io_r_522_b : _GEN_17861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17863 = 10'h20b == r_count_23_io_out ? io_r_523_b : _GEN_17862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17864 = 10'h20c == r_count_23_io_out ? io_r_524_b : _GEN_17863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17865 = 10'h20d == r_count_23_io_out ? io_r_525_b : _GEN_17864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17866 = 10'h20e == r_count_23_io_out ? io_r_526_b : _GEN_17865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17867 = 10'h20f == r_count_23_io_out ? io_r_527_b : _GEN_17866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17868 = 10'h210 == r_count_23_io_out ? io_r_528_b : _GEN_17867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17869 = 10'h211 == r_count_23_io_out ? io_r_529_b : _GEN_17868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17870 = 10'h212 == r_count_23_io_out ? io_r_530_b : _GEN_17869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17871 = 10'h213 == r_count_23_io_out ? io_r_531_b : _GEN_17870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17872 = 10'h214 == r_count_23_io_out ? io_r_532_b : _GEN_17871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17873 = 10'h215 == r_count_23_io_out ? io_r_533_b : _GEN_17872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17874 = 10'h216 == r_count_23_io_out ? io_r_534_b : _GEN_17873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17875 = 10'h217 == r_count_23_io_out ? io_r_535_b : _GEN_17874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17876 = 10'h218 == r_count_23_io_out ? io_r_536_b : _GEN_17875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17877 = 10'h219 == r_count_23_io_out ? io_r_537_b : _GEN_17876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17878 = 10'h21a == r_count_23_io_out ? io_r_538_b : _GEN_17877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17879 = 10'h21b == r_count_23_io_out ? io_r_539_b : _GEN_17878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17880 = 10'h21c == r_count_23_io_out ? io_r_540_b : _GEN_17879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17881 = 10'h21d == r_count_23_io_out ? io_r_541_b : _GEN_17880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17882 = 10'h21e == r_count_23_io_out ? io_r_542_b : _GEN_17881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17883 = 10'h21f == r_count_23_io_out ? io_r_543_b : _GEN_17882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17884 = 10'h220 == r_count_23_io_out ? io_r_544_b : _GEN_17883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17885 = 10'h221 == r_count_23_io_out ? io_r_545_b : _GEN_17884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17886 = 10'h222 == r_count_23_io_out ? io_r_546_b : _GEN_17885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17887 = 10'h223 == r_count_23_io_out ? io_r_547_b : _GEN_17886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17888 = 10'h224 == r_count_23_io_out ? io_r_548_b : _GEN_17887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17889 = 10'h225 == r_count_23_io_out ? io_r_549_b : _GEN_17888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17890 = 10'h226 == r_count_23_io_out ? io_r_550_b : _GEN_17889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17891 = 10'h227 == r_count_23_io_out ? io_r_551_b : _GEN_17890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17892 = 10'h228 == r_count_23_io_out ? io_r_552_b : _GEN_17891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17893 = 10'h229 == r_count_23_io_out ? io_r_553_b : _GEN_17892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17894 = 10'h22a == r_count_23_io_out ? io_r_554_b : _GEN_17893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17895 = 10'h22b == r_count_23_io_out ? io_r_555_b : _GEN_17894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17896 = 10'h22c == r_count_23_io_out ? io_r_556_b : _GEN_17895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17897 = 10'h22d == r_count_23_io_out ? io_r_557_b : _GEN_17896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17898 = 10'h22e == r_count_23_io_out ? io_r_558_b : _GEN_17897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17899 = 10'h22f == r_count_23_io_out ? io_r_559_b : _GEN_17898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17900 = 10'h230 == r_count_23_io_out ? io_r_560_b : _GEN_17899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17901 = 10'h231 == r_count_23_io_out ? io_r_561_b : _GEN_17900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17902 = 10'h232 == r_count_23_io_out ? io_r_562_b : _GEN_17901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17903 = 10'h233 == r_count_23_io_out ? io_r_563_b : _GEN_17902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17904 = 10'h234 == r_count_23_io_out ? io_r_564_b : _GEN_17903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17905 = 10'h235 == r_count_23_io_out ? io_r_565_b : _GEN_17904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17906 = 10'h236 == r_count_23_io_out ? io_r_566_b : _GEN_17905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17907 = 10'h237 == r_count_23_io_out ? io_r_567_b : _GEN_17906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17908 = 10'h238 == r_count_23_io_out ? io_r_568_b : _GEN_17907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17909 = 10'h239 == r_count_23_io_out ? io_r_569_b : _GEN_17908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17910 = 10'h23a == r_count_23_io_out ? io_r_570_b : _GEN_17909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17911 = 10'h23b == r_count_23_io_out ? io_r_571_b : _GEN_17910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17912 = 10'h23c == r_count_23_io_out ? io_r_572_b : _GEN_17911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17913 = 10'h23d == r_count_23_io_out ? io_r_573_b : _GEN_17912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17914 = 10'h23e == r_count_23_io_out ? io_r_574_b : _GEN_17913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17915 = 10'h23f == r_count_23_io_out ? io_r_575_b : _GEN_17914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17916 = 10'h240 == r_count_23_io_out ? io_r_576_b : _GEN_17915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17917 = 10'h241 == r_count_23_io_out ? io_r_577_b : _GEN_17916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17918 = 10'h242 == r_count_23_io_out ? io_r_578_b : _GEN_17917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17919 = 10'h243 == r_count_23_io_out ? io_r_579_b : _GEN_17918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17920 = 10'h244 == r_count_23_io_out ? io_r_580_b : _GEN_17919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17921 = 10'h245 == r_count_23_io_out ? io_r_581_b : _GEN_17920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17922 = 10'h246 == r_count_23_io_out ? io_r_582_b : _GEN_17921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17923 = 10'h247 == r_count_23_io_out ? io_r_583_b : _GEN_17922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17924 = 10'h248 == r_count_23_io_out ? io_r_584_b : _GEN_17923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17925 = 10'h249 == r_count_23_io_out ? io_r_585_b : _GEN_17924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17926 = 10'h24a == r_count_23_io_out ? io_r_586_b : _GEN_17925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17927 = 10'h24b == r_count_23_io_out ? io_r_587_b : _GEN_17926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17928 = 10'h24c == r_count_23_io_out ? io_r_588_b : _GEN_17927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17929 = 10'h24d == r_count_23_io_out ? io_r_589_b : _GEN_17928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17930 = 10'h24e == r_count_23_io_out ? io_r_590_b : _GEN_17929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17931 = 10'h24f == r_count_23_io_out ? io_r_591_b : _GEN_17930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17932 = 10'h250 == r_count_23_io_out ? io_r_592_b : _GEN_17931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17933 = 10'h251 == r_count_23_io_out ? io_r_593_b : _GEN_17932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17934 = 10'h252 == r_count_23_io_out ? io_r_594_b : _GEN_17933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17935 = 10'h253 == r_count_23_io_out ? io_r_595_b : _GEN_17934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17936 = 10'h254 == r_count_23_io_out ? io_r_596_b : _GEN_17935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17937 = 10'h255 == r_count_23_io_out ? io_r_597_b : _GEN_17936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17938 = 10'h256 == r_count_23_io_out ? io_r_598_b : _GEN_17937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17939 = 10'h257 == r_count_23_io_out ? io_r_599_b : _GEN_17938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17940 = 10'h258 == r_count_23_io_out ? io_r_600_b : _GEN_17939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17941 = 10'h259 == r_count_23_io_out ? io_r_601_b : _GEN_17940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17942 = 10'h25a == r_count_23_io_out ? io_r_602_b : _GEN_17941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17943 = 10'h25b == r_count_23_io_out ? io_r_603_b : _GEN_17942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17944 = 10'h25c == r_count_23_io_out ? io_r_604_b : _GEN_17943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17945 = 10'h25d == r_count_23_io_out ? io_r_605_b : _GEN_17944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17946 = 10'h25e == r_count_23_io_out ? io_r_606_b : _GEN_17945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17947 = 10'h25f == r_count_23_io_out ? io_r_607_b : _GEN_17946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17948 = 10'h260 == r_count_23_io_out ? io_r_608_b : _GEN_17947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17949 = 10'h261 == r_count_23_io_out ? io_r_609_b : _GEN_17948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17950 = 10'h262 == r_count_23_io_out ? io_r_610_b : _GEN_17949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17951 = 10'h263 == r_count_23_io_out ? io_r_611_b : _GEN_17950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17952 = 10'h264 == r_count_23_io_out ? io_r_612_b : _GEN_17951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17953 = 10'h265 == r_count_23_io_out ? io_r_613_b : _GEN_17952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17954 = 10'h266 == r_count_23_io_out ? io_r_614_b : _GEN_17953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17955 = 10'h267 == r_count_23_io_out ? io_r_615_b : _GEN_17954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17956 = 10'h268 == r_count_23_io_out ? io_r_616_b : _GEN_17955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17957 = 10'h269 == r_count_23_io_out ? io_r_617_b : _GEN_17956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17958 = 10'h26a == r_count_23_io_out ? io_r_618_b : _GEN_17957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17959 = 10'h26b == r_count_23_io_out ? io_r_619_b : _GEN_17958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17960 = 10'h26c == r_count_23_io_out ? io_r_620_b : _GEN_17959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17961 = 10'h26d == r_count_23_io_out ? io_r_621_b : _GEN_17960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17962 = 10'h26e == r_count_23_io_out ? io_r_622_b : _GEN_17961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17963 = 10'h26f == r_count_23_io_out ? io_r_623_b : _GEN_17962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17964 = 10'h270 == r_count_23_io_out ? io_r_624_b : _GEN_17963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17965 = 10'h271 == r_count_23_io_out ? io_r_625_b : _GEN_17964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17966 = 10'h272 == r_count_23_io_out ? io_r_626_b : _GEN_17965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17967 = 10'h273 == r_count_23_io_out ? io_r_627_b : _GEN_17966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17968 = 10'h274 == r_count_23_io_out ? io_r_628_b : _GEN_17967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17969 = 10'h275 == r_count_23_io_out ? io_r_629_b : _GEN_17968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17970 = 10'h276 == r_count_23_io_out ? io_r_630_b : _GEN_17969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17971 = 10'h277 == r_count_23_io_out ? io_r_631_b : _GEN_17970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17972 = 10'h278 == r_count_23_io_out ? io_r_632_b : _GEN_17971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17973 = 10'h279 == r_count_23_io_out ? io_r_633_b : _GEN_17972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17974 = 10'h27a == r_count_23_io_out ? io_r_634_b : _GEN_17973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17975 = 10'h27b == r_count_23_io_out ? io_r_635_b : _GEN_17974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17976 = 10'h27c == r_count_23_io_out ? io_r_636_b : _GEN_17975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17977 = 10'h27d == r_count_23_io_out ? io_r_637_b : _GEN_17976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17978 = 10'h27e == r_count_23_io_out ? io_r_638_b : _GEN_17977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17979 = 10'h27f == r_count_23_io_out ? io_r_639_b : _GEN_17978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17980 = 10'h280 == r_count_23_io_out ? io_r_640_b : _GEN_17979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17981 = 10'h281 == r_count_23_io_out ? io_r_641_b : _GEN_17980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17982 = 10'h282 == r_count_23_io_out ? io_r_642_b : _GEN_17981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17983 = 10'h283 == r_count_23_io_out ? io_r_643_b : _GEN_17982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17984 = 10'h284 == r_count_23_io_out ? io_r_644_b : _GEN_17983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17985 = 10'h285 == r_count_23_io_out ? io_r_645_b : _GEN_17984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17986 = 10'h286 == r_count_23_io_out ? io_r_646_b : _GEN_17985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17987 = 10'h287 == r_count_23_io_out ? io_r_647_b : _GEN_17986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17988 = 10'h288 == r_count_23_io_out ? io_r_648_b : _GEN_17987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17989 = 10'h289 == r_count_23_io_out ? io_r_649_b : _GEN_17988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17990 = 10'h28a == r_count_23_io_out ? io_r_650_b : _GEN_17989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17991 = 10'h28b == r_count_23_io_out ? io_r_651_b : _GEN_17990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17992 = 10'h28c == r_count_23_io_out ? io_r_652_b : _GEN_17991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17993 = 10'h28d == r_count_23_io_out ? io_r_653_b : _GEN_17992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17994 = 10'h28e == r_count_23_io_out ? io_r_654_b : _GEN_17993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17995 = 10'h28f == r_count_23_io_out ? io_r_655_b : _GEN_17994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17996 = 10'h290 == r_count_23_io_out ? io_r_656_b : _GEN_17995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17997 = 10'h291 == r_count_23_io_out ? io_r_657_b : _GEN_17996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17998 = 10'h292 == r_count_23_io_out ? io_r_658_b : _GEN_17997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17999 = 10'h293 == r_count_23_io_out ? io_r_659_b : _GEN_17998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18000 = 10'h294 == r_count_23_io_out ? io_r_660_b : _GEN_17999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18001 = 10'h295 == r_count_23_io_out ? io_r_661_b : _GEN_18000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18002 = 10'h296 == r_count_23_io_out ? io_r_662_b : _GEN_18001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18003 = 10'h297 == r_count_23_io_out ? io_r_663_b : _GEN_18002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18004 = 10'h298 == r_count_23_io_out ? io_r_664_b : _GEN_18003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18005 = 10'h299 == r_count_23_io_out ? io_r_665_b : _GEN_18004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18006 = 10'h29a == r_count_23_io_out ? io_r_666_b : _GEN_18005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18007 = 10'h29b == r_count_23_io_out ? io_r_667_b : _GEN_18006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18008 = 10'h29c == r_count_23_io_out ? io_r_668_b : _GEN_18007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18009 = 10'h29d == r_count_23_io_out ? io_r_669_b : _GEN_18008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18010 = 10'h29e == r_count_23_io_out ? io_r_670_b : _GEN_18009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18011 = 10'h29f == r_count_23_io_out ? io_r_671_b : _GEN_18010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18012 = 10'h2a0 == r_count_23_io_out ? io_r_672_b : _GEN_18011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18013 = 10'h2a1 == r_count_23_io_out ? io_r_673_b : _GEN_18012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18014 = 10'h2a2 == r_count_23_io_out ? io_r_674_b : _GEN_18013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18015 = 10'h2a3 == r_count_23_io_out ? io_r_675_b : _GEN_18014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18016 = 10'h2a4 == r_count_23_io_out ? io_r_676_b : _GEN_18015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18017 = 10'h2a5 == r_count_23_io_out ? io_r_677_b : _GEN_18016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18018 = 10'h2a6 == r_count_23_io_out ? io_r_678_b : _GEN_18017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18019 = 10'h2a7 == r_count_23_io_out ? io_r_679_b : _GEN_18018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18020 = 10'h2a8 == r_count_23_io_out ? io_r_680_b : _GEN_18019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18021 = 10'h2a9 == r_count_23_io_out ? io_r_681_b : _GEN_18020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18022 = 10'h2aa == r_count_23_io_out ? io_r_682_b : _GEN_18021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18023 = 10'h2ab == r_count_23_io_out ? io_r_683_b : _GEN_18022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18024 = 10'h2ac == r_count_23_io_out ? io_r_684_b : _GEN_18023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18025 = 10'h2ad == r_count_23_io_out ? io_r_685_b : _GEN_18024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18026 = 10'h2ae == r_count_23_io_out ? io_r_686_b : _GEN_18025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18027 = 10'h2af == r_count_23_io_out ? io_r_687_b : _GEN_18026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18028 = 10'h2b0 == r_count_23_io_out ? io_r_688_b : _GEN_18027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18029 = 10'h2b1 == r_count_23_io_out ? io_r_689_b : _GEN_18028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18030 = 10'h2b2 == r_count_23_io_out ? io_r_690_b : _GEN_18029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18031 = 10'h2b3 == r_count_23_io_out ? io_r_691_b : _GEN_18030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18032 = 10'h2b4 == r_count_23_io_out ? io_r_692_b : _GEN_18031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18033 = 10'h2b5 == r_count_23_io_out ? io_r_693_b : _GEN_18032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18034 = 10'h2b6 == r_count_23_io_out ? io_r_694_b : _GEN_18033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18035 = 10'h2b7 == r_count_23_io_out ? io_r_695_b : _GEN_18034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18036 = 10'h2b8 == r_count_23_io_out ? io_r_696_b : _GEN_18035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18037 = 10'h2b9 == r_count_23_io_out ? io_r_697_b : _GEN_18036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18038 = 10'h2ba == r_count_23_io_out ? io_r_698_b : _GEN_18037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18039 = 10'h2bb == r_count_23_io_out ? io_r_699_b : _GEN_18038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18040 = 10'h2bc == r_count_23_io_out ? io_r_700_b : _GEN_18039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18041 = 10'h2bd == r_count_23_io_out ? io_r_701_b : _GEN_18040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18042 = 10'h2be == r_count_23_io_out ? io_r_702_b : _GEN_18041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18043 = 10'h2bf == r_count_23_io_out ? io_r_703_b : _GEN_18042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18044 = 10'h2c0 == r_count_23_io_out ? io_r_704_b : _GEN_18043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18045 = 10'h2c1 == r_count_23_io_out ? io_r_705_b : _GEN_18044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18046 = 10'h2c2 == r_count_23_io_out ? io_r_706_b : _GEN_18045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18047 = 10'h2c3 == r_count_23_io_out ? io_r_707_b : _GEN_18046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18048 = 10'h2c4 == r_count_23_io_out ? io_r_708_b : _GEN_18047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18049 = 10'h2c5 == r_count_23_io_out ? io_r_709_b : _GEN_18048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18050 = 10'h2c6 == r_count_23_io_out ? io_r_710_b : _GEN_18049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18051 = 10'h2c7 == r_count_23_io_out ? io_r_711_b : _GEN_18050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18052 = 10'h2c8 == r_count_23_io_out ? io_r_712_b : _GEN_18051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18053 = 10'h2c9 == r_count_23_io_out ? io_r_713_b : _GEN_18052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18054 = 10'h2ca == r_count_23_io_out ? io_r_714_b : _GEN_18053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18055 = 10'h2cb == r_count_23_io_out ? io_r_715_b : _GEN_18054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18056 = 10'h2cc == r_count_23_io_out ? io_r_716_b : _GEN_18055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18057 = 10'h2cd == r_count_23_io_out ? io_r_717_b : _GEN_18056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18058 = 10'h2ce == r_count_23_io_out ? io_r_718_b : _GEN_18057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18059 = 10'h2cf == r_count_23_io_out ? io_r_719_b : _GEN_18058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18060 = 10'h2d0 == r_count_23_io_out ? io_r_720_b : _GEN_18059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18061 = 10'h2d1 == r_count_23_io_out ? io_r_721_b : _GEN_18060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18062 = 10'h2d2 == r_count_23_io_out ? io_r_722_b : _GEN_18061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18063 = 10'h2d3 == r_count_23_io_out ? io_r_723_b : _GEN_18062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18064 = 10'h2d4 == r_count_23_io_out ? io_r_724_b : _GEN_18063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18065 = 10'h2d5 == r_count_23_io_out ? io_r_725_b : _GEN_18064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18066 = 10'h2d6 == r_count_23_io_out ? io_r_726_b : _GEN_18065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18067 = 10'h2d7 == r_count_23_io_out ? io_r_727_b : _GEN_18066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18068 = 10'h2d8 == r_count_23_io_out ? io_r_728_b : _GEN_18067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18069 = 10'h2d9 == r_count_23_io_out ? io_r_729_b : _GEN_18068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18070 = 10'h2da == r_count_23_io_out ? io_r_730_b : _GEN_18069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18071 = 10'h2db == r_count_23_io_out ? io_r_731_b : _GEN_18070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18072 = 10'h2dc == r_count_23_io_out ? io_r_732_b : _GEN_18071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18073 = 10'h2dd == r_count_23_io_out ? io_r_733_b : _GEN_18072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18074 = 10'h2de == r_count_23_io_out ? io_r_734_b : _GEN_18073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18075 = 10'h2df == r_count_23_io_out ? io_r_735_b : _GEN_18074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18076 = 10'h2e0 == r_count_23_io_out ? io_r_736_b : _GEN_18075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18077 = 10'h2e1 == r_count_23_io_out ? io_r_737_b : _GEN_18076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18078 = 10'h2e2 == r_count_23_io_out ? io_r_738_b : _GEN_18077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18079 = 10'h2e3 == r_count_23_io_out ? io_r_739_b : _GEN_18078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18080 = 10'h2e4 == r_count_23_io_out ? io_r_740_b : _GEN_18079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18081 = 10'h2e5 == r_count_23_io_out ? io_r_741_b : _GEN_18080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18082 = 10'h2e6 == r_count_23_io_out ? io_r_742_b : _GEN_18081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18083 = 10'h2e7 == r_count_23_io_out ? io_r_743_b : _GEN_18082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18084 = 10'h2e8 == r_count_23_io_out ? io_r_744_b : _GEN_18083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18085 = 10'h2e9 == r_count_23_io_out ? io_r_745_b : _GEN_18084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18086 = 10'h2ea == r_count_23_io_out ? io_r_746_b : _GEN_18085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18087 = 10'h2eb == r_count_23_io_out ? io_r_747_b : _GEN_18086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18088 = 10'h2ec == r_count_23_io_out ? io_r_748_b : _GEN_18087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18091 = 10'h1 == r_count_24_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18092 = 10'h2 == r_count_24_io_out ? io_r_2_b : _GEN_18091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18093 = 10'h3 == r_count_24_io_out ? io_r_3_b : _GEN_18092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18094 = 10'h4 == r_count_24_io_out ? io_r_4_b : _GEN_18093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18095 = 10'h5 == r_count_24_io_out ? io_r_5_b : _GEN_18094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18096 = 10'h6 == r_count_24_io_out ? io_r_6_b : _GEN_18095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18097 = 10'h7 == r_count_24_io_out ? io_r_7_b : _GEN_18096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18098 = 10'h8 == r_count_24_io_out ? io_r_8_b : _GEN_18097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18099 = 10'h9 == r_count_24_io_out ? io_r_9_b : _GEN_18098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18100 = 10'ha == r_count_24_io_out ? io_r_10_b : _GEN_18099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18101 = 10'hb == r_count_24_io_out ? io_r_11_b : _GEN_18100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18102 = 10'hc == r_count_24_io_out ? io_r_12_b : _GEN_18101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18103 = 10'hd == r_count_24_io_out ? io_r_13_b : _GEN_18102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18104 = 10'he == r_count_24_io_out ? io_r_14_b : _GEN_18103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18105 = 10'hf == r_count_24_io_out ? io_r_15_b : _GEN_18104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18106 = 10'h10 == r_count_24_io_out ? io_r_16_b : _GEN_18105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18107 = 10'h11 == r_count_24_io_out ? io_r_17_b : _GEN_18106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18108 = 10'h12 == r_count_24_io_out ? io_r_18_b : _GEN_18107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18109 = 10'h13 == r_count_24_io_out ? io_r_19_b : _GEN_18108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18110 = 10'h14 == r_count_24_io_out ? io_r_20_b : _GEN_18109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18111 = 10'h15 == r_count_24_io_out ? io_r_21_b : _GEN_18110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18112 = 10'h16 == r_count_24_io_out ? io_r_22_b : _GEN_18111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18113 = 10'h17 == r_count_24_io_out ? io_r_23_b : _GEN_18112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18114 = 10'h18 == r_count_24_io_out ? io_r_24_b : _GEN_18113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18115 = 10'h19 == r_count_24_io_out ? io_r_25_b : _GEN_18114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18116 = 10'h1a == r_count_24_io_out ? io_r_26_b : _GEN_18115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18117 = 10'h1b == r_count_24_io_out ? io_r_27_b : _GEN_18116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18118 = 10'h1c == r_count_24_io_out ? io_r_28_b : _GEN_18117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18119 = 10'h1d == r_count_24_io_out ? io_r_29_b : _GEN_18118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18120 = 10'h1e == r_count_24_io_out ? io_r_30_b : _GEN_18119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18121 = 10'h1f == r_count_24_io_out ? io_r_31_b : _GEN_18120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18122 = 10'h20 == r_count_24_io_out ? io_r_32_b : _GEN_18121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18123 = 10'h21 == r_count_24_io_out ? io_r_33_b : _GEN_18122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18124 = 10'h22 == r_count_24_io_out ? io_r_34_b : _GEN_18123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18125 = 10'h23 == r_count_24_io_out ? io_r_35_b : _GEN_18124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18126 = 10'h24 == r_count_24_io_out ? io_r_36_b : _GEN_18125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18127 = 10'h25 == r_count_24_io_out ? io_r_37_b : _GEN_18126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18128 = 10'h26 == r_count_24_io_out ? io_r_38_b : _GEN_18127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18129 = 10'h27 == r_count_24_io_out ? io_r_39_b : _GEN_18128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18130 = 10'h28 == r_count_24_io_out ? io_r_40_b : _GEN_18129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18131 = 10'h29 == r_count_24_io_out ? io_r_41_b : _GEN_18130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18132 = 10'h2a == r_count_24_io_out ? io_r_42_b : _GEN_18131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18133 = 10'h2b == r_count_24_io_out ? io_r_43_b : _GEN_18132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18134 = 10'h2c == r_count_24_io_out ? io_r_44_b : _GEN_18133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18135 = 10'h2d == r_count_24_io_out ? io_r_45_b : _GEN_18134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18136 = 10'h2e == r_count_24_io_out ? io_r_46_b : _GEN_18135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18137 = 10'h2f == r_count_24_io_out ? io_r_47_b : _GEN_18136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18138 = 10'h30 == r_count_24_io_out ? io_r_48_b : _GEN_18137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18139 = 10'h31 == r_count_24_io_out ? io_r_49_b : _GEN_18138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18140 = 10'h32 == r_count_24_io_out ? io_r_50_b : _GEN_18139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18141 = 10'h33 == r_count_24_io_out ? io_r_51_b : _GEN_18140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18142 = 10'h34 == r_count_24_io_out ? io_r_52_b : _GEN_18141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18143 = 10'h35 == r_count_24_io_out ? io_r_53_b : _GEN_18142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18144 = 10'h36 == r_count_24_io_out ? io_r_54_b : _GEN_18143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18145 = 10'h37 == r_count_24_io_out ? io_r_55_b : _GEN_18144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18146 = 10'h38 == r_count_24_io_out ? io_r_56_b : _GEN_18145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18147 = 10'h39 == r_count_24_io_out ? io_r_57_b : _GEN_18146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18148 = 10'h3a == r_count_24_io_out ? io_r_58_b : _GEN_18147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18149 = 10'h3b == r_count_24_io_out ? io_r_59_b : _GEN_18148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18150 = 10'h3c == r_count_24_io_out ? io_r_60_b : _GEN_18149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18151 = 10'h3d == r_count_24_io_out ? io_r_61_b : _GEN_18150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18152 = 10'h3e == r_count_24_io_out ? io_r_62_b : _GEN_18151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18153 = 10'h3f == r_count_24_io_out ? io_r_63_b : _GEN_18152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18154 = 10'h40 == r_count_24_io_out ? io_r_64_b : _GEN_18153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18155 = 10'h41 == r_count_24_io_out ? io_r_65_b : _GEN_18154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18156 = 10'h42 == r_count_24_io_out ? io_r_66_b : _GEN_18155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18157 = 10'h43 == r_count_24_io_out ? io_r_67_b : _GEN_18156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18158 = 10'h44 == r_count_24_io_out ? io_r_68_b : _GEN_18157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18159 = 10'h45 == r_count_24_io_out ? io_r_69_b : _GEN_18158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18160 = 10'h46 == r_count_24_io_out ? io_r_70_b : _GEN_18159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18161 = 10'h47 == r_count_24_io_out ? io_r_71_b : _GEN_18160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18162 = 10'h48 == r_count_24_io_out ? io_r_72_b : _GEN_18161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18163 = 10'h49 == r_count_24_io_out ? io_r_73_b : _GEN_18162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18164 = 10'h4a == r_count_24_io_out ? io_r_74_b : _GEN_18163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18165 = 10'h4b == r_count_24_io_out ? io_r_75_b : _GEN_18164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18166 = 10'h4c == r_count_24_io_out ? io_r_76_b : _GEN_18165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18167 = 10'h4d == r_count_24_io_out ? io_r_77_b : _GEN_18166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18168 = 10'h4e == r_count_24_io_out ? io_r_78_b : _GEN_18167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18169 = 10'h4f == r_count_24_io_out ? io_r_79_b : _GEN_18168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18170 = 10'h50 == r_count_24_io_out ? io_r_80_b : _GEN_18169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18171 = 10'h51 == r_count_24_io_out ? io_r_81_b : _GEN_18170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18172 = 10'h52 == r_count_24_io_out ? io_r_82_b : _GEN_18171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18173 = 10'h53 == r_count_24_io_out ? io_r_83_b : _GEN_18172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18174 = 10'h54 == r_count_24_io_out ? io_r_84_b : _GEN_18173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18175 = 10'h55 == r_count_24_io_out ? io_r_85_b : _GEN_18174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18176 = 10'h56 == r_count_24_io_out ? io_r_86_b : _GEN_18175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18177 = 10'h57 == r_count_24_io_out ? io_r_87_b : _GEN_18176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18178 = 10'h58 == r_count_24_io_out ? io_r_88_b : _GEN_18177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18179 = 10'h59 == r_count_24_io_out ? io_r_89_b : _GEN_18178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18180 = 10'h5a == r_count_24_io_out ? io_r_90_b : _GEN_18179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18181 = 10'h5b == r_count_24_io_out ? io_r_91_b : _GEN_18180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18182 = 10'h5c == r_count_24_io_out ? io_r_92_b : _GEN_18181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18183 = 10'h5d == r_count_24_io_out ? io_r_93_b : _GEN_18182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18184 = 10'h5e == r_count_24_io_out ? io_r_94_b : _GEN_18183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18185 = 10'h5f == r_count_24_io_out ? io_r_95_b : _GEN_18184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18186 = 10'h60 == r_count_24_io_out ? io_r_96_b : _GEN_18185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18187 = 10'h61 == r_count_24_io_out ? io_r_97_b : _GEN_18186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18188 = 10'h62 == r_count_24_io_out ? io_r_98_b : _GEN_18187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18189 = 10'h63 == r_count_24_io_out ? io_r_99_b : _GEN_18188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18190 = 10'h64 == r_count_24_io_out ? io_r_100_b : _GEN_18189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18191 = 10'h65 == r_count_24_io_out ? io_r_101_b : _GEN_18190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18192 = 10'h66 == r_count_24_io_out ? io_r_102_b : _GEN_18191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18193 = 10'h67 == r_count_24_io_out ? io_r_103_b : _GEN_18192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18194 = 10'h68 == r_count_24_io_out ? io_r_104_b : _GEN_18193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18195 = 10'h69 == r_count_24_io_out ? io_r_105_b : _GEN_18194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18196 = 10'h6a == r_count_24_io_out ? io_r_106_b : _GEN_18195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18197 = 10'h6b == r_count_24_io_out ? io_r_107_b : _GEN_18196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18198 = 10'h6c == r_count_24_io_out ? io_r_108_b : _GEN_18197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18199 = 10'h6d == r_count_24_io_out ? io_r_109_b : _GEN_18198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18200 = 10'h6e == r_count_24_io_out ? io_r_110_b : _GEN_18199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18201 = 10'h6f == r_count_24_io_out ? io_r_111_b : _GEN_18200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18202 = 10'h70 == r_count_24_io_out ? io_r_112_b : _GEN_18201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18203 = 10'h71 == r_count_24_io_out ? io_r_113_b : _GEN_18202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18204 = 10'h72 == r_count_24_io_out ? io_r_114_b : _GEN_18203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18205 = 10'h73 == r_count_24_io_out ? io_r_115_b : _GEN_18204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18206 = 10'h74 == r_count_24_io_out ? io_r_116_b : _GEN_18205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18207 = 10'h75 == r_count_24_io_out ? io_r_117_b : _GEN_18206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18208 = 10'h76 == r_count_24_io_out ? io_r_118_b : _GEN_18207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18209 = 10'h77 == r_count_24_io_out ? io_r_119_b : _GEN_18208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18210 = 10'h78 == r_count_24_io_out ? io_r_120_b : _GEN_18209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18211 = 10'h79 == r_count_24_io_out ? io_r_121_b : _GEN_18210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18212 = 10'h7a == r_count_24_io_out ? io_r_122_b : _GEN_18211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18213 = 10'h7b == r_count_24_io_out ? io_r_123_b : _GEN_18212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18214 = 10'h7c == r_count_24_io_out ? io_r_124_b : _GEN_18213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18215 = 10'h7d == r_count_24_io_out ? io_r_125_b : _GEN_18214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18216 = 10'h7e == r_count_24_io_out ? io_r_126_b : _GEN_18215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18217 = 10'h7f == r_count_24_io_out ? io_r_127_b : _GEN_18216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18218 = 10'h80 == r_count_24_io_out ? io_r_128_b : _GEN_18217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18219 = 10'h81 == r_count_24_io_out ? io_r_129_b : _GEN_18218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18220 = 10'h82 == r_count_24_io_out ? io_r_130_b : _GEN_18219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18221 = 10'h83 == r_count_24_io_out ? io_r_131_b : _GEN_18220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18222 = 10'h84 == r_count_24_io_out ? io_r_132_b : _GEN_18221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18223 = 10'h85 == r_count_24_io_out ? io_r_133_b : _GEN_18222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18224 = 10'h86 == r_count_24_io_out ? io_r_134_b : _GEN_18223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18225 = 10'h87 == r_count_24_io_out ? io_r_135_b : _GEN_18224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18226 = 10'h88 == r_count_24_io_out ? io_r_136_b : _GEN_18225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18227 = 10'h89 == r_count_24_io_out ? io_r_137_b : _GEN_18226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18228 = 10'h8a == r_count_24_io_out ? io_r_138_b : _GEN_18227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18229 = 10'h8b == r_count_24_io_out ? io_r_139_b : _GEN_18228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18230 = 10'h8c == r_count_24_io_out ? io_r_140_b : _GEN_18229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18231 = 10'h8d == r_count_24_io_out ? io_r_141_b : _GEN_18230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18232 = 10'h8e == r_count_24_io_out ? io_r_142_b : _GEN_18231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18233 = 10'h8f == r_count_24_io_out ? io_r_143_b : _GEN_18232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18234 = 10'h90 == r_count_24_io_out ? io_r_144_b : _GEN_18233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18235 = 10'h91 == r_count_24_io_out ? io_r_145_b : _GEN_18234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18236 = 10'h92 == r_count_24_io_out ? io_r_146_b : _GEN_18235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18237 = 10'h93 == r_count_24_io_out ? io_r_147_b : _GEN_18236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18238 = 10'h94 == r_count_24_io_out ? io_r_148_b : _GEN_18237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18239 = 10'h95 == r_count_24_io_out ? io_r_149_b : _GEN_18238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18240 = 10'h96 == r_count_24_io_out ? io_r_150_b : _GEN_18239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18241 = 10'h97 == r_count_24_io_out ? io_r_151_b : _GEN_18240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18242 = 10'h98 == r_count_24_io_out ? io_r_152_b : _GEN_18241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18243 = 10'h99 == r_count_24_io_out ? io_r_153_b : _GEN_18242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18244 = 10'h9a == r_count_24_io_out ? io_r_154_b : _GEN_18243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18245 = 10'h9b == r_count_24_io_out ? io_r_155_b : _GEN_18244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18246 = 10'h9c == r_count_24_io_out ? io_r_156_b : _GEN_18245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18247 = 10'h9d == r_count_24_io_out ? io_r_157_b : _GEN_18246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18248 = 10'h9e == r_count_24_io_out ? io_r_158_b : _GEN_18247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18249 = 10'h9f == r_count_24_io_out ? io_r_159_b : _GEN_18248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18250 = 10'ha0 == r_count_24_io_out ? io_r_160_b : _GEN_18249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18251 = 10'ha1 == r_count_24_io_out ? io_r_161_b : _GEN_18250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18252 = 10'ha2 == r_count_24_io_out ? io_r_162_b : _GEN_18251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18253 = 10'ha3 == r_count_24_io_out ? io_r_163_b : _GEN_18252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18254 = 10'ha4 == r_count_24_io_out ? io_r_164_b : _GEN_18253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18255 = 10'ha5 == r_count_24_io_out ? io_r_165_b : _GEN_18254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18256 = 10'ha6 == r_count_24_io_out ? io_r_166_b : _GEN_18255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18257 = 10'ha7 == r_count_24_io_out ? io_r_167_b : _GEN_18256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18258 = 10'ha8 == r_count_24_io_out ? io_r_168_b : _GEN_18257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18259 = 10'ha9 == r_count_24_io_out ? io_r_169_b : _GEN_18258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18260 = 10'haa == r_count_24_io_out ? io_r_170_b : _GEN_18259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18261 = 10'hab == r_count_24_io_out ? io_r_171_b : _GEN_18260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18262 = 10'hac == r_count_24_io_out ? io_r_172_b : _GEN_18261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18263 = 10'had == r_count_24_io_out ? io_r_173_b : _GEN_18262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18264 = 10'hae == r_count_24_io_out ? io_r_174_b : _GEN_18263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18265 = 10'haf == r_count_24_io_out ? io_r_175_b : _GEN_18264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18266 = 10'hb0 == r_count_24_io_out ? io_r_176_b : _GEN_18265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18267 = 10'hb1 == r_count_24_io_out ? io_r_177_b : _GEN_18266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18268 = 10'hb2 == r_count_24_io_out ? io_r_178_b : _GEN_18267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18269 = 10'hb3 == r_count_24_io_out ? io_r_179_b : _GEN_18268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18270 = 10'hb4 == r_count_24_io_out ? io_r_180_b : _GEN_18269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18271 = 10'hb5 == r_count_24_io_out ? io_r_181_b : _GEN_18270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18272 = 10'hb6 == r_count_24_io_out ? io_r_182_b : _GEN_18271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18273 = 10'hb7 == r_count_24_io_out ? io_r_183_b : _GEN_18272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18274 = 10'hb8 == r_count_24_io_out ? io_r_184_b : _GEN_18273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18275 = 10'hb9 == r_count_24_io_out ? io_r_185_b : _GEN_18274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18276 = 10'hba == r_count_24_io_out ? io_r_186_b : _GEN_18275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18277 = 10'hbb == r_count_24_io_out ? io_r_187_b : _GEN_18276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18278 = 10'hbc == r_count_24_io_out ? io_r_188_b : _GEN_18277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18279 = 10'hbd == r_count_24_io_out ? io_r_189_b : _GEN_18278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18280 = 10'hbe == r_count_24_io_out ? io_r_190_b : _GEN_18279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18281 = 10'hbf == r_count_24_io_out ? io_r_191_b : _GEN_18280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18282 = 10'hc0 == r_count_24_io_out ? io_r_192_b : _GEN_18281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18283 = 10'hc1 == r_count_24_io_out ? io_r_193_b : _GEN_18282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18284 = 10'hc2 == r_count_24_io_out ? io_r_194_b : _GEN_18283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18285 = 10'hc3 == r_count_24_io_out ? io_r_195_b : _GEN_18284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18286 = 10'hc4 == r_count_24_io_out ? io_r_196_b : _GEN_18285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18287 = 10'hc5 == r_count_24_io_out ? io_r_197_b : _GEN_18286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18288 = 10'hc6 == r_count_24_io_out ? io_r_198_b : _GEN_18287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18289 = 10'hc7 == r_count_24_io_out ? io_r_199_b : _GEN_18288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18290 = 10'hc8 == r_count_24_io_out ? io_r_200_b : _GEN_18289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18291 = 10'hc9 == r_count_24_io_out ? io_r_201_b : _GEN_18290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18292 = 10'hca == r_count_24_io_out ? io_r_202_b : _GEN_18291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18293 = 10'hcb == r_count_24_io_out ? io_r_203_b : _GEN_18292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18294 = 10'hcc == r_count_24_io_out ? io_r_204_b : _GEN_18293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18295 = 10'hcd == r_count_24_io_out ? io_r_205_b : _GEN_18294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18296 = 10'hce == r_count_24_io_out ? io_r_206_b : _GEN_18295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18297 = 10'hcf == r_count_24_io_out ? io_r_207_b : _GEN_18296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18298 = 10'hd0 == r_count_24_io_out ? io_r_208_b : _GEN_18297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18299 = 10'hd1 == r_count_24_io_out ? io_r_209_b : _GEN_18298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18300 = 10'hd2 == r_count_24_io_out ? io_r_210_b : _GEN_18299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18301 = 10'hd3 == r_count_24_io_out ? io_r_211_b : _GEN_18300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18302 = 10'hd4 == r_count_24_io_out ? io_r_212_b : _GEN_18301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18303 = 10'hd5 == r_count_24_io_out ? io_r_213_b : _GEN_18302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18304 = 10'hd6 == r_count_24_io_out ? io_r_214_b : _GEN_18303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18305 = 10'hd7 == r_count_24_io_out ? io_r_215_b : _GEN_18304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18306 = 10'hd8 == r_count_24_io_out ? io_r_216_b : _GEN_18305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18307 = 10'hd9 == r_count_24_io_out ? io_r_217_b : _GEN_18306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18308 = 10'hda == r_count_24_io_out ? io_r_218_b : _GEN_18307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18309 = 10'hdb == r_count_24_io_out ? io_r_219_b : _GEN_18308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18310 = 10'hdc == r_count_24_io_out ? io_r_220_b : _GEN_18309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18311 = 10'hdd == r_count_24_io_out ? io_r_221_b : _GEN_18310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18312 = 10'hde == r_count_24_io_out ? io_r_222_b : _GEN_18311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18313 = 10'hdf == r_count_24_io_out ? io_r_223_b : _GEN_18312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18314 = 10'he0 == r_count_24_io_out ? io_r_224_b : _GEN_18313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18315 = 10'he1 == r_count_24_io_out ? io_r_225_b : _GEN_18314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18316 = 10'he2 == r_count_24_io_out ? io_r_226_b : _GEN_18315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18317 = 10'he3 == r_count_24_io_out ? io_r_227_b : _GEN_18316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18318 = 10'he4 == r_count_24_io_out ? io_r_228_b : _GEN_18317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18319 = 10'he5 == r_count_24_io_out ? io_r_229_b : _GEN_18318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18320 = 10'he6 == r_count_24_io_out ? io_r_230_b : _GEN_18319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18321 = 10'he7 == r_count_24_io_out ? io_r_231_b : _GEN_18320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18322 = 10'he8 == r_count_24_io_out ? io_r_232_b : _GEN_18321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18323 = 10'he9 == r_count_24_io_out ? io_r_233_b : _GEN_18322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18324 = 10'hea == r_count_24_io_out ? io_r_234_b : _GEN_18323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18325 = 10'heb == r_count_24_io_out ? io_r_235_b : _GEN_18324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18326 = 10'hec == r_count_24_io_out ? io_r_236_b : _GEN_18325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18327 = 10'hed == r_count_24_io_out ? io_r_237_b : _GEN_18326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18328 = 10'hee == r_count_24_io_out ? io_r_238_b : _GEN_18327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18329 = 10'hef == r_count_24_io_out ? io_r_239_b : _GEN_18328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18330 = 10'hf0 == r_count_24_io_out ? io_r_240_b : _GEN_18329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18331 = 10'hf1 == r_count_24_io_out ? io_r_241_b : _GEN_18330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18332 = 10'hf2 == r_count_24_io_out ? io_r_242_b : _GEN_18331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18333 = 10'hf3 == r_count_24_io_out ? io_r_243_b : _GEN_18332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18334 = 10'hf4 == r_count_24_io_out ? io_r_244_b : _GEN_18333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18335 = 10'hf5 == r_count_24_io_out ? io_r_245_b : _GEN_18334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18336 = 10'hf6 == r_count_24_io_out ? io_r_246_b : _GEN_18335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18337 = 10'hf7 == r_count_24_io_out ? io_r_247_b : _GEN_18336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18338 = 10'hf8 == r_count_24_io_out ? io_r_248_b : _GEN_18337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18339 = 10'hf9 == r_count_24_io_out ? io_r_249_b : _GEN_18338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18340 = 10'hfa == r_count_24_io_out ? io_r_250_b : _GEN_18339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18341 = 10'hfb == r_count_24_io_out ? io_r_251_b : _GEN_18340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18342 = 10'hfc == r_count_24_io_out ? io_r_252_b : _GEN_18341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18343 = 10'hfd == r_count_24_io_out ? io_r_253_b : _GEN_18342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18344 = 10'hfe == r_count_24_io_out ? io_r_254_b : _GEN_18343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18345 = 10'hff == r_count_24_io_out ? io_r_255_b : _GEN_18344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18346 = 10'h100 == r_count_24_io_out ? io_r_256_b : _GEN_18345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18347 = 10'h101 == r_count_24_io_out ? io_r_257_b : _GEN_18346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18348 = 10'h102 == r_count_24_io_out ? io_r_258_b : _GEN_18347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18349 = 10'h103 == r_count_24_io_out ? io_r_259_b : _GEN_18348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18350 = 10'h104 == r_count_24_io_out ? io_r_260_b : _GEN_18349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18351 = 10'h105 == r_count_24_io_out ? io_r_261_b : _GEN_18350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18352 = 10'h106 == r_count_24_io_out ? io_r_262_b : _GEN_18351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18353 = 10'h107 == r_count_24_io_out ? io_r_263_b : _GEN_18352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18354 = 10'h108 == r_count_24_io_out ? io_r_264_b : _GEN_18353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18355 = 10'h109 == r_count_24_io_out ? io_r_265_b : _GEN_18354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18356 = 10'h10a == r_count_24_io_out ? io_r_266_b : _GEN_18355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18357 = 10'h10b == r_count_24_io_out ? io_r_267_b : _GEN_18356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18358 = 10'h10c == r_count_24_io_out ? io_r_268_b : _GEN_18357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18359 = 10'h10d == r_count_24_io_out ? io_r_269_b : _GEN_18358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18360 = 10'h10e == r_count_24_io_out ? io_r_270_b : _GEN_18359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18361 = 10'h10f == r_count_24_io_out ? io_r_271_b : _GEN_18360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18362 = 10'h110 == r_count_24_io_out ? io_r_272_b : _GEN_18361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18363 = 10'h111 == r_count_24_io_out ? io_r_273_b : _GEN_18362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18364 = 10'h112 == r_count_24_io_out ? io_r_274_b : _GEN_18363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18365 = 10'h113 == r_count_24_io_out ? io_r_275_b : _GEN_18364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18366 = 10'h114 == r_count_24_io_out ? io_r_276_b : _GEN_18365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18367 = 10'h115 == r_count_24_io_out ? io_r_277_b : _GEN_18366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18368 = 10'h116 == r_count_24_io_out ? io_r_278_b : _GEN_18367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18369 = 10'h117 == r_count_24_io_out ? io_r_279_b : _GEN_18368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18370 = 10'h118 == r_count_24_io_out ? io_r_280_b : _GEN_18369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18371 = 10'h119 == r_count_24_io_out ? io_r_281_b : _GEN_18370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18372 = 10'h11a == r_count_24_io_out ? io_r_282_b : _GEN_18371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18373 = 10'h11b == r_count_24_io_out ? io_r_283_b : _GEN_18372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18374 = 10'h11c == r_count_24_io_out ? io_r_284_b : _GEN_18373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18375 = 10'h11d == r_count_24_io_out ? io_r_285_b : _GEN_18374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18376 = 10'h11e == r_count_24_io_out ? io_r_286_b : _GEN_18375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18377 = 10'h11f == r_count_24_io_out ? io_r_287_b : _GEN_18376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18378 = 10'h120 == r_count_24_io_out ? io_r_288_b : _GEN_18377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18379 = 10'h121 == r_count_24_io_out ? io_r_289_b : _GEN_18378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18380 = 10'h122 == r_count_24_io_out ? io_r_290_b : _GEN_18379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18381 = 10'h123 == r_count_24_io_out ? io_r_291_b : _GEN_18380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18382 = 10'h124 == r_count_24_io_out ? io_r_292_b : _GEN_18381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18383 = 10'h125 == r_count_24_io_out ? io_r_293_b : _GEN_18382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18384 = 10'h126 == r_count_24_io_out ? io_r_294_b : _GEN_18383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18385 = 10'h127 == r_count_24_io_out ? io_r_295_b : _GEN_18384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18386 = 10'h128 == r_count_24_io_out ? io_r_296_b : _GEN_18385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18387 = 10'h129 == r_count_24_io_out ? io_r_297_b : _GEN_18386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18388 = 10'h12a == r_count_24_io_out ? io_r_298_b : _GEN_18387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18389 = 10'h12b == r_count_24_io_out ? io_r_299_b : _GEN_18388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18390 = 10'h12c == r_count_24_io_out ? io_r_300_b : _GEN_18389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18391 = 10'h12d == r_count_24_io_out ? io_r_301_b : _GEN_18390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18392 = 10'h12e == r_count_24_io_out ? io_r_302_b : _GEN_18391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18393 = 10'h12f == r_count_24_io_out ? io_r_303_b : _GEN_18392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18394 = 10'h130 == r_count_24_io_out ? io_r_304_b : _GEN_18393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18395 = 10'h131 == r_count_24_io_out ? io_r_305_b : _GEN_18394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18396 = 10'h132 == r_count_24_io_out ? io_r_306_b : _GEN_18395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18397 = 10'h133 == r_count_24_io_out ? io_r_307_b : _GEN_18396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18398 = 10'h134 == r_count_24_io_out ? io_r_308_b : _GEN_18397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18399 = 10'h135 == r_count_24_io_out ? io_r_309_b : _GEN_18398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18400 = 10'h136 == r_count_24_io_out ? io_r_310_b : _GEN_18399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18401 = 10'h137 == r_count_24_io_out ? io_r_311_b : _GEN_18400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18402 = 10'h138 == r_count_24_io_out ? io_r_312_b : _GEN_18401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18403 = 10'h139 == r_count_24_io_out ? io_r_313_b : _GEN_18402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18404 = 10'h13a == r_count_24_io_out ? io_r_314_b : _GEN_18403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18405 = 10'h13b == r_count_24_io_out ? io_r_315_b : _GEN_18404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18406 = 10'h13c == r_count_24_io_out ? io_r_316_b : _GEN_18405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18407 = 10'h13d == r_count_24_io_out ? io_r_317_b : _GEN_18406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18408 = 10'h13e == r_count_24_io_out ? io_r_318_b : _GEN_18407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18409 = 10'h13f == r_count_24_io_out ? io_r_319_b : _GEN_18408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18410 = 10'h140 == r_count_24_io_out ? io_r_320_b : _GEN_18409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18411 = 10'h141 == r_count_24_io_out ? io_r_321_b : _GEN_18410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18412 = 10'h142 == r_count_24_io_out ? io_r_322_b : _GEN_18411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18413 = 10'h143 == r_count_24_io_out ? io_r_323_b : _GEN_18412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18414 = 10'h144 == r_count_24_io_out ? io_r_324_b : _GEN_18413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18415 = 10'h145 == r_count_24_io_out ? io_r_325_b : _GEN_18414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18416 = 10'h146 == r_count_24_io_out ? io_r_326_b : _GEN_18415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18417 = 10'h147 == r_count_24_io_out ? io_r_327_b : _GEN_18416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18418 = 10'h148 == r_count_24_io_out ? io_r_328_b : _GEN_18417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18419 = 10'h149 == r_count_24_io_out ? io_r_329_b : _GEN_18418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18420 = 10'h14a == r_count_24_io_out ? io_r_330_b : _GEN_18419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18421 = 10'h14b == r_count_24_io_out ? io_r_331_b : _GEN_18420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18422 = 10'h14c == r_count_24_io_out ? io_r_332_b : _GEN_18421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18423 = 10'h14d == r_count_24_io_out ? io_r_333_b : _GEN_18422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18424 = 10'h14e == r_count_24_io_out ? io_r_334_b : _GEN_18423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18425 = 10'h14f == r_count_24_io_out ? io_r_335_b : _GEN_18424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18426 = 10'h150 == r_count_24_io_out ? io_r_336_b : _GEN_18425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18427 = 10'h151 == r_count_24_io_out ? io_r_337_b : _GEN_18426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18428 = 10'h152 == r_count_24_io_out ? io_r_338_b : _GEN_18427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18429 = 10'h153 == r_count_24_io_out ? io_r_339_b : _GEN_18428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18430 = 10'h154 == r_count_24_io_out ? io_r_340_b : _GEN_18429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18431 = 10'h155 == r_count_24_io_out ? io_r_341_b : _GEN_18430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18432 = 10'h156 == r_count_24_io_out ? io_r_342_b : _GEN_18431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18433 = 10'h157 == r_count_24_io_out ? io_r_343_b : _GEN_18432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18434 = 10'h158 == r_count_24_io_out ? io_r_344_b : _GEN_18433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18435 = 10'h159 == r_count_24_io_out ? io_r_345_b : _GEN_18434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18436 = 10'h15a == r_count_24_io_out ? io_r_346_b : _GEN_18435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18437 = 10'h15b == r_count_24_io_out ? io_r_347_b : _GEN_18436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18438 = 10'h15c == r_count_24_io_out ? io_r_348_b : _GEN_18437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18439 = 10'h15d == r_count_24_io_out ? io_r_349_b : _GEN_18438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18440 = 10'h15e == r_count_24_io_out ? io_r_350_b : _GEN_18439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18441 = 10'h15f == r_count_24_io_out ? io_r_351_b : _GEN_18440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18442 = 10'h160 == r_count_24_io_out ? io_r_352_b : _GEN_18441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18443 = 10'h161 == r_count_24_io_out ? io_r_353_b : _GEN_18442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18444 = 10'h162 == r_count_24_io_out ? io_r_354_b : _GEN_18443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18445 = 10'h163 == r_count_24_io_out ? io_r_355_b : _GEN_18444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18446 = 10'h164 == r_count_24_io_out ? io_r_356_b : _GEN_18445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18447 = 10'h165 == r_count_24_io_out ? io_r_357_b : _GEN_18446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18448 = 10'h166 == r_count_24_io_out ? io_r_358_b : _GEN_18447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18449 = 10'h167 == r_count_24_io_out ? io_r_359_b : _GEN_18448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18450 = 10'h168 == r_count_24_io_out ? io_r_360_b : _GEN_18449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18451 = 10'h169 == r_count_24_io_out ? io_r_361_b : _GEN_18450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18452 = 10'h16a == r_count_24_io_out ? io_r_362_b : _GEN_18451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18453 = 10'h16b == r_count_24_io_out ? io_r_363_b : _GEN_18452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18454 = 10'h16c == r_count_24_io_out ? io_r_364_b : _GEN_18453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18455 = 10'h16d == r_count_24_io_out ? io_r_365_b : _GEN_18454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18456 = 10'h16e == r_count_24_io_out ? io_r_366_b : _GEN_18455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18457 = 10'h16f == r_count_24_io_out ? io_r_367_b : _GEN_18456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18458 = 10'h170 == r_count_24_io_out ? io_r_368_b : _GEN_18457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18459 = 10'h171 == r_count_24_io_out ? io_r_369_b : _GEN_18458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18460 = 10'h172 == r_count_24_io_out ? io_r_370_b : _GEN_18459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18461 = 10'h173 == r_count_24_io_out ? io_r_371_b : _GEN_18460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18462 = 10'h174 == r_count_24_io_out ? io_r_372_b : _GEN_18461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18463 = 10'h175 == r_count_24_io_out ? io_r_373_b : _GEN_18462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18464 = 10'h176 == r_count_24_io_out ? io_r_374_b : _GEN_18463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18465 = 10'h177 == r_count_24_io_out ? io_r_375_b : _GEN_18464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18466 = 10'h178 == r_count_24_io_out ? io_r_376_b : _GEN_18465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18467 = 10'h179 == r_count_24_io_out ? io_r_377_b : _GEN_18466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18468 = 10'h17a == r_count_24_io_out ? io_r_378_b : _GEN_18467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18469 = 10'h17b == r_count_24_io_out ? io_r_379_b : _GEN_18468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18470 = 10'h17c == r_count_24_io_out ? io_r_380_b : _GEN_18469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18471 = 10'h17d == r_count_24_io_out ? io_r_381_b : _GEN_18470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18472 = 10'h17e == r_count_24_io_out ? io_r_382_b : _GEN_18471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18473 = 10'h17f == r_count_24_io_out ? io_r_383_b : _GEN_18472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18474 = 10'h180 == r_count_24_io_out ? io_r_384_b : _GEN_18473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18475 = 10'h181 == r_count_24_io_out ? io_r_385_b : _GEN_18474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18476 = 10'h182 == r_count_24_io_out ? io_r_386_b : _GEN_18475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18477 = 10'h183 == r_count_24_io_out ? io_r_387_b : _GEN_18476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18478 = 10'h184 == r_count_24_io_out ? io_r_388_b : _GEN_18477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18479 = 10'h185 == r_count_24_io_out ? io_r_389_b : _GEN_18478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18480 = 10'h186 == r_count_24_io_out ? io_r_390_b : _GEN_18479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18481 = 10'h187 == r_count_24_io_out ? io_r_391_b : _GEN_18480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18482 = 10'h188 == r_count_24_io_out ? io_r_392_b : _GEN_18481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18483 = 10'h189 == r_count_24_io_out ? io_r_393_b : _GEN_18482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18484 = 10'h18a == r_count_24_io_out ? io_r_394_b : _GEN_18483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18485 = 10'h18b == r_count_24_io_out ? io_r_395_b : _GEN_18484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18486 = 10'h18c == r_count_24_io_out ? io_r_396_b : _GEN_18485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18487 = 10'h18d == r_count_24_io_out ? io_r_397_b : _GEN_18486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18488 = 10'h18e == r_count_24_io_out ? io_r_398_b : _GEN_18487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18489 = 10'h18f == r_count_24_io_out ? io_r_399_b : _GEN_18488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18490 = 10'h190 == r_count_24_io_out ? io_r_400_b : _GEN_18489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18491 = 10'h191 == r_count_24_io_out ? io_r_401_b : _GEN_18490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18492 = 10'h192 == r_count_24_io_out ? io_r_402_b : _GEN_18491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18493 = 10'h193 == r_count_24_io_out ? io_r_403_b : _GEN_18492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18494 = 10'h194 == r_count_24_io_out ? io_r_404_b : _GEN_18493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18495 = 10'h195 == r_count_24_io_out ? io_r_405_b : _GEN_18494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18496 = 10'h196 == r_count_24_io_out ? io_r_406_b : _GEN_18495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18497 = 10'h197 == r_count_24_io_out ? io_r_407_b : _GEN_18496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18498 = 10'h198 == r_count_24_io_out ? io_r_408_b : _GEN_18497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18499 = 10'h199 == r_count_24_io_out ? io_r_409_b : _GEN_18498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18500 = 10'h19a == r_count_24_io_out ? io_r_410_b : _GEN_18499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18501 = 10'h19b == r_count_24_io_out ? io_r_411_b : _GEN_18500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18502 = 10'h19c == r_count_24_io_out ? io_r_412_b : _GEN_18501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18503 = 10'h19d == r_count_24_io_out ? io_r_413_b : _GEN_18502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18504 = 10'h19e == r_count_24_io_out ? io_r_414_b : _GEN_18503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18505 = 10'h19f == r_count_24_io_out ? io_r_415_b : _GEN_18504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18506 = 10'h1a0 == r_count_24_io_out ? io_r_416_b : _GEN_18505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18507 = 10'h1a1 == r_count_24_io_out ? io_r_417_b : _GEN_18506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18508 = 10'h1a2 == r_count_24_io_out ? io_r_418_b : _GEN_18507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18509 = 10'h1a3 == r_count_24_io_out ? io_r_419_b : _GEN_18508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18510 = 10'h1a4 == r_count_24_io_out ? io_r_420_b : _GEN_18509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18511 = 10'h1a5 == r_count_24_io_out ? io_r_421_b : _GEN_18510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18512 = 10'h1a6 == r_count_24_io_out ? io_r_422_b : _GEN_18511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18513 = 10'h1a7 == r_count_24_io_out ? io_r_423_b : _GEN_18512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18514 = 10'h1a8 == r_count_24_io_out ? io_r_424_b : _GEN_18513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18515 = 10'h1a9 == r_count_24_io_out ? io_r_425_b : _GEN_18514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18516 = 10'h1aa == r_count_24_io_out ? io_r_426_b : _GEN_18515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18517 = 10'h1ab == r_count_24_io_out ? io_r_427_b : _GEN_18516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18518 = 10'h1ac == r_count_24_io_out ? io_r_428_b : _GEN_18517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18519 = 10'h1ad == r_count_24_io_out ? io_r_429_b : _GEN_18518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18520 = 10'h1ae == r_count_24_io_out ? io_r_430_b : _GEN_18519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18521 = 10'h1af == r_count_24_io_out ? io_r_431_b : _GEN_18520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18522 = 10'h1b0 == r_count_24_io_out ? io_r_432_b : _GEN_18521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18523 = 10'h1b1 == r_count_24_io_out ? io_r_433_b : _GEN_18522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18524 = 10'h1b2 == r_count_24_io_out ? io_r_434_b : _GEN_18523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18525 = 10'h1b3 == r_count_24_io_out ? io_r_435_b : _GEN_18524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18526 = 10'h1b4 == r_count_24_io_out ? io_r_436_b : _GEN_18525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18527 = 10'h1b5 == r_count_24_io_out ? io_r_437_b : _GEN_18526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18528 = 10'h1b6 == r_count_24_io_out ? io_r_438_b : _GEN_18527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18529 = 10'h1b7 == r_count_24_io_out ? io_r_439_b : _GEN_18528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18530 = 10'h1b8 == r_count_24_io_out ? io_r_440_b : _GEN_18529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18531 = 10'h1b9 == r_count_24_io_out ? io_r_441_b : _GEN_18530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18532 = 10'h1ba == r_count_24_io_out ? io_r_442_b : _GEN_18531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18533 = 10'h1bb == r_count_24_io_out ? io_r_443_b : _GEN_18532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18534 = 10'h1bc == r_count_24_io_out ? io_r_444_b : _GEN_18533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18535 = 10'h1bd == r_count_24_io_out ? io_r_445_b : _GEN_18534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18536 = 10'h1be == r_count_24_io_out ? io_r_446_b : _GEN_18535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18537 = 10'h1bf == r_count_24_io_out ? io_r_447_b : _GEN_18536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18538 = 10'h1c0 == r_count_24_io_out ? io_r_448_b : _GEN_18537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18539 = 10'h1c1 == r_count_24_io_out ? io_r_449_b : _GEN_18538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18540 = 10'h1c2 == r_count_24_io_out ? io_r_450_b : _GEN_18539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18541 = 10'h1c3 == r_count_24_io_out ? io_r_451_b : _GEN_18540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18542 = 10'h1c4 == r_count_24_io_out ? io_r_452_b : _GEN_18541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18543 = 10'h1c5 == r_count_24_io_out ? io_r_453_b : _GEN_18542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18544 = 10'h1c6 == r_count_24_io_out ? io_r_454_b : _GEN_18543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18545 = 10'h1c7 == r_count_24_io_out ? io_r_455_b : _GEN_18544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18546 = 10'h1c8 == r_count_24_io_out ? io_r_456_b : _GEN_18545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18547 = 10'h1c9 == r_count_24_io_out ? io_r_457_b : _GEN_18546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18548 = 10'h1ca == r_count_24_io_out ? io_r_458_b : _GEN_18547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18549 = 10'h1cb == r_count_24_io_out ? io_r_459_b : _GEN_18548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18550 = 10'h1cc == r_count_24_io_out ? io_r_460_b : _GEN_18549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18551 = 10'h1cd == r_count_24_io_out ? io_r_461_b : _GEN_18550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18552 = 10'h1ce == r_count_24_io_out ? io_r_462_b : _GEN_18551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18553 = 10'h1cf == r_count_24_io_out ? io_r_463_b : _GEN_18552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18554 = 10'h1d0 == r_count_24_io_out ? io_r_464_b : _GEN_18553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18555 = 10'h1d1 == r_count_24_io_out ? io_r_465_b : _GEN_18554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18556 = 10'h1d2 == r_count_24_io_out ? io_r_466_b : _GEN_18555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18557 = 10'h1d3 == r_count_24_io_out ? io_r_467_b : _GEN_18556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18558 = 10'h1d4 == r_count_24_io_out ? io_r_468_b : _GEN_18557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18559 = 10'h1d5 == r_count_24_io_out ? io_r_469_b : _GEN_18558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18560 = 10'h1d6 == r_count_24_io_out ? io_r_470_b : _GEN_18559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18561 = 10'h1d7 == r_count_24_io_out ? io_r_471_b : _GEN_18560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18562 = 10'h1d8 == r_count_24_io_out ? io_r_472_b : _GEN_18561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18563 = 10'h1d9 == r_count_24_io_out ? io_r_473_b : _GEN_18562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18564 = 10'h1da == r_count_24_io_out ? io_r_474_b : _GEN_18563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18565 = 10'h1db == r_count_24_io_out ? io_r_475_b : _GEN_18564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18566 = 10'h1dc == r_count_24_io_out ? io_r_476_b : _GEN_18565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18567 = 10'h1dd == r_count_24_io_out ? io_r_477_b : _GEN_18566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18568 = 10'h1de == r_count_24_io_out ? io_r_478_b : _GEN_18567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18569 = 10'h1df == r_count_24_io_out ? io_r_479_b : _GEN_18568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18570 = 10'h1e0 == r_count_24_io_out ? io_r_480_b : _GEN_18569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18571 = 10'h1e1 == r_count_24_io_out ? io_r_481_b : _GEN_18570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18572 = 10'h1e2 == r_count_24_io_out ? io_r_482_b : _GEN_18571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18573 = 10'h1e3 == r_count_24_io_out ? io_r_483_b : _GEN_18572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18574 = 10'h1e4 == r_count_24_io_out ? io_r_484_b : _GEN_18573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18575 = 10'h1e5 == r_count_24_io_out ? io_r_485_b : _GEN_18574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18576 = 10'h1e6 == r_count_24_io_out ? io_r_486_b : _GEN_18575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18577 = 10'h1e7 == r_count_24_io_out ? io_r_487_b : _GEN_18576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18578 = 10'h1e8 == r_count_24_io_out ? io_r_488_b : _GEN_18577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18579 = 10'h1e9 == r_count_24_io_out ? io_r_489_b : _GEN_18578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18580 = 10'h1ea == r_count_24_io_out ? io_r_490_b : _GEN_18579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18581 = 10'h1eb == r_count_24_io_out ? io_r_491_b : _GEN_18580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18582 = 10'h1ec == r_count_24_io_out ? io_r_492_b : _GEN_18581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18583 = 10'h1ed == r_count_24_io_out ? io_r_493_b : _GEN_18582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18584 = 10'h1ee == r_count_24_io_out ? io_r_494_b : _GEN_18583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18585 = 10'h1ef == r_count_24_io_out ? io_r_495_b : _GEN_18584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18586 = 10'h1f0 == r_count_24_io_out ? io_r_496_b : _GEN_18585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18587 = 10'h1f1 == r_count_24_io_out ? io_r_497_b : _GEN_18586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18588 = 10'h1f2 == r_count_24_io_out ? io_r_498_b : _GEN_18587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18589 = 10'h1f3 == r_count_24_io_out ? io_r_499_b : _GEN_18588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18590 = 10'h1f4 == r_count_24_io_out ? io_r_500_b : _GEN_18589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18591 = 10'h1f5 == r_count_24_io_out ? io_r_501_b : _GEN_18590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18592 = 10'h1f6 == r_count_24_io_out ? io_r_502_b : _GEN_18591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18593 = 10'h1f7 == r_count_24_io_out ? io_r_503_b : _GEN_18592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18594 = 10'h1f8 == r_count_24_io_out ? io_r_504_b : _GEN_18593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18595 = 10'h1f9 == r_count_24_io_out ? io_r_505_b : _GEN_18594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18596 = 10'h1fa == r_count_24_io_out ? io_r_506_b : _GEN_18595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18597 = 10'h1fb == r_count_24_io_out ? io_r_507_b : _GEN_18596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18598 = 10'h1fc == r_count_24_io_out ? io_r_508_b : _GEN_18597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18599 = 10'h1fd == r_count_24_io_out ? io_r_509_b : _GEN_18598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18600 = 10'h1fe == r_count_24_io_out ? io_r_510_b : _GEN_18599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18601 = 10'h1ff == r_count_24_io_out ? io_r_511_b : _GEN_18600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18602 = 10'h200 == r_count_24_io_out ? io_r_512_b : _GEN_18601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18603 = 10'h201 == r_count_24_io_out ? io_r_513_b : _GEN_18602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18604 = 10'h202 == r_count_24_io_out ? io_r_514_b : _GEN_18603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18605 = 10'h203 == r_count_24_io_out ? io_r_515_b : _GEN_18604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18606 = 10'h204 == r_count_24_io_out ? io_r_516_b : _GEN_18605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18607 = 10'h205 == r_count_24_io_out ? io_r_517_b : _GEN_18606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18608 = 10'h206 == r_count_24_io_out ? io_r_518_b : _GEN_18607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18609 = 10'h207 == r_count_24_io_out ? io_r_519_b : _GEN_18608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18610 = 10'h208 == r_count_24_io_out ? io_r_520_b : _GEN_18609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18611 = 10'h209 == r_count_24_io_out ? io_r_521_b : _GEN_18610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18612 = 10'h20a == r_count_24_io_out ? io_r_522_b : _GEN_18611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18613 = 10'h20b == r_count_24_io_out ? io_r_523_b : _GEN_18612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18614 = 10'h20c == r_count_24_io_out ? io_r_524_b : _GEN_18613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18615 = 10'h20d == r_count_24_io_out ? io_r_525_b : _GEN_18614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18616 = 10'h20e == r_count_24_io_out ? io_r_526_b : _GEN_18615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18617 = 10'h20f == r_count_24_io_out ? io_r_527_b : _GEN_18616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18618 = 10'h210 == r_count_24_io_out ? io_r_528_b : _GEN_18617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18619 = 10'h211 == r_count_24_io_out ? io_r_529_b : _GEN_18618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18620 = 10'h212 == r_count_24_io_out ? io_r_530_b : _GEN_18619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18621 = 10'h213 == r_count_24_io_out ? io_r_531_b : _GEN_18620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18622 = 10'h214 == r_count_24_io_out ? io_r_532_b : _GEN_18621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18623 = 10'h215 == r_count_24_io_out ? io_r_533_b : _GEN_18622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18624 = 10'h216 == r_count_24_io_out ? io_r_534_b : _GEN_18623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18625 = 10'h217 == r_count_24_io_out ? io_r_535_b : _GEN_18624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18626 = 10'h218 == r_count_24_io_out ? io_r_536_b : _GEN_18625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18627 = 10'h219 == r_count_24_io_out ? io_r_537_b : _GEN_18626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18628 = 10'h21a == r_count_24_io_out ? io_r_538_b : _GEN_18627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18629 = 10'h21b == r_count_24_io_out ? io_r_539_b : _GEN_18628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18630 = 10'h21c == r_count_24_io_out ? io_r_540_b : _GEN_18629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18631 = 10'h21d == r_count_24_io_out ? io_r_541_b : _GEN_18630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18632 = 10'h21e == r_count_24_io_out ? io_r_542_b : _GEN_18631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18633 = 10'h21f == r_count_24_io_out ? io_r_543_b : _GEN_18632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18634 = 10'h220 == r_count_24_io_out ? io_r_544_b : _GEN_18633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18635 = 10'h221 == r_count_24_io_out ? io_r_545_b : _GEN_18634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18636 = 10'h222 == r_count_24_io_out ? io_r_546_b : _GEN_18635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18637 = 10'h223 == r_count_24_io_out ? io_r_547_b : _GEN_18636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18638 = 10'h224 == r_count_24_io_out ? io_r_548_b : _GEN_18637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18639 = 10'h225 == r_count_24_io_out ? io_r_549_b : _GEN_18638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18640 = 10'h226 == r_count_24_io_out ? io_r_550_b : _GEN_18639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18641 = 10'h227 == r_count_24_io_out ? io_r_551_b : _GEN_18640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18642 = 10'h228 == r_count_24_io_out ? io_r_552_b : _GEN_18641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18643 = 10'h229 == r_count_24_io_out ? io_r_553_b : _GEN_18642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18644 = 10'h22a == r_count_24_io_out ? io_r_554_b : _GEN_18643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18645 = 10'h22b == r_count_24_io_out ? io_r_555_b : _GEN_18644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18646 = 10'h22c == r_count_24_io_out ? io_r_556_b : _GEN_18645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18647 = 10'h22d == r_count_24_io_out ? io_r_557_b : _GEN_18646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18648 = 10'h22e == r_count_24_io_out ? io_r_558_b : _GEN_18647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18649 = 10'h22f == r_count_24_io_out ? io_r_559_b : _GEN_18648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18650 = 10'h230 == r_count_24_io_out ? io_r_560_b : _GEN_18649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18651 = 10'h231 == r_count_24_io_out ? io_r_561_b : _GEN_18650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18652 = 10'h232 == r_count_24_io_out ? io_r_562_b : _GEN_18651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18653 = 10'h233 == r_count_24_io_out ? io_r_563_b : _GEN_18652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18654 = 10'h234 == r_count_24_io_out ? io_r_564_b : _GEN_18653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18655 = 10'h235 == r_count_24_io_out ? io_r_565_b : _GEN_18654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18656 = 10'h236 == r_count_24_io_out ? io_r_566_b : _GEN_18655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18657 = 10'h237 == r_count_24_io_out ? io_r_567_b : _GEN_18656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18658 = 10'h238 == r_count_24_io_out ? io_r_568_b : _GEN_18657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18659 = 10'h239 == r_count_24_io_out ? io_r_569_b : _GEN_18658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18660 = 10'h23a == r_count_24_io_out ? io_r_570_b : _GEN_18659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18661 = 10'h23b == r_count_24_io_out ? io_r_571_b : _GEN_18660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18662 = 10'h23c == r_count_24_io_out ? io_r_572_b : _GEN_18661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18663 = 10'h23d == r_count_24_io_out ? io_r_573_b : _GEN_18662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18664 = 10'h23e == r_count_24_io_out ? io_r_574_b : _GEN_18663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18665 = 10'h23f == r_count_24_io_out ? io_r_575_b : _GEN_18664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18666 = 10'h240 == r_count_24_io_out ? io_r_576_b : _GEN_18665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18667 = 10'h241 == r_count_24_io_out ? io_r_577_b : _GEN_18666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18668 = 10'h242 == r_count_24_io_out ? io_r_578_b : _GEN_18667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18669 = 10'h243 == r_count_24_io_out ? io_r_579_b : _GEN_18668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18670 = 10'h244 == r_count_24_io_out ? io_r_580_b : _GEN_18669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18671 = 10'h245 == r_count_24_io_out ? io_r_581_b : _GEN_18670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18672 = 10'h246 == r_count_24_io_out ? io_r_582_b : _GEN_18671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18673 = 10'h247 == r_count_24_io_out ? io_r_583_b : _GEN_18672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18674 = 10'h248 == r_count_24_io_out ? io_r_584_b : _GEN_18673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18675 = 10'h249 == r_count_24_io_out ? io_r_585_b : _GEN_18674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18676 = 10'h24a == r_count_24_io_out ? io_r_586_b : _GEN_18675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18677 = 10'h24b == r_count_24_io_out ? io_r_587_b : _GEN_18676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18678 = 10'h24c == r_count_24_io_out ? io_r_588_b : _GEN_18677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18679 = 10'h24d == r_count_24_io_out ? io_r_589_b : _GEN_18678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18680 = 10'h24e == r_count_24_io_out ? io_r_590_b : _GEN_18679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18681 = 10'h24f == r_count_24_io_out ? io_r_591_b : _GEN_18680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18682 = 10'h250 == r_count_24_io_out ? io_r_592_b : _GEN_18681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18683 = 10'h251 == r_count_24_io_out ? io_r_593_b : _GEN_18682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18684 = 10'h252 == r_count_24_io_out ? io_r_594_b : _GEN_18683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18685 = 10'h253 == r_count_24_io_out ? io_r_595_b : _GEN_18684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18686 = 10'h254 == r_count_24_io_out ? io_r_596_b : _GEN_18685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18687 = 10'h255 == r_count_24_io_out ? io_r_597_b : _GEN_18686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18688 = 10'h256 == r_count_24_io_out ? io_r_598_b : _GEN_18687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18689 = 10'h257 == r_count_24_io_out ? io_r_599_b : _GEN_18688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18690 = 10'h258 == r_count_24_io_out ? io_r_600_b : _GEN_18689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18691 = 10'h259 == r_count_24_io_out ? io_r_601_b : _GEN_18690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18692 = 10'h25a == r_count_24_io_out ? io_r_602_b : _GEN_18691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18693 = 10'h25b == r_count_24_io_out ? io_r_603_b : _GEN_18692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18694 = 10'h25c == r_count_24_io_out ? io_r_604_b : _GEN_18693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18695 = 10'h25d == r_count_24_io_out ? io_r_605_b : _GEN_18694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18696 = 10'h25e == r_count_24_io_out ? io_r_606_b : _GEN_18695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18697 = 10'h25f == r_count_24_io_out ? io_r_607_b : _GEN_18696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18698 = 10'h260 == r_count_24_io_out ? io_r_608_b : _GEN_18697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18699 = 10'h261 == r_count_24_io_out ? io_r_609_b : _GEN_18698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18700 = 10'h262 == r_count_24_io_out ? io_r_610_b : _GEN_18699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18701 = 10'h263 == r_count_24_io_out ? io_r_611_b : _GEN_18700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18702 = 10'h264 == r_count_24_io_out ? io_r_612_b : _GEN_18701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18703 = 10'h265 == r_count_24_io_out ? io_r_613_b : _GEN_18702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18704 = 10'h266 == r_count_24_io_out ? io_r_614_b : _GEN_18703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18705 = 10'h267 == r_count_24_io_out ? io_r_615_b : _GEN_18704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18706 = 10'h268 == r_count_24_io_out ? io_r_616_b : _GEN_18705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18707 = 10'h269 == r_count_24_io_out ? io_r_617_b : _GEN_18706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18708 = 10'h26a == r_count_24_io_out ? io_r_618_b : _GEN_18707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18709 = 10'h26b == r_count_24_io_out ? io_r_619_b : _GEN_18708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18710 = 10'h26c == r_count_24_io_out ? io_r_620_b : _GEN_18709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18711 = 10'h26d == r_count_24_io_out ? io_r_621_b : _GEN_18710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18712 = 10'h26e == r_count_24_io_out ? io_r_622_b : _GEN_18711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18713 = 10'h26f == r_count_24_io_out ? io_r_623_b : _GEN_18712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18714 = 10'h270 == r_count_24_io_out ? io_r_624_b : _GEN_18713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18715 = 10'h271 == r_count_24_io_out ? io_r_625_b : _GEN_18714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18716 = 10'h272 == r_count_24_io_out ? io_r_626_b : _GEN_18715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18717 = 10'h273 == r_count_24_io_out ? io_r_627_b : _GEN_18716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18718 = 10'h274 == r_count_24_io_out ? io_r_628_b : _GEN_18717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18719 = 10'h275 == r_count_24_io_out ? io_r_629_b : _GEN_18718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18720 = 10'h276 == r_count_24_io_out ? io_r_630_b : _GEN_18719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18721 = 10'h277 == r_count_24_io_out ? io_r_631_b : _GEN_18720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18722 = 10'h278 == r_count_24_io_out ? io_r_632_b : _GEN_18721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18723 = 10'h279 == r_count_24_io_out ? io_r_633_b : _GEN_18722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18724 = 10'h27a == r_count_24_io_out ? io_r_634_b : _GEN_18723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18725 = 10'h27b == r_count_24_io_out ? io_r_635_b : _GEN_18724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18726 = 10'h27c == r_count_24_io_out ? io_r_636_b : _GEN_18725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18727 = 10'h27d == r_count_24_io_out ? io_r_637_b : _GEN_18726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18728 = 10'h27e == r_count_24_io_out ? io_r_638_b : _GEN_18727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18729 = 10'h27f == r_count_24_io_out ? io_r_639_b : _GEN_18728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18730 = 10'h280 == r_count_24_io_out ? io_r_640_b : _GEN_18729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18731 = 10'h281 == r_count_24_io_out ? io_r_641_b : _GEN_18730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18732 = 10'h282 == r_count_24_io_out ? io_r_642_b : _GEN_18731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18733 = 10'h283 == r_count_24_io_out ? io_r_643_b : _GEN_18732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18734 = 10'h284 == r_count_24_io_out ? io_r_644_b : _GEN_18733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18735 = 10'h285 == r_count_24_io_out ? io_r_645_b : _GEN_18734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18736 = 10'h286 == r_count_24_io_out ? io_r_646_b : _GEN_18735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18737 = 10'h287 == r_count_24_io_out ? io_r_647_b : _GEN_18736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18738 = 10'h288 == r_count_24_io_out ? io_r_648_b : _GEN_18737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18739 = 10'h289 == r_count_24_io_out ? io_r_649_b : _GEN_18738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18740 = 10'h28a == r_count_24_io_out ? io_r_650_b : _GEN_18739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18741 = 10'h28b == r_count_24_io_out ? io_r_651_b : _GEN_18740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18742 = 10'h28c == r_count_24_io_out ? io_r_652_b : _GEN_18741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18743 = 10'h28d == r_count_24_io_out ? io_r_653_b : _GEN_18742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18744 = 10'h28e == r_count_24_io_out ? io_r_654_b : _GEN_18743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18745 = 10'h28f == r_count_24_io_out ? io_r_655_b : _GEN_18744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18746 = 10'h290 == r_count_24_io_out ? io_r_656_b : _GEN_18745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18747 = 10'h291 == r_count_24_io_out ? io_r_657_b : _GEN_18746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18748 = 10'h292 == r_count_24_io_out ? io_r_658_b : _GEN_18747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18749 = 10'h293 == r_count_24_io_out ? io_r_659_b : _GEN_18748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18750 = 10'h294 == r_count_24_io_out ? io_r_660_b : _GEN_18749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18751 = 10'h295 == r_count_24_io_out ? io_r_661_b : _GEN_18750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18752 = 10'h296 == r_count_24_io_out ? io_r_662_b : _GEN_18751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18753 = 10'h297 == r_count_24_io_out ? io_r_663_b : _GEN_18752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18754 = 10'h298 == r_count_24_io_out ? io_r_664_b : _GEN_18753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18755 = 10'h299 == r_count_24_io_out ? io_r_665_b : _GEN_18754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18756 = 10'h29a == r_count_24_io_out ? io_r_666_b : _GEN_18755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18757 = 10'h29b == r_count_24_io_out ? io_r_667_b : _GEN_18756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18758 = 10'h29c == r_count_24_io_out ? io_r_668_b : _GEN_18757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18759 = 10'h29d == r_count_24_io_out ? io_r_669_b : _GEN_18758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18760 = 10'h29e == r_count_24_io_out ? io_r_670_b : _GEN_18759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18761 = 10'h29f == r_count_24_io_out ? io_r_671_b : _GEN_18760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18762 = 10'h2a0 == r_count_24_io_out ? io_r_672_b : _GEN_18761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18763 = 10'h2a1 == r_count_24_io_out ? io_r_673_b : _GEN_18762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18764 = 10'h2a2 == r_count_24_io_out ? io_r_674_b : _GEN_18763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18765 = 10'h2a3 == r_count_24_io_out ? io_r_675_b : _GEN_18764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18766 = 10'h2a4 == r_count_24_io_out ? io_r_676_b : _GEN_18765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18767 = 10'h2a5 == r_count_24_io_out ? io_r_677_b : _GEN_18766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18768 = 10'h2a6 == r_count_24_io_out ? io_r_678_b : _GEN_18767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18769 = 10'h2a7 == r_count_24_io_out ? io_r_679_b : _GEN_18768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18770 = 10'h2a8 == r_count_24_io_out ? io_r_680_b : _GEN_18769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18771 = 10'h2a9 == r_count_24_io_out ? io_r_681_b : _GEN_18770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18772 = 10'h2aa == r_count_24_io_out ? io_r_682_b : _GEN_18771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18773 = 10'h2ab == r_count_24_io_out ? io_r_683_b : _GEN_18772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18774 = 10'h2ac == r_count_24_io_out ? io_r_684_b : _GEN_18773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18775 = 10'h2ad == r_count_24_io_out ? io_r_685_b : _GEN_18774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18776 = 10'h2ae == r_count_24_io_out ? io_r_686_b : _GEN_18775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18777 = 10'h2af == r_count_24_io_out ? io_r_687_b : _GEN_18776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18778 = 10'h2b0 == r_count_24_io_out ? io_r_688_b : _GEN_18777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18779 = 10'h2b1 == r_count_24_io_out ? io_r_689_b : _GEN_18778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18780 = 10'h2b2 == r_count_24_io_out ? io_r_690_b : _GEN_18779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18781 = 10'h2b3 == r_count_24_io_out ? io_r_691_b : _GEN_18780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18782 = 10'h2b4 == r_count_24_io_out ? io_r_692_b : _GEN_18781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18783 = 10'h2b5 == r_count_24_io_out ? io_r_693_b : _GEN_18782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18784 = 10'h2b6 == r_count_24_io_out ? io_r_694_b : _GEN_18783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18785 = 10'h2b7 == r_count_24_io_out ? io_r_695_b : _GEN_18784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18786 = 10'h2b8 == r_count_24_io_out ? io_r_696_b : _GEN_18785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18787 = 10'h2b9 == r_count_24_io_out ? io_r_697_b : _GEN_18786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18788 = 10'h2ba == r_count_24_io_out ? io_r_698_b : _GEN_18787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18789 = 10'h2bb == r_count_24_io_out ? io_r_699_b : _GEN_18788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18790 = 10'h2bc == r_count_24_io_out ? io_r_700_b : _GEN_18789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18791 = 10'h2bd == r_count_24_io_out ? io_r_701_b : _GEN_18790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18792 = 10'h2be == r_count_24_io_out ? io_r_702_b : _GEN_18791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18793 = 10'h2bf == r_count_24_io_out ? io_r_703_b : _GEN_18792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18794 = 10'h2c0 == r_count_24_io_out ? io_r_704_b : _GEN_18793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18795 = 10'h2c1 == r_count_24_io_out ? io_r_705_b : _GEN_18794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18796 = 10'h2c2 == r_count_24_io_out ? io_r_706_b : _GEN_18795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18797 = 10'h2c3 == r_count_24_io_out ? io_r_707_b : _GEN_18796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18798 = 10'h2c4 == r_count_24_io_out ? io_r_708_b : _GEN_18797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18799 = 10'h2c5 == r_count_24_io_out ? io_r_709_b : _GEN_18798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18800 = 10'h2c6 == r_count_24_io_out ? io_r_710_b : _GEN_18799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18801 = 10'h2c7 == r_count_24_io_out ? io_r_711_b : _GEN_18800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18802 = 10'h2c8 == r_count_24_io_out ? io_r_712_b : _GEN_18801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18803 = 10'h2c9 == r_count_24_io_out ? io_r_713_b : _GEN_18802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18804 = 10'h2ca == r_count_24_io_out ? io_r_714_b : _GEN_18803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18805 = 10'h2cb == r_count_24_io_out ? io_r_715_b : _GEN_18804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18806 = 10'h2cc == r_count_24_io_out ? io_r_716_b : _GEN_18805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18807 = 10'h2cd == r_count_24_io_out ? io_r_717_b : _GEN_18806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18808 = 10'h2ce == r_count_24_io_out ? io_r_718_b : _GEN_18807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18809 = 10'h2cf == r_count_24_io_out ? io_r_719_b : _GEN_18808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18810 = 10'h2d0 == r_count_24_io_out ? io_r_720_b : _GEN_18809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18811 = 10'h2d1 == r_count_24_io_out ? io_r_721_b : _GEN_18810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18812 = 10'h2d2 == r_count_24_io_out ? io_r_722_b : _GEN_18811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18813 = 10'h2d3 == r_count_24_io_out ? io_r_723_b : _GEN_18812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18814 = 10'h2d4 == r_count_24_io_out ? io_r_724_b : _GEN_18813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18815 = 10'h2d5 == r_count_24_io_out ? io_r_725_b : _GEN_18814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18816 = 10'h2d6 == r_count_24_io_out ? io_r_726_b : _GEN_18815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18817 = 10'h2d7 == r_count_24_io_out ? io_r_727_b : _GEN_18816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18818 = 10'h2d8 == r_count_24_io_out ? io_r_728_b : _GEN_18817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18819 = 10'h2d9 == r_count_24_io_out ? io_r_729_b : _GEN_18818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18820 = 10'h2da == r_count_24_io_out ? io_r_730_b : _GEN_18819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18821 = 10'h2db == r_count_24_io_out ? io_r_731_b : _GEN_18820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18822 = 10'h2dc == r_count_24_io_out ? io_r_732_b : _GEN_18821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18823 = 10'h2dd == r_count_24_io_out ? io_r_733_b : _GEN_18822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18824 = 10'h2de == r_count_24_io_out ? io_r_734_b : _GEN_18823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18825 = 10'h2df == r_count_24_io_out ? io_r_735_b : _GEN_18824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18826 = 10'h2e0 == r_count_24_io_out ? io_r_736_b : _GEN_18825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18827 = 10'h2e1 == r_count_24_io_out ? io_r_737_b : _GEN_18826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18828 = 10'h2e2 == r_count_24_io_out ? io_r_738_b : _GEN_18827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18829 = 10'h2e3 == r_count_24_io_out ? io_r_739_b : _GEN_18828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18830 = 10'h2e4 == r_count_24_io_out ? io_r_740_b : _GEN_18829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18831 = 10'h2e5 == r_count_24_io_out ? io_r_741_b : _GEN_18830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18832 = 10'h2e6 == r_count_24_io_out ? io_r_742_b : _GEN_18831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18833 = 10'h2e7 == r_count_24_io_out ? io_r_743_b : _GEN_18832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18834 = 10'h2e8 == r_count_24_io_out ? io_r_744_b : _GEN_18833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18835 = 10'h2e9 == r_count_24_io_out ? io_r_745_b : _GEN_18834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18836 = 10'h2ea == r_count_24_io_out ? io_r_746_b : _GEN_18835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18837 = 10'h2eb == r_count_24_io_out ? io_r_747_b : _GEN_18836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18838 = 10'h2ec == r_count_24_io_out ? io_r_748_b : _GEN_18837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18841 = 10'h1 == r_count_25_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18842 = 10'h2 == r_count_25_io_out ? io_r_2_b : _GEN_18841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18843 = 10'h3 == r_count_25_io_out ? io_r_3_b : _GEN_18842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18844 = 10'h4 == r_count_25_io_out ? io_r_4_b : _GEN_18843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18845 = 10'h5 == r_count_25_io_out ? io_r_5_b : _GEN_18844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18846 = 10'h6 == r_count_25_io_out ? io_r_6_b : _GEN_18845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18847 = 10'h7 == r_count_25_io_out ? io_r_7_b : _GEN_18846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18848 = 10'h8 == r_count_25_io_out ? io_r_8_b : _GEN_18847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18849 = 10'h9 == r_count_25_io_out ? io_r_9_b : _GEN_18848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18850 = 10'ha == r_count_25_io_out ? io_r_10_b : _GEN_18849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18851 = 10'hb == r_count_25_io_out ? io_r_11_b : _GEN_18850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18852 = 10'hc == r_count_25_io_out ? io_r_12_b : _GEN_18851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18853 = 10'hd == r_count_25_io_out ? io_r_13_b : _GEN_18852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18854 = 10'he == r_count_25_io_out ? io_r_14_b : _GEN_18853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18855 = 10'hf == r_count_25_io_out ? io_r_15_b : _GEN_18854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18856 = 10'h10 == r_count_25_io_out ? io_r_16_b : _GEN_18855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18857 = 10'h11 == r_count_25_io_out ? io_r_17_b : _GEN_18856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18858 = 10'h12 == r_count_25_io_out ? io_r_18_b : _GEN_18857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18859 = 10'h13 == r_count_25_io_out ? io_r_19_b : _GEN_18858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18860 = 10'h14 == r_count_25_io_out ? io_r_20_b : _GEN_18859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18861 = 10'h15 == r_count_25_io_out ? io_r_21_b : _GEN_18860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18862 = 10'h16 == r_count_25_io_out ? io_r_22_b : _GEN_18861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18863 = 10'h17 == r_count_25_io_out ? io_r_23_b : _GEN_18862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18864 = 10'h18 == r_count_25_io_out ? io_r_24_b : _GEN_18863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18865 = 10'h19 == r_count_25_io_out ? io_r_25_b : _GEN_18864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18866 = 10'h1a == r_count_25_io_out ? io_r_26_b : _GEN_18865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18867 = 10'h1b == r_count_25_io_out ? io_r_27_b : _GEN_18866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18868 = 10'h1c == r_count_25_io_out ? io_r_28_b : _GEN_18867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18869 = 10'h1d == r_count_25_io_out ? io_r_29_b : _GEN_18868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18870 = 10'h1e == r_count_25_io_out ? io_r_30_b : _GEN_18869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18871 = 10'h1f == r_count_25_io_out ? io_r_31_b : _GEN_18870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18872 = 10'h20 == r_count_25_io_out ? io_r_32_b : _GEN_18871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18873 = 10'h21 == r_count_25_io_out ? io_r_33_b : _GEN_18872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18874 = 10'h22 == r_count_25_io_out ? io_r_34_b : _GEN_18873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18875 = 10'h23 == r_count_25_io_out ? io_r_35_b : _GEN_18874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18876 = 10'h24 == r_count_25_io_out ? io_r_36_b : _GEN_18875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18877 = 10'h25 == r_count_25_io_out ? io_r_37_b : _GEN_18876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18878 = 10'h26 == r_count_25_io_out ? io_r_38_b : _GEN_18877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18879 = 10'h27 == r_count_25_io_out ? io_r_39_b : _GEN_18878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18880 = 10'h28 == r_count_25_io_out ? io_r_40_b : _GEN_18879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18881 = 10'h29 == r_count_25_io_out ? io_r_41_b : _GEN_18880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18882 = 10'h2a == r_count_25_io_out ? io_r_42_b : _GEN_18881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18883 = 10'h2b == r_count_25_io_out ? io_r_43_b : _GEN_18882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18884 = 10'h2c == r_count_25_io_out ? io_r_44_b : _GEN_18883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18885 = 10'h2d == r_count_25_io_out ? io_r_45_b : _GEN_18884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18886 = 10'h2e == r_count_25_io_out ? io_r_46_b : _GEN_18885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18887 = 10'h2f == r_count_25_io_out ? io_r_47_b : _GEN_18886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18888 = 10'h30 == r_count_25_io_out ? io_r_48_b : _GEN_18887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18889 = 10'h31 == r_count_25_io_out ? io_r_49_b : _GEN_18888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18890 = 10'h32 == r_count_25_io_out ? io_r_50_b : _GEN_18889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18891 = 10'h33 == r_count_25_io_out ? io_r_51_b : _GEN_18890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18892 = 10'h34 == r_count_25_io_out ? io_r_52_b : _GEN_18891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18893 = 10'h35 == r_count_25_io_out ? io_r_53_b : _GEN_18892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18894 = 10'h36 == r_count_25_io_out ? io_r_54_b : _GEN_18893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18895 = 10'h37 == r_count_25_io_out ? io_r_55_b : _GEN_18894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18896 = 10'h38 == r_count_25_io_out ? io_r_56_b : _GEN_18895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18897 = 10'h39 == r_count_25_io_out ? io_r_57_b : _GEN_18896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18898 = 10'h3a == r_count_25_io_out ? io_r_58_b : _GEN_18897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18899 = 10'h3b == r_count_25_io_out ? io_r_59_b : _GEN_18898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18900 = 10'h3c == r_count_25_io_out ? io_r_60_b : _GEN_18899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18901 = 10'h3d == r_count_25_io_out ? io_r_61_b : _GEN_18900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18902 = 10'h3e == r_count_25_io_out ? io_r_62_b : _GEN_18901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18903 = 10'h3f == r_count_25_io_out ? io_r_63_b : _GEN_18902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18904 = 10'h40 == r_count_25_io_out ? io_r_64_b : _GEN_18903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18905 = 10'h41 == r_count_25_io_out ? io_r_65_b : _GEN_18904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18906 = 10'h42 == r_count_25_io_out ? io_r_66_b : _GEN_18905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18907 = 10'h43 == r_count_25_io_out ? io_r_67_b : _GEN_18906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18908 = 10'h44 == r_count_25_io_out ? io_r_68_b : _GEN_18907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18909 = 10'h45 == r_count_25_io_out ? io_r_69_b : _GEN_18908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18910 = 10'h46 == r_count_25_io_out ? io_r_70_b : _GEN_18909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18911 = 10'h47 == r_count_25_io_out ? io_r_71_b : _GEN_18910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18912 = 10'h48 == r_count_25_io_out ? io_r_72_b : _GEN_18911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18913 = 10'h49 == r_count_25_io_out ? io_r_73_b : _GEN_18912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18914 = 10'h4a == r_count_25_io_out ? io_r_74_b : _GEN_18913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18915 = 10'h4b == r_count_25_io_out ? io_r_75_b : _GEN_18914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18916 = 10'h4c == r_count_25_io_out ? io_r_76_b : _GEN_18915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18917 = 10'h4d == r_count_25_io_out ? io_r_77_b : _GEN_18916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18918 = 10'h4e == r_count_25_io_out ? io_r_78_b : _GEN_18917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18919 = 10'h4f == r_count_25_io_out ? io_r_79_b : _GEN_18918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18920 = 10'h50 == r_count_25_io_out ? io_r_80_b : _GEN_18919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18921 = 10'h51 == r_count_25_io_out ? io_r_81_b : _GEN_18920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18922 = 10'h52 == r_count_25_io_out ? io_r_82_b : _GEN_18921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18923 = 10'h53 == r_count_25_io_out ? io_r_83_b : _GEN_18922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18924 = 10'h54 == r_count_25_io_out ? io_r_84_b : _GEN_18923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18925 = 10'h55 == r_count_25_io_out ? io_r_85_b : _GEN_18924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18926 = 10'h56 == r_count_25_io_out ? io_r_86_b : _GEN_18925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18927 = 10'h57 == r_count_25_io_out ? io_r_87_b : _GEN_18926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18928 = 10'h58 == r_count_25_io_out ? io_r_88_b : _GEN_18927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18929 = 10'h59 == r_count_25_io_out ? io_r_89_b : _GEN_18928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18930 = 10'h5a == r_count_25_io_out ? io_r_90_b : _GEN_18929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18931 = 10'h5b == r_count_25_io_out ? io_r_91_b : _GEN_18930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18932 = 10'h5c == r_count_25_io_out ? io_r_92_b : _GEN_18931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18933 = 10'h5d == r_count_25_io_out ? io_r_93_b : _GEN_18932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18934 = 10'h5e == r_count_25_io_out ? io_r_94_b : _GEN_18933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18935 = 10'h5f == r_count_25_io_out ? io_r_95_b : _GEN_18934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18936 = 10'h60 == r_count_25_io_out ? io_r_96_b : _GEN_18935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18937 = 10'h61 == r_count_25_io_out ? io_r_97_b : _GEN_18936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18938 = 10'h62 == r_count_25_io_out ? io_r_98_b : _GEN_18937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18939 = 10'h63 == r_count_25_io_out ? io_r_99_b : _GEN_18938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18940 = 10'h64 == r_count_25_io_out ? io_r_100_b : _GEN_18939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18941 = 10'h65 == r_count_25_io_out ? io_r_101_b : _GEN_18940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18942 = 10'h66 == r_count_25_io_out ? io_r_102_b : _GEN_18941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18943 = 10'h67 == r_count_25_io_out ? io_r_103_b : _GEN_18942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18944 = 10'h68 == r_count_25_io_out ? io_r_104_b : _GEN_18943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18945 = 10'h69 == r_count_25_io_out ? io_r_105_b : _GEN_18944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18946 = 10'h6a == r_count_25_io_out ? io_r_106_b : _GEN_18945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18947 = 10'h6b == r_count_25_io_out ? io_r_107_b : _GEN_18946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18948 = 10'h6c == r_count_25_io_out ? io_r_108_b : _GEN_18947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18949 = 10'h6d == r_count_25_io_out ? io_r_109_b : _GEN_18948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18950 = 10'h6e == r_count_25_io_out ? io_r_110_b : _GEN_18949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18951 = 10'h6f == r_count_25_io_out ? io_r_111_b : _GEN_18950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18952 = 10'h70 == r_count_25_io_out ? io_r_112_b : _GEN_18951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18953 = 10'h71 == r_count_25_io_out ? io_r_113_b : _GEN_18952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18954 = 10'h72 == r_count_25_io_out ? io_r_114_b : _GEN_18953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18955 = 10'h73 == r_count_25_io_out ? io_r_115_b : _GEN_18954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18956 = 10'h74 == r_count_25_io_out ? io_r_116_b : _GEN_18955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18957 = 10'h75 == r_count_25_io_out ? io_r_117_b : _GEN_18956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18958 = 10'h76 == r_count_25_io_out ? io_r_118_b : _GEN_18957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18959 = 10'h77 == r_count_25_io_out ? io_r_119_b : _GEN_18958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18960 = 10'h78 == r_count_25_io_out ? io_r_120_b : _GEN_18959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18961 = 10'h79 == r_count_25_io_out ? io_r_121_b : _GEN_18960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18962 = 10'h7a == r_count_25_io_out ? io_r_122_b : _GEN_18961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18963 = 10'h7b == r_count_25_io_out ? io_r_123_b : _GEN_18962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18964 = 10'h7c == r_count_25_io_out ? io_r_124_b : _GEN_18963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18965 = 10'h7d == r_count_25_io_out ? io_r_125_b : _GEN_18964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18966 = 10'h7e == r_count_25_io_out ? io_r_126_b : _GEN_18965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18967 = 10'h7f == r_count_25_io_out ? io_r_127_b : _GEN_18966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18968 = 10'h80 == r_count_25_io_out ? io_r_128_b : _GEN_18967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18969 = 10'h81 == r_count_25_io_out ? io_r_129_b : _GEN_18968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18970 = 10'h82 == r_count_25_io_out ? io_r_130_b : _GEN_18969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18971 = 10'h83 == r_count_25_io_out ? io_r_131_b : _GEN_18970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18972 = 10'h84 == r_count_25_io_out ? io_r_132_b : _GEN_18971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18973 = 10'h85 == r_count_25_io_out ? io_r_133_b : _GEN_18972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18974 = 10'h86 == r_count_25_io_out ? io_r_134_b : _GEN_18973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18975 = 10'h87 == r_count_25_io_out ? io_r_135_b : _GEN_18974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18976 = 10'h88 == r_count_25_io_out ? io_r_136_b : _GEN_18975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18977 = 10'h89 == r_count_25_io_out ? io_r_137_b : _GEN_18976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18978 = 10'h8a == r_count_25_io_out ? io_r_138_b : _GEN_18977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18979 = 10'h8b == r_count_25_io_out ? io_r_139_b : _GEN_18978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18980 = 10'h8c == r_count_25_io_out ? io_r_140_b : _GEN_18979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18981 = 10'h8d == r_count_25_io_out ? io_r_141_b : _GEN_18980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18982 = 10'h8e == r_count_25_io_out ? io_r_142_b : _GEN_18981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18983 = 10'h8f == r_count_25_io_out ? io_r_143_b : _GEN_18982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18984 = 10'h90 == r_count_25_io_out ? io_r_144_b : _GEN_18983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18985 = 10'h91 == r_count_25_io_out ? io_r_145_b : _GEN_18984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18986 = 10'h92 == r_count_25_io_out ? io_r_146_b : _GEN_18985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18987 = 10'h93 == r_count_25_io_out ? io_r_147_b : _GEN_18986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18988 = 10'h94 == r_count_25_io_out ? io_r_148_b : _GEN_18987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18989 = 10'h95 == r_count_25_io_out ? io_r_149_b : _GEN_18988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18990 = 10'h96 == r_count_25_io_out ? io_r_150_b : _GEN_18989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18991 = 10'h97 == r_count_25_io_out ? io_r_151_b : _GEN_18990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18992 = 10'h98 == r_count_25_io_out ? io_r_152_b : _GEN_18991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18993 = 10'h99 == r_count_25_io_out ? io_r_153_b : _GEN_18992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18994 = 10'h9a == r_count_25_io_out ? io_r_154_b : _GEN_18993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18995 = 10'h9b == r_count_25_io_out ? io_r_155_b : _GEN_18994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18996 = 10'h9c == r_count_25_io_out ? io_r_156_b : _GEN_18995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18997 = 10'h9d == r_count_25_io_out ? io_r_157_b : _GEN_18996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18998 = 10'h9e == r_count_25_io_out ? io_r_158_b : _GEN_18997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18999 = 10'h9f == r_count_25_io_out ? io_r_159_b : _GEN_18998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19000 = 10'ha0 == r_count_25_io_out ? io_r_160_b : _GEN_18999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19001 = 10'ha1 == r_count_25_io_out ? io_r_161_b : _GEN_19000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19002 = 10'ha2 == r_count_25_io_out ? io_r_162_b : _GEN_19001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19003 = 10'ha3 == r_count_25_io_out ? io_r_163_b : _GEN_19002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19004 = 10'ha4 == r_count_25_io_out ? io_r_164_b : _GEN_19003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19005 = 10'ha5 == r_count_25_io_out ? io_r_165_b : _GEN_19004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19006 = 10'ha6 == r_count_25_io_out ? io_r_166_b : _GEN_19005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19007 = 10'ha7 == r_count_25_io_out ? io_r_167_b : _GEN_19006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19008 = 10'ha8 == r_count_25_io_out ? io_r_168_b : _GEN_19007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19009 = 10'ha9 == r_count_25_io_out ? io_r_169_b : _GEN_19008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19010 = 10'haa == r_count_25_io_out ? io_r_170_b : _GEN_19009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19011 = 10'hab == r_count_25_io_out ? io_r_171_b : _GEN_19010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19012 = 10'hac == r_count_25_io_out ? io_r_172_b : _GEN_19011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19013 = 10'had == r_count_25_io_out ? io_r_173_b : _GEN_19012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19014 = 10'hae == r_count_25_io_out ? io_r_174_b : _GEN_19013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19015 = 10'haf == r_count_25_io_out ? io_r_175_b : _GEN_19014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19016 = 10'hb0 == r_count_25_io_out ? io_r_176_b : _GEN_19015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19017 = 10'hb1 == r_count_25_io_out ? io_r_177_b : _GEN_19016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19018 = 10'hb2 == r_count_25_io_out ? io_r_178_b : _GEN_19017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19019 = 10'hb3 == r_count_25_io_out ? io_r_179_b : _GEN_19018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19020 = 10'hb4 == r_count_25_io_out ? io_r_180_b : _GEN_19019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19021 = 10'hb5 == r_count_25_io_out ? io_r_181_b : _GEN_19020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19022 = 10'hb6 == r_count_25_io_out ? io_r_182_b : _GEN_19021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19023 = 10'hb7 == r_count_25_io_out ? io_r_183_b : _GEN_19022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19024 = 10'hb8 == r_count_25_io_out ? io_r_184_b : _GEN_19023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19025 = 10'hb9 == r_count_25_io_out ? io_r_185_b : _GEN_19024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19026 = 10'hba == r_count_25_io_out ? io_r_186_b : _GEN_19025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19027 = 10'hbb == r_count_25_io_out ? io_r_187_b : _GEN_19026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19028 = 10'hbc == r_count_25_io_out ? io_r_188_b : _GEN_19027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19029 = 10'hbd == r_count_25_io_out ? io_r_189_b : _GEN_19028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19030 = 10'hbe == r_count_25_io_out ? io_r_190_b : _GEN_19029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19031 = 10'hbf == r_count_25_io_out ? io_r_191_b : _GEN_19030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19032 = 10'hc0 == r_count_25_io_out ? io_r_192_b : _GEN_19031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19033 = 10'hc1 == r_count_25_io_out ? io_r_193_b : _GEN_19032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19034 = 10'hc2 == r_count_25_io_out ? io_r_194_b : _GEN_19033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19035 = 10'hc3 == r_count_25_io_out ? io_r_195_b : _GEN_19034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19036 = 10'hc4 == r_count_25_io_out ? io_r_196_b : _GEN_19035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19037 = 10'hc5 == r_count_25_io_out ? io_r_197_b : _GEN_19036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19038 = 10'hc6 == r_count_25_io_out ? io_r_198_b : _GEN_19037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19039 = 10'hc7 == r_count_25_io_out ? io_r_199_b : _GEN_19038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19040 = 10'hc8 == r_count_25_io_out ? io_r_200_b : _GEN_19039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19041 = 10'hc9 == r_count_25_io_out ? io_r_201_b : _GEN_19040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19042 = 10'hca == r_count_25_io_out ? io_r_202_b : _GEN_19041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19043 = 10'hcb == r_count_25_io_out ? io_r_203_b : _GEN_19042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19044 = 10'hcc == r_count_25_io_out ? io_r_204_b : _GEN_19043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19045 = 10'hcd == r_count_25_io_out ? io_r_205_b : _GEN_19044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19046 = 10'hce == r_count_25_io_out ? io_r_206_b : _GEN_19045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19047 = 10'hcf == r_count_25_io_out ? io_r_207_b : _GEN_19046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19048 = 10'hd0 == r_count_25_io_out ? io_r_208_b : _GEN_19047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19049 = 10'hd1 == r_count_25_io_out ? io_r_209_b : _GEN_19048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19050 = 10'hd2 == r_count_25_io_out ? io_r_210_b : _GEN_19049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19051 = 10'hd3 == r_count_25_io_out ? io_r_211_b : _GEN_19050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19052 = 10'hd4 == r_count_25_io_out ? io_r_212_b : _GEN_19051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19053 = 10'hd5 == r_count_25_io_out ? io_r_213_b : _GEN_19052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19054 = 10'hd6 == r_count_25_io_out ? io_r_214_b : _GEN_19053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19055 = 10'hd7 == r_count_25_io_out ? io_r_215_b : _GEN_19054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19056 = 10'hd8 == r_count_25_io_out ? io_r_216_b : _GEN_19055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19057 = 10'hd9 == r_count_25_io_out ? io_r_217_b : _GEN_19056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19058 = 10'hda == r_count_25_io_out ? io_r_218_b : _GEN_19057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19059 = 10'hdb == r_count_25_io_out ? io_r_219_b : _GEN_19058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19060 = 10'hdc == r_count_25_io_out ? io_r_220_b : _GEN_19059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19061 = 10'hdd == r_count_25_io_out ? io_r_221_b : _GEN_19060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19062 = 10'hde == r_count_25_io_out ? io_r_222_b : _GEN_19061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19063 = 10'hdf == r_count_25_io_out ? io_r_223_b : _GEN_19062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19064 = 10'he0 == r_count_25_io_out ? io_r_224_b : _GEN_19063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19065 = 10'he1 == r_count_25_io_out ? io_r_225_b : _GEN_19064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19066 = 10'he2 == r_count_25_io_out ? io_r_226_b : _GEN_19065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19067 = 10'he3 == r_count_25_io_out ? io_r_227_b : _GEN_19066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19068 = 10'he4 == r_count_25_io_out ? io_r_228_b : _GEN_19067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19069 = 10'he5 == r_count_25_io_out ? io_r_229_b : _GEN_19068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19070 = 10'he6 == r_count_25_io_out ? io_r_230_b : _GEN_19069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19071 = 10'he7 == r_count_25_io_out ? io_r_231_b : _GEN_19070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19072 = 10'he8 == r_count_25_io_out ? io_r_232_b : _GEN_19071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19073 = 10'he9 == r_count_25_io_out ? io_r_233_b : _GEN_19072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19074 = 10'hea == r_count_25_io_out ? io_r_234_b : _GEN_19073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19075 = 10'heb == r_count_25_io_out ? io_r_235_b : _GEN_19074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19076 = 10'hec == r_count_25_io_out ? io_r_236_b : _GEN_19075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19077 = 10'hed == r_count_25_io_out ? io_r_237_b : _GEN_19076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19078 = 10'hee == r_count_25_io_out ? io_r_238_b : _GEN_19077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19079 = 10'hef == r_count_25_io_out ? io_r_239_b : _GEN_19078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19080 = 10'hf0 == r_count_25_io_out ? io_r_240_b : _GEN_19079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19081 = 10'hf1 == r_count_25_io_out ? io_r_241_b : _GEN_19080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19082 = 10'hf2 == r_count_25_io_out ? io_r_242_b : _GEN_19081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19083 = 10'hf3 == r_count_25_io_out ? io_r_243_b : _GEN_19082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19084 = 10'hf4 == r_count_25_io_out ? io_r_244_b : _GEN_19083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19085 = 10'hf5 == r_count_25_io_out ? io_r_245_b : _GEN_19084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19086 = 10'hf6 == r_count_25_io_out ? io_r_246_b : _GEN_19085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19087 = 10'hf7 == r_count_25_io_out ? io_r_247_b : _GEN_19086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19088 = 10'hf8 == r_count_25_io_out ? io_r_248_b : _GEN_19087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19089 = 10'hf9 == r_count_25_io_out ? io_r_249_b : _GEN_19088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19090 = 10'hfa == r_count_25_io_out ? io_r_250_b : _GEN_19089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19091 = 10'hfb == r_count_25_io_out ? io_r_251_b : _GEN_19090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19092 = 10'hfc == r_count_25_io_out ? io_r_252_b : _GEN_19091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19093 = 10'hfd == r_count_25_io_out ? io_r_253_b : _GEN_19092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19094 = 10'hfe == r_count_25_io_out ? io_r_254_b : _GEN_19093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19095 = 10'hff == r_count_25_io_out ? io_r_255_b : _GEN_19094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19096 = 10'h100 == r_count_25_io_out ? io_r_256_b : _GEN_19095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19097 = 10'h101 == r_count_25_io_out ? io_r_257_b : _GEN_19096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19098 = 10'h102 == r_count_25_io_out ? io_r_258_b : _GEN_19097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19099 = 10'h103 == r_count_25_io_out ? io_r_259_b : _GEN_19098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19100 = 10'h104 == r_count_25_io_out ? io_r_260_b : _GEN_19099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19101 = 10'h105 == r_count_25_io_out ? io_r_261_b : _GEN_19100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19102 = 10'h106 == r_count_25_io_out ? io_r_262_b : _GEN_19101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19103 = 10'h107 == r_count_25_io_out ? io_r_263_b : _GEN_19102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19104 = 10'h108 == r_count_25_io_out ? io_r_264_b : _GEN_19103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19105 = 10'h109 == r_count_25_io_out ? io_r_265_b : _GEN_19104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19106 = 10'h10a == r_count_25_io_out ? io_r_266_b : _GEN_19105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19107 = 10'h10b == r_count_25_io_out ? io_r_267_b : _GEN_19106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19108 = 10'h10c == r_count_25_io_out ? io_r_268_b : _GEN_19107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19109 = 10'h10d == r_count_25_io_out ? io_r_269_b : _GEN_19108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19110 = 10'h10e == r_count_25_io_out ? io_r_270_b : _GEN_19109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19111 = 10'h10f == r_count_25_io_out ? io_r_271_b : _GEN_19110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19112 = 10'h110 == r_count_25_io_out ? io_r_272_b : _GEN_19111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19113 = 10'h111 == r_count_25_io_out ? io_r_273_b : _GEN_19112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19114 = 10'h112 == r_count_25_io_out ? io_r_274_b : _GEN_19113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19115 = 10'h113 == r_count_25_io_out ? io_r_275_b : _GEN_19114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19116 = 10'h114 == r_count_25_io_out ? io_r_276_b : _GEN_19115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19117 = 10'h115 == r_count_25_io_out ? io_r_277_b : _GEN_19116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19118 = 10'h116 == r_count_25_io_out ? io_r_278_b : _GEN_19117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19119 = 10'h117 == r_count_25_io_out ? io_r_279_b : _GEN_19118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19120 = 10'h118 == r_count_25_io_out ? io_r_280_b : _GEN_19119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19121 = 10'h119 == r_count_25_io_out ? io_r_281_b : _GEN_19120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19122 = 10'h11a == r_count_25_io_out ? io_r_282_b : _GEN_19121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19123 = 10'h11b == r_count_25_io_out ? io_r_283_b : _GEN_19122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19124 = 10'h11c == r_count_25_io_out ? io_r_284_b : _GEN_19123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19125 = 10'h11d == r_count_25_io_out ? io_r_285_b : _GEN_19124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19126 = 10'h11e == r_count_25_io_out ? io_r_286_b : _GEN_19125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19127 = 10'h11f == r_count_25_io_out ? io_r_287_b : _GEN_19126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19128 = 10'h120 == r_count_25_io_out ? io_r_288_b : _GEN_19127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19129 = 10'h121 == r_count_25_io_out ? io_r_289_b : _GEN_19128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19130 = 10'h122 == r_count_25_io_out ? io_r_290_b : _GEN_19129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19131 = 10'h123 == r_count_25_io_out ? io_r_291_b : _GEN_19130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19132 = 10'h124 == r_count_25_io_out ? io_r_292_b : _GEN_19131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19133 = 10'h125 == r_count_25_io_out ? io_r_293_b : _GEN_19132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19134 = 10'h126 == r_count_25_io_out ? io_r_294_b : _GEN_19133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19135 = 10'h127 == r_count_25_io_out ? io_r_295_b : _GEN_19134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19136 = 10'h128 == r_count_25_io_out ? io_r_296_b : _GEN_19135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19137 = 10'h129 == r_count_25_io_out ? io_r_297_b : _GEN_19136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19138 = 10'h12a == r_count_25_io_out ? io_r_298_b : _GEN_19137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19139 = 10'h12b == r_count_25_io_out ? io_r_299_b : _GEN_19138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19140 = 10'h12c == r_count_25_io_out ? io_r_300_b : _GEN_19139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19141 = 10'h12d == r_count_25_io_out ? io_r_301_b : _GEN_19140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19142 = 10'h12e == r_count_25_io_out ? io_r_302_b : _GEN_19141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19143 = 10'h12f == r_count_25_io_out ? io_r_303_b : _GEN_19142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19144 = 10'h130 == r_count_25_io_out ? io_r_304_b : _GEN_19143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19145 = 10'h131 == r_count_25_io_out ? io_r_305_b : _GEN_19144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19146 = 10'h132 == r_count_25_io_out ? io_r_306_b : _GEN_19145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19147 = 10'h133 == r_count_25_io_out ? io_r_307_b : _GEN_19146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19148 = 10'h134 == r_count_25_io_out ? io_r_308_b : _GEN_19147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19149 = 10'h135 == r_count_25_io_out ? io_r_309_b : _GEN_19148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19150 = 10'h136 == r_count_25_io_out ? io_r_310_b : _GEN_19149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19151 = 10'h137 == r_count_25_io_out ? io_r_311_b : _GEN_19150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19152 = 10'h138 == r_count_25_io_out ? io_r_312_b : _GEN_19151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19153 = 10'h139 == r_count_25_io_out ? io_r_313_b : _GEN_19152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19154 = 10'h13a == r_count_25_io_out ? io_r_314_b : _GEN_19153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19155 = 10'h13b == r_count_25_io_out ? io_r_315_b : _GEN_19154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19156 = 10'h13c == r_count_25_io_out ? io_r_316_b : _GEN_19155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19157 = 10'h13d == r_count_25_io_out ? io_r_317_b : _GEN_19156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19158 = 10'h13e == r_count_25_io_out ? io_r_318_b : _GEN_19157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19159 = 10'h13f == r_count_25_io_out ? io_r_319_b : _GEN_19158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19160 = 10'h140 == r_count_25_io_out ? io_r_320_b : _GEN_19159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19161 = 10'h141 == r_count_25_io_out ? io_r_321_b : _GEN_19160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19162 = 10'h142 == r_count_25_io_out ? io_r_322_b : _GEN_19161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19163 = 10'h143 == r_count_25_io_out ? io_r_323_b : _GEN_19162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19164 = 10'h144 == r_count_25_io_out ? io_r_324_b : _GEN_19163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19165 = 10'h145 == r_count_25_io_out ? io_r_325_b : _GEN_19164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19166 = 10'h146 == r_count_25_io_out ? io_r_326_b : _GEN_19165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19167 = 10'h147 == r_count_25_io_out ? io_r_327_b : _GEN_19166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19168 = 10'h148 == r_count_25_io_out ? io_r_328_b : _GEN_19167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19169 = 10'h149 == r_count_25_io_out ? io_r_329_b : _GEN_19168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19170 = 10'h14a == r_count_25_io_out ? io_r_330_b : _GEN_19169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19171 = 10'h14b == r_count_25_io_out ? io_r_331_b : _GEN_19170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19172 = 10'h14c == r_count_25_io_out ? io_r_332_b : _GEN_19171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19173 = 10'h14d == r_count_25_io_out ? io_r_333_b : _GEN_19172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19174 = 10'h14e == r_count_25_io_out ? io_r_334_b : _GEN_19173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19175 = 10'h14f == r_count_25_io_out ? io_r_335_b : _GEN_19174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19176 = 10'h150 == r_count_25_io_out ? io_r_336_b : _GEN_19175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19177 = 10'h151 == r_count_25_io_out ? io_r_337_b : _GEN_19176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19178 = 10'h152 == r_count_25_io_out ? io_r_338_b : _GEN_19177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19179 = 10'h153 == r_count_25_io_out ? io_r_339_b : _GEN_19178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19180 = 10'h154 == r_count_25_io_out ? io_r_340_b : _GEN_19179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19181 = 10'h155 == r_count_25_io_out ? io_r_341_b : _GEN_19180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19182 = 10'h156 == r_count_25_io_out ? io_r_342_b : _GEN_19181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19183 = 10'h157 == r_count_25_io_out ? io_r_343_b : _GEN_19182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19184 = 10'h158 == r_count_25_io_out ? io_r_344_b : _GEN_19183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19185 = 10'h159 == r_count_25_io_out ? io_r_345_b : _GEN_19184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19186 = 10'h15a == r_count_25_io_out ? io_r_346_b : _GEN_19185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19187 = 10'h15b == r_count_25_io_out ? io_r_347_b : _GEN_19186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19188 = 10'h15c == r_count_25_io_out ? io_r_348_b : _GEN_19187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19189 = 10'h15d == r_count_25_io_out ? io_r_349_b : _GEN_19188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19190 = 10'h15e == r_count_25_io_out ? io_r_350_b : _GEN_19189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19191 = 10'h15f == r_count_25_io_out ? io_r_351_b : _GEN_19190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19192 = 10'h160 == r_count_25_io_out ? io_r_352_b : _GEN_19191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19193 = 10'h161 == r_count_25_io_out ? io_r_353_b : _GEN_19192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19194 = 10'h162 == r_count_25_io_out ? io_r_354_b : _GEN_19193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19195 = 10'h163 == r_count_25_io_out ? io_r_355_b : _GEN_19194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19196 = 10'h164 == r_count_25_io_out ? io_r_356_b : _GEN_19195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19197 = 10'h165 == r_count_25_io_out ? io_r_357_b : _GEN_19196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19198 = 10'h166 == r_count_25_io_out ? io_r_358_b : _GEN_19197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19199 = 10'h167 == r_count_25_io_out ? io_r_359_b : _GEN_19198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19200 = 10'h168 == r_count_25_io_out ? io_r_360_b : _GEN_19199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19201 = 10'h169 == r_count_25_io_out ? io_r_361_b : _GEN_19200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19202 = 10'h16a == r_count_25_io_out ? io_r_362_b : _GEN_19201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19203 = 10'h16b == r_count_25_io_out ? io_r_363_b : _GEN_19202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19204 = 10'h16c == r_count_25_io_out ? io_r_364_b : _GEN_19203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19205 = 10'h16d == r_count_25_io_out ? io_r_365_b : _GEN_19204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19206 = 10'h16e == r_count_25_io_out ? io_r_366_b : _GEN_19205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19207 = 10'h16f == r_count_25_io_out ? io_r_367_b : _GEN_19206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19208 = 10'h170 == r_count_25_io_out ? io_r_368_b : _GEN_19207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19209 = 10'h171 == r_count_25_io_out ? io_r_369_b : _GEN_19208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19210 = 10'h172 == r_count_25_io_out ? io_r_370_b : _GEN_19209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19211 = 10'h173 == r_count_25_io_out ? io_r_371_b : _GEN_19210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19212 = 10'h174 == r_count_25_io_out ? io_r_372_b : _GEN_19211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19213 = 10'h175 == r_count_25_io_out ? io_r_373_b : _GEN_19212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19214 = 10'h176 == r_count_25_io_out ? io_r_374_b : _GEN_19213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19215 = 10'h177 == r_count_25_io_out ? io_r_375_b : _GEN_19214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19216 = 10'h178 == r_count_25_io_out ? io_r_376_b : _GEN_19215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19217 = 10'h179 == r_count_25_io_out ? io_r_377_b : _GEN_19216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19218 = 10'h17a == r_count_25_io_out ? io_r_378_b : _GEN_19217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19219 = 10'h17b == r_count_25_io_out ? io_r_379_b : _GEN_19218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19220 = 10'h17c == r_count_25_io_out ? io_r_380_b : _GEN_19219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19221 = 10'h17d == r_count_25_io_out ? io_r_381_b : _GEN_19220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19222 = 10'h17e == r_count_25_io_out ? io_r_382_b : _GEN_19221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19223 = 10'h17f == r_count_25_io_out ? io_r_383_b : _GEN_19222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19224 = 10'h180 == r_count_25_io_out ? io_r_384_b : _GEN_19223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19225 = 10'h181 == r_count_25_io_out ? io_r_385_b : _GEN_19224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19226 = 10'h182 == r_count_25_io_out ? io_r_386_b : _GEN_19225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19227 = 10'h183 == r_count_25_io_out ? io_r_387_b : _GEN_19226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19228 = 10'h184 == r_count_25_io_out ? io_r_388_b : _GEN_19227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19229 = 10'h185 == r_count_25_io_out ? io_r_389_b : _GEN_19228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19230 = 10'h186 == r_count_25_io_out ? io_r_390_b : _GEN_19229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19231 = 10'h187 == r_count_25_io_out ? io_r_391_b : _GEN_19230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19232 = 10'h188 == r_count_25_io_out ? io_r_392_b : _GEN_19231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19233 = 10'h189 == r_count_25_io_out ? io_r_393_b : _GEN_19232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19234 = 10'h18a == r_count_25_io_out ? io_r_394_b : _GEN_19233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19235 = 10'h18b == r_count_25_io_out ? io_r_395_b : _GEN_19234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19236 = 10'h18c == r_count_25_io_out ? io_r_396_b : _GEN_19235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19237 = 10'h18d == r_count_25_io_out ? io_r_397_b : _GEN_19236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19238 = 10'h18e == r_count_25_io_out ? io_r_398_b : _GEN_19237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19239 = 10'h18f == r_count_25_io_out ? io_r_399_b : _GEN_19238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19240 = 10'h190 == r_count_25_io_out ? io_r_400_b : _GEN_19239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19241 = 10'h191 == r_count_25_io_out ? io_r_401_b : _GEN_19240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19242 = 10'h192 == r_count_25_io_out ? io_r_402_b : _GEN_19241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19243 = 10'h193 == r_count_25_io_out ? io_r_403_b : _GEN_19242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19244 = 10'h194 == r_count_25_io_out ? io_r_404_b : _GEN_19243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19245 = 10'h195 == r_count_25_io_out ? io_r_405_b : _GEN_19244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19246 = 10'h196 == r_count_25_io_out ? io_r_406_b : _GEN_19245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19247 = 10'h197 == r_count_25_io_out ? io_r_407_b : _GEN_19246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19248 = 10'h198 == r_count_25_io_out ? io_r_408_b : _GEN_19247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19249 = 10'h199 == r_count_25_io_out ? io_r_409_b : _GEN_19248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19250 = 10'h19a == r_count_25_io_out ? io_r_410_b : _GEN_19249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19251 = 10'h19b == r_count_25_io_out ? io_r_411_b : _GEN_19250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19252 = 10'h19c == r_count_25_io_out ? io_r_412_b : _GEN_19251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19253 = 10'h19d == r_count_25_io_out ? io_r_413_b : _GEN_19252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19254 = 10'h19e == r_count_25_io_out ? io_r_414_b : _GEN_19253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19255 = 10'h19f == r_count_25_io_out ? io_r_415_b : _GEN_19254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19256 = 10'h1a0 == r_count_25_io_out ? io_r_416_b : _GEN_19255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19257 = 10'h1a1 == r_count_25_io_out ? io_r_417_b : _GEN_19256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19258 = 10'h1a2 == r_count_25_io_out ? io_r_418_b : _GEN_19257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19259 = 10'h1a3 == r_count_25_io_out ? io_r_419_b : _GEN_19258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19260 = 10'h1a4 == r_count_25_io_out ? io_r_420_b : _GEN_19259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19261 = 10'h1a5 == r_count_25_io_out ? io_r_421_b : _GEN_19260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19262 = 10'h1a6 == r_count_25_io_out ? io_r_422_b : _GEN_19261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19263 = 10'h1a7 == r_count_25_io_out ? io_r_423_b : _GEN_19262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19264 = 10'h1a8 == r_count_25_io_out ? io_r_424_b : _GEN_19263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19265 = 10'h1a9 == r_count_25_io_out ? io_r_425_b : _GEN_19264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19266 = 10'h1aa == r_count_25_io_out ? io_r_426_b : _GEN_19265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19267 = 10'h1ab == r_count_25_io_out ? io_r_427_b : _GEN_19266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19268 = 10'h1ac == r_count_25_io_out ? io_r_428_b : _GEN_19267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19269 = 10'h1ad == r_count_25_io_out ? io_r_429_b : _GEN_19268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19270 = 10'h1ae == r_count_25_io_out ? io_r_430_b : _GEN_19269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19271 = 10'h1af == r_count_25_io_out ? io_r_431_b : _GEN_19270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19272 = 10'h1b0 == r_count_25_io_out ? io_r_432_b : _GEN_19271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19273 = 10'h1b1 == r_count_25_io_out ? io_r_433_b : _GEN_19272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19274 = 10'h1b2 == r_count_25_io_out ? io_r_434_b : _GEN_19273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19275 = 10'h1b3 == r_count_25_io_out ? io_r_435_b : _GEN_19274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19276 = 10'h1b4 == r_count_25_io_out ? io_r_436_b : _GEN_19275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19277 = 10'h1b5 == r_count_25_io_out ? io_r_437_b : _GEN_19276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19278 = 10'h1b6 == r_count_25_io_out ? io_r_438_b : _GEN_19277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19279 = 10'h1b7 == r_count_25_io_out ? io_r_439_b : _GEN_19278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19280 = 10'h1b8 == r_count_25_io_out ? io_r_440_b : _GEN_19279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19281 = 10'h1b9 == r_count_25_io_out ? io_r_441_b : _GEN_19280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19282 = 10'h1ba == r_count_25_io_out ? io_r_442_b : _GEN_19281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19283 = 10'h1bb == r_count_25_io_out ? io_r_443_b : _GEN_19282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19284 = 10'h1bc == r_count_25_io_out ? io_r_444_b : _GEN_19283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19285 = 10'h1bd == r_count_25_io_out ? io_r_445_b : _GEN_19284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19286 = 10'h1be == r_count_25_io_out ? io_r_446_b : _GEN_19285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19287 = 10'h1bf == r_count_25_io_out ? io_r_447_b : _GEN_19286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19288 = 10'h1c0 == r_count_25_io_out ? io_r_448_b : _GEN_19287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19289 = 10'h1c1 == r_count_25_io_out ? io_r_449_b : _GEN_19288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19290 = 10'h1c2 == r_count_25_io_out ? io_r_450_b : _GEN_19289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19291 = 10'h1c3 == r_count_25_io_out ? io_r_451_b : _GEN_19290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19292 = 10'h1c4 == r_count_25_io_out ? io_r_452_b : _GEN_19291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19293 = 10'h1c5 == r_count_25_io_out ? io_r_453_b : _GEN_19292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19294 = 10'h1c6 == r_count_25_io_out ? io_r_454_b : _GEN_19293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19295 = 10'h1c7 == r_count_25_io_out ? io_r_455_b : _GEN_19294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19296 = 10'h1c8 == r_count_25_io_out ? io_r_456_b : _GEN_19295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19297 = 10'h1c9 == r_count_25_io_out ? io_r_457_b : _GEN_19296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19298 = 10'h1ca == r_count_25_io_out ? io_r_458_b : _GEN_19297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19299 = 10'h1cb == r_count_25_io_out ? io_r_459_b : _GEN_19298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19300 = 10'h1cc == r_count_25_io_out ? io_r_460_b : _GEN_19299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19301 = 10'h1cd == r_count_25_io_out ? io_r_461_b : _GEN_19300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19302 = 10'h1ce == r_count_25_io_out ? io_r_462_b : _GEN_19301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19303 = 10'h1cf == r_count_25_io_out ? io_r_463_b : _GEN_19302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19304 = 10'h1d0 == r_count_25_io_out ? io_r_464_b : _GEN_19303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19305 = 10'h1d1 == r_count_25_io_out ? io_r_465_b : _GEN_19304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19306 = 10'h1d2 == r_count_25_io_out ? io_r_466_b : _GEN_19305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19307 = 10'h1d3 == r_count_25_io_out ? io_r_467_b : _GEN_19306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19308 = 10'h1d4 == r_count_25_io_out ? io_r_468_b : _GEN_19307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19309 = 10'h1d5 == r_count_25_io_out ? io_r_469_b : _GEN_19308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19310 = 10'h1d6 == r_count_25_io_out ? io_r_470_b : _GEN_19309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19311 = 10'h1d7 == r_count_25_io_out ? io_r_471_b : _GEN_19310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19312 = 10'h1d8 == r_count_25_io_out ? io_r_472_b : _GEN_19311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19313 = 10'h1d9 == r_count_25_io_out ? io_r_473_b : _GEN_19312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19314 = 10'h1da == r_count_25_io_out ? io_r_474_b : _GEN_19313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19315 = 10'h1db == r_count_25_io_out ? io_r_475_b : _GEN_19314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19316 = 10'h1dc == r_count_25_io_out ? io_r_476_b : _GEN_19315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19317 = 10'h1dd == r_count_25_io_out ? io_r_477_b : _GEN_19316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19318 = 10'h1de == r_count_25_io_out ? io_r_478_b : _GEN_19317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19319 = 10'h1df == r_count_25_io_out ? io_r_479_b : _GEN_19318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19320 = 10'h1e0 == r_count_25_io_out ? io_r_480_b : _GEN_19319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19321 = 10'h1e1 == r_count_25_io_out ? io_r_481_b : _GEN_19320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19322 = 10'h1e2 == r_count_25_io_out ? io_r_482_b : _GEN_19321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19323 = 10'h1e3 == r_count_25_io_out ? io_r_483_b : _GEN_19322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19324 = 10'h1e4 == r_count_25_io_out ? io_r_484_b : _GEN_19323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19325 = 10'h1e5 == r_count_25_io_out ? io_r_485_b : _GEN_19324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19326 = 10'h1e6 == r_count_25_io_out ? io_r_486_b : _GEN_19325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19327 = 10'h1e7 == r_count_25_io_out ? io_r_487_b : _GEN_19326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19328 = 10'h1e8 == r_count_25_io_out ? io_r_488_b : _GEN_19327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19329 = 10'h1e9 == r_count_25_io_out ? io_r_489_b : _GEN_19328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19330 = 10'h1ea == r_count_25_io_out ? io_r_490_b : _GEN_19329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19331 = 10'h1eb == r_count_25_io_out ? io_r_491_b : _GEN_19330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19332 = 10'h1ec == r_count_25_io_out ? io_r_492_b : _GEN_19331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19333 = 10'h1ed == r_count_25_io_out ? io_r_493_b : _GEN_19332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19334 = 10'h1ee == r_count_25_io_out ? io_r_494_b : _GEN_19333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19335 = 10'h1ef == r_count_25_io_out ? io_r_495_b : _GEN_19334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19336 = 10'h1f0 == r_count_25_io_out ? io_r_496_b : _GEN_19335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19337 = 10'h1f1 == r_count_25_io_out ? io_r_497_b : _GEN_19336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19338 = 10'h1f2 == r_count_25_io_out ? io_r_498_b : _GEN_19337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19339 = 10'h1f3 == r_count_25_io_out ? io_r_499_b : _GEN_19338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19340 = 10'h1f4 == r_count_25_io_out ? io_r_500_b : _GEN_19339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19341 = 10'h1f5 == r_count_25_io_out ? io_r_501_b : _GEN_19340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19342 = 10'h1f6 == r_count_25_io_out ? io_r_502_b : _GEN_19341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19343 = 10'h1f7 == r_count_25_io_out ? io_r_503_b : _GEN_19342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19344 = 10'h1f8 == r_count_25_io_out ? io_r_504_b : _GEN_19343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19345 = 10'h1f9 == r_count_25_io_out ? io_r_505_b : _GEN_19344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19346 = 10'h1fa == r_count_25_io_out ? io_r_506_b : _GEN_19345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19347 = 10'h1fb == r_count_25_io_out ? io_r_507_b : _GEN_19346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19348 = 10'h1fc == r_count_25_io_out ? io_r_508_b : _GEN_19347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19349 = 10'h1fd == r_count_25_io_out ? io_r_509_b : _GEN_19348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19350 = 10'h1fe == r_count_25_io_out ? io_r_510_b : _GEN_19349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19351 = 10'h1ff == r_count_25_io_out ? io_r_511_b : _GEN_19350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19352 = 10'h200 == r_count_25_io_out ? io_r_512_b : _GEN_19351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19353 = 10'h201 == r_count_25_io_out ? io_r_513_b : _GEN_19352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19354 = 10'h202 == r_count_25_io_out ? io_r_514_b : _GEN_19353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19355 = 10'h203 == r_count_25_io_out ? io_r_515_b : _GEN_19354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19356 = 10'h204 == r_count_25_io_out ? io_r_516_b : _GEN_19355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19357 = 10'h205 == r_count_25_io_out ? io_r_517_b : _GEN_19356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19358 = 10'h206 == r_count_25_io_out ? io_r_518_b : _GEN_19357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19359 = 10'h207 == r_count_25_io_out ? io_r_519_b : _GEN_19358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19360 = 10'h208 == r_count_25_io_out ? io_r_520_b : _GEN_19359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19361 = 10'h209 == r_count_25_io_out ? io_r_521_b : _GEN_19360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19362 = 10'h20a == r_count_25_io_out ? io_r_522_b : _GEN_19361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19363 = 10'h20b == r_count_25_io_out ? io_r_523_b : _GEN_19362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19364 = 10'h20c == r_count_25_io_out ? io_r_524_b : _GEN_19363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19365 = 10'h20d == r_count_25_io_out ? io_r_525_b : _GEN_19364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19366 = 10'h20e == r_count_25_io_out ? io_r_526_b : _GEN_19365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19367 = 10'h20f == r_count_25_io_out ? io_r_527_b : _GEN_19366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19368 = 10'h210 == r_count_25_io_out ? io_r_528_b : _GEN_19367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19369 = 10'h211 == r_count_25_io_out ? io_r_529_b : _GEN_19368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19370 = 10'h212 == r_count_25_io_out ? io_r_530_b : _GEN_19369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19371 = 10'h213 == r_count_25_io_out ? io_r_531_b : _GEN_19370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19372 = 10'h214 == r_count_25_io_out ? io_r_532_b : _GEN_19371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19373 = 10'h215 == r_count_25_io_out ? io_r_533_b : _GEN_19372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19374 = 10'h216 == r_count_25_io_out ? io_r_534_b : _GEN_19373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19375 = 10'h217 == r_count_25_io_out ? io_r_535_b : _GEN_19374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19376 = 10'h218 == r_count_25_io_out ? io_r_536_b : _GEN_19375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19377 = 10'h219 == r_count_25_io_out ? io_r_537_b : _GEN_19376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19378 = 10'h21a == r_count_25_io_out ? io_r_538_b : _GEN_19377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19379 = 10'h21b == r_count_25_io_out ? io_r_539_b : _GEN_19378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19380 = 10'h21c == r_count_25_io_out ? io_r_540_b : _GEN_19379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19381 = 10'h21d == r_count_25_io_out ? io_r_541_b : _GEN_19380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19382 = 10'h21e == r_count_25_io_out ? io_r_542_b : _GEN_19381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19383 = 10'h21f == r_count_25_io_out ? io_r_543_b : _GEN_19382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19384 = 10'h220 == r_count_25_io_out ? io_r_544_b : _GEN_19383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19385 = 10'h221 == r_count_25_io_out ? io_r_545_b : _GEN_19384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19386 = 10'h222 == r_count_25_io_out ? io_r_546_b : _GEN_19385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19387 = 10'h223 == r_count_25_io_out ? io_r_547_b : _GEN_19386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19388 = 10'h224 == r_count_25_io_out ? io_r_548_b : _GEN_19387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19389 = 10'h225 == r_count_25_io_out ? io_r_549_b : _GEN_19388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19390 = 10'h226 == r_count_25_io_out ? io_r_550_b : _GEN_19389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19391 = 10'h227 == r_count_25_io_out ? io_r_551_b : _GEN_19390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19392 = 10'h228 == r_count_25_io_out ? io_r_552_b : _GEN_19391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19393 = 10'h229 == r_count_25_io_out ? io_r_553_b : _GEN_19392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19394 = 10'h22a == r_count_25_io_out ? io_r_554_b : _GEN_19393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19395 = 10'h22b == r_count_25_io_out ? io_r_555_b : _GEN_19394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19396 = 10'h22c == r_count_25_io_out ? io_r_556_b : _GEN_19395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19397 = 10'h22d == r_count_25_io_out ? io_r_557_b : _GEN_19396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19398 = 10'h22e == r_count_25_io_out ? io_r_558_b : _GEN_19397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19399 = 10'h22f == r_count_25_io_out ? io_r_559_b : _GEN_19398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19400 = 10'h230 == r_count_25_io_out ? io_r_560_b : _GEN_19399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19401 = 10'h231 == r_count_25_io_out ? io_r_561_b : _GEN_19400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19402 = 10'h232 == r_count_25_io_out ? io_r_562_b : _GEN_19401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19403 = 10'h233 == r_count_25_io_out ? io_r_563_b : _GEN_19402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19404 = 10'h234 == r_count_25_io_out ? io_r_564_b : _GEN_19403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19405 = 10'h235 == r_count_25_io_out ? io_r_565_b : _GEN_19404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19406 = 10'h236 == r_count_25_io_out ? io_r_566_b : _GEN_19405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19407 = 10'h237 == r_count_25_io_out ? io_r_567_b : _GEN_19406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19408 = 10'h238 == r_count_25_io_out ? io_r_568_b : _GEN_19407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19409 = 10'h239 == r_count_25_io_out ? io_r_569_b : _GEN_19408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19410 = 10'h23a == r_count_25_io_out ? io_r_570_b : _GEN_19409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19411 = 10'h23b == r_count_25_io_out ? io_r_571_b : _GEN_19410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19412 = 10'h23c == r_count_25_io_out ? io_r_572_b : _GEN_19411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19413 = 10'h23d == r_count_25_io_out ? io_r_573_b : _GEN_19412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19414 = 10'h23e == r_count_25_io_out ? io_r_574_b : _GEN_19413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19415 = 10'h23f == r_count_25_io_out ? io_r_575_b : _GEN_19414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19416 = 10'h240 == r_count_25_io_out ? io_r_576_b : _GEN_19415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19417 = 10'h241 == r_count_25_io_out ? io_r_577_b : _GEN_19416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19418 = 10'h242 == r_count_25_io_out ? io_r_578_b : _GEN_19417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19419 = 10'h243 == r_count_25_io_out ? io_r_579_b : _GEN_19418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19420 = 10'h244 == r_count_25_io_out ? io_r_580_b : _GEN_19419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19421 = 10'h245 == r_count_25_io_out ? io_r_581_b : _GEN_19420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19422 = 10'h246 == r_count_25_io_out ? io_r_582_b : _GEN_19421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19423 = 10'h247 == r_count_25_io_out ? io_r_583_b : _GEN_19422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19424 = 10'h248 == r_count_25_io_out ? io_r_584_b : _GEN_19423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19425 = 10'h249 == r_count_25_io_out ? io_r_585_b : _GEN_19424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19426 = 10'h24a == r_count_25_io_out ? io_r_586_b : _GEN_19425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19427 = 10'h24b == r_count_25_io_out ? io_r_587_b : _GEN_19426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19428 = 10'h24c == r_count_25_io_out ? io_r_588_b : _GEN_19427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19429 = 10'h24d == r_count_25_io_out ? io_r_589_b : _GEN_19428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19430 = 10'h24e == r_count_25_io_out ? io_r_590_b : _GEN_19429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19431 = 10'h24f == r_count_25_io_out ? io_r_591_b : _GEN_19430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19432 = 10'h250 == r_count_25_io_out ? io_r_592_b : _GEN_19431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19433 = 10'h251 == r_count_25_io_out ? io_r_593_b : _GEN_19432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19434 = 10'h252 == r_count_25_io_out ? io_r_594_b : _GEN_19433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19435 = 10'h253 == r_count_25_io_out ? io_r_595_b : _GEN_19434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19436 = 10'h254 == r_count_25_io_out ? io_r_596_b : _GEN_19435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19437 = 10'h255 == r_count_25_io_out ? io_r_597_b : _GEN_19436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19438 = 10'h256 == r_count_25_io_out ? io_r_598_b : _GEN_19437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19439 = 10'h257 == r_count_25_io_out ? io_r_599_b : _GEN_19438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19440 = 10'h258 == r_count_25_io_out ? io_r_600_b : _GEN_19439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19441 = 10'h259 == r_count_25_io_out ? io_r_601_b : _GEN_19440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19442 = 10'h25a == r_count_25_io_out ? io_r_602_b : _GEN_19441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19443 = 10'h25b == r_count_25_io_out ? io_r_603_b : _GEN_19442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19444 = 10'h25c == r_count_25_io_out ? io_r_604_b : _GEN_19443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19445 = 10'h25d == r_count_25_io_out ? io_r_605_b : _GEN_19444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19446 = 10'h25e == r_count_25_io_out ? io_r_606_b : _GEN_19445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19447 = 10'h25f == r_count_25_io_out ? io_r_607_b : _GEN_19446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19448 = 10'h260 == r_count_25_io_out ? io_r_608_b : _GEN_19447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19449 = 10'h261 == r_count_25_io_out ? io_r_609_b : _GEN_19448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19450 = 10'h262 == r_count_25_io_out ? io_r_610_b : _GEN_19449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19451 = 10'h263 == r_count_25_io_out ? io_r_611_b : _GEN_19450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19452 = 10'h264 == r_count_25_io_out ? io_r_612_b : _GEN_19451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19453 = 10'h265 == r_count_25_io_out ? io_r_613_b : _GEN_19452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19454 = 10'h266 == r_count_25_io_out ? io_r_614_b : _GEN_19453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19455 = 10'h267 == r_count_25_io_out ? io_r_615_b : _GEN_19454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19456 = 10'h268 == r_count_25_io_out ? io_r_616_b : _GEN_19455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19457 = 10'h269 == r_count_25_io_out ? io_r_617_b : _GEN_19456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19458 = 10'h26a == r_count_25_io_out ? io_r_618_b : _GEN_19457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19459 = 10'h26b == r_count_25_io_out ? io_r_619_b : _GEN_19458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19460 = 10'h26c == r_count_25_io_out ? io_r_620_b : _GEN_19459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19461 = 10'h26d == r_count_25_io_out ? io_r_621_b : _GEN_19460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19462 = 10'h26e == r_count_25_io_out ? io_r_622_b : _GEN_19461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19463 = 10'h26f == r_count_25_io_out ? io_r_623_b : _GEN_19462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19464 = 10'h270 == r_count_25_io_out ? io_r_624_b : _GEN_19463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19465 = 10'h271 == r_count_25_io_out ? io_r_625_b : _GEN_19464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19466 = 10'h272 == r_count_25_io_out ? io_r_626_b : _GEN_19465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19467 = 10'h273 == r_count_25_io_out ? io_r_627_b : _GEN_19466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19468 = 10'h274 == r_count_25_io_out ? io_r_628_b : _GEN_19467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19469 = 10'h275 == r_count_25_io_out ? io_r_629_b : _GEN_19468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19470 = 10'h276 == r_count_25_io_out ? io_r_630_b : _GEN_19469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19471 = 10'h277 == r_count_25_io_out ? io_r_631_b : _GEN_19470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19472 = 10'h278 == r_count_25_io_out ? io_r_632_b : _GEN_19471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19473 = 10'h279 == r_count_25_io_out ? io_r_633_b : _GEN_19472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19474 = 10'h27a == r_count_25_io_out ? io_r_634_b : _GEN_19473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19475 = 10'h27b == r_count_25_io_out ? io_r_635_b : _GEN_19474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19476 = 10'h27c == r_count_25_io_out ? io_r_636_b : _GEN_19475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19477 = 10'h27d == r_count_25_io_out ? io_r_637_b : _GEN_19476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19478 = 10'h27e == r_count_25_io_out ? io_r_638_b : _GEN_19477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19479 = 10'h27f == r_count_25_io_out ? io_r_639_b : _GEN_19478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19480 = 10'h280 == r_count_25_io_out ? io_r_640_b : _GEN_19479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19481 = 10'h281 == r_count_25_io_out ? io_r_641_b : _GEN_19480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19482 = 10'h282 == r_count_25_io_out ? io_r_642_b : _GEN_19481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19483 = 10'h283 == r_count_25_io_out ? io_r_643_b : _GEN_19482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19484 = 10'h284 == r_count_25_io_out ? io_r_644_b : _GEN_19483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19485 = 10'h285 == r_count_25_io_out ? io_r_645_b : _GEN_19484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19486 = 10'h286 == r_count_25_io_out ? io_r_646_b : _GEN_19485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19487 = 10'h287 == r_count_25_io_out ? io_r_647_b : _GEN_19486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19488 = 10'h288 == r_count_25_io_out ? io_r_648_b : _GEN_19487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19489 = 10'h289 == r_count_25_io_out ? io_r_649_b : _GEN_19488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19490 = 10'h28a == r_count_25_io_out ? io_r_650_b : _GEN_19489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19491 = 10'h28b == r_count_25_io_out ? io_r_651_b : _GEN_19490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19492 = 10'h28c == r_count_25_io_out ? io_r_652_b : _GEN_19491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19493 = 10'h28d == r_count_25_io_out ? io_r_653_b : _GEN_19492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19494 = 10'h28e == r_count_25_io_out ? io_r_654_b : _GEN_19493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19495 = 10'h28f == r_count_25_io_out ? io_r_655_b : _GEN_19494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19496 = 10'h290 == r_count_25_io_out ? io_r_656_b : _GEN_19495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19497 = 10'h291 == r_count_25_io_out ? io_r_657_b : _GEN_19496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19498 = 10'h292 == r_count_25_io_out ? io_r_658_b : _GEN_19497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19499 = 10'h293 == r_count_25_io_out ? io_r_659_b : _GEN_19498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19500 = 10'h294 == r_count_25_io_out ? io_r_660_b : _GEN_19499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19501 = 10'h295 == r_count_25_io_out ? io_r_661_b : _GEN_19500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19502 = 10'h296 == r_count_25_io_out ? io_r_662_b : _GEN_19501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19503 = 10'h297 == r_count_25_io_out ? io_r_663_b : _GEN_19502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19504 = 10'h298 == r_count_25_io_out ? io_r_664_b : _GEN_19503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19505 = 10'h299 == r_count_25_io_out ? io_r_665_b : _GEN_19504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19506 = 10'h29a == r_count_25_io_out ? io_r_666_b : _GEN_19505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19507 = 10'h29b == r_count_25_io_out ? io_r_667_b : _GEN_19506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19508 = 10'h29c == r_count_25_io_out ? io_r_668_b : _GEN_19507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19509 = 10'h29d == r_count_25_io_out ? io_r_669_b : _GEN_19508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19510 = 10'h29e == r_count_25_io_out ? io_r_670_b : _GEN_19509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19511 = 10'h29f == r_count_25_io_out ? io_r_671_b : _GEN_19510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19512 = 10'h2a0 == r_count_25_io_out ? io_r_672_b : _GEN_19511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19513 = 10'h2a1 == r_count_25_io_out ? io_r_673_b : _GEN_19512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19514 = 10'h2a2 == r_count_25_io_out ? io_r_674_b : _GEN_19513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19515 = 10'h2a3 == r_count_25_io_out ? io_r_675_b : _GEN_19514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19516 = 10'h2a4 == r_count_25_io_out ? io_r_676_b : _GEN_19515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19517 = 10'h2a5 == r_count_25_io_out ? io_r_677_b : _GEN_19516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19518 = 10'h2a6 == r_count_25_io_out ? io_r_678_b : _GEN_19517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19519 = 10'h2a7 == r_count_25_io_out ? io_r_679_b : _GEN_19518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19520 = 10'h2a8 == r_count_25_io_out ? io_r_680_b : _GEN_19519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19521 = 10'h2a9 == r_count_25_io_out ? io_r_681_b : _GEN_19520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19522 = 10'h2aa == r_count_25_io_out ? io_r_682_b : _GEN_19521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19523 = 10'h2ab == r_count_25_io_out ? io_r_683_b : _GEN_19522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19524 = 10'h2ac == r_count_25_io_out ? io_r_684_b : _GEN_19523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19525 = 10'h2ad == r_count_25_io_out ? io_r_685_b : _GEN_19524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19526 = 10'h2ae == r_count_25_io_out ? io_r_686_b : _GEN_19525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19527 = 10'h2af == r_count_25_io_out ? io_r_687_b : _GEN_19526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19528 = 10'h2b0 == r_count_25_io_out ? io_r_688_b : _GEN_19527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19529 = 10'h2b1 == r_count_25_io_out ? io_r_689_b : _GEN_19528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19530 = 10'h2b2 == r_count_25_io_out ? io_r_690_b : _GEN_19529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19531 = 10'h2b3 == r_count_25_io_out ? io_r_691_b : _GEN_19530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19532 = 10'h2b4 == r_count_25_io_out ? io_r_692_b : _GEN_19531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19533 = 10'h2b5 == r_count_25_io_out ? io_r_693_b : _GEN_19532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19534 = 10'h2b6 == r_count_25_io_out ? io_r_694_b : _GEN_19533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19535 = 10'h2b7 == r_count_25_io_out ? io_r_695_b : _GEN_19534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19536 = 10'h2b8 == r_count_25_io_out ? io_r_696_b : _GEN_19535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19537 = 10'h2b9 == r_count_25_io_out ? io_r_697_b : _GEN_19536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19538 = 10'h2ba == r_count_25_io_out ? io_r_698_b : _GEN_19537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19539 = 10'h2bb == r_count_25_io_out ? io_r_699_b : _GEN_19538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19540 = 10'h2bc == r_count_25_io_out ? io_r_700_b : _GEN_19539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19541 = 10'h2bd == r_count_25_io_out ? io_r_701_b : _GEN_19540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19542 = 10'h2be == r_count_25_io_out ? io_r_702_b : _GEN_19541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19543 = 10'h2bf == r_count_25_io_out ? io_r_703_b : _GEN_19542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19544 = 10'h2c0 == r_count_25_io_out ? io_r_704_b : _GEN_19543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19545 = 10'h2c1 == r_count_25_io_out ? io_r_705_b : _GEN_19544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19546 = 10'h2c2 == r_count_25_io_out ? io_r_706_b : _GEN_19545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19547 = 10'h2c3 == r_count_25_io_out ? io_r_707_b : _GEN_19546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19548 = 10'h2c4 == r_count_25_io_out ? io_r_708_b : _GEN_19547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19549 = 10'h2c5 == r_count_25_io_out ? io_r_709_b : _GEN_19548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19550 = 10'h2c6 == r_count_25_io_out ? io_r_710_b : _GEN_19549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19551 = 10'h2c7 == r_count_25_io_out ? io_r_711_b : _GEN_19550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19552 = 10'h2c8 == r_count_25_io_out ? io_r_712_b : _GEN_19551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19553 = 10'h2c9 == r_count_25_io_out ? io_r_713_b : _GEN_19552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19554 = 10'h2ca == r_count_25_io_out ? io_r_714_b : _GEN_19553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19555 = 10'h2cb == r_count_25_io_out ? io_r_715_b : _GEN_19554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19556 = 10'h2cc == r_count_25_io_out ? io_r_716_b : _GEN_19555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19557 = 10'h2cd == r_count_25_io_out ? io_r_717_b : _GEN_19556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19558 = 10'h2ce == r_count_25_io_out ? io_r_718_b : _GEN_19557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19559 = 10'h2cf == r_count_25_io_out ? io_r_719_b : _GEN_19558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19560 = 10'h2d0 == r_count_25_io_out ? io_r_720_b : _GEN_19559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19561 = 10'h2d1 == r_count_25_io_out ? io_r_721_b : _GEN_19560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19562 = 10'h2d2 == r_count_25_io_out ? io_r_722_b : _GEN_19561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19563 = 10'h2d3 == r_count_25_io_out ? io_r_723_b : _GEN_19562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19564 = 10'h2d4 == r_count_25_io_out ? io_r_724_b : _GEN_19563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19565 = 10'h2d5 == r_count_25_io_out ? io_r_725_b : _GEN_19564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19566 = 10'h2d6 == r_count_25_io_out ? io_r_726_b : _GEN_19565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19567 = 10'h2d7 == r_count_25_io_out ? io_r_727_b : _GEN_19566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19568 = 10'h2d8 == r_count_25_io_out ? io_r_728_b : _GEN_19567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19569 = 10'h2d9 == r_count_25_io_out ? io_r_729_b : _GEN_19568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19570 = 10'h2da == r_count_25_io_out ? io_r_730_b : _GEN_19569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19571 = 10'h2db == r_count_25_io_out ? io_r_731_b : _GEN_19570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19572 = 10'h2dc == r_count_25_io_out ? io_r_732_b : _GEN_19571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19573 = 10'h2dd == r_count_25_io_out ? io_r_733_b : _GEN_19572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19574 = 10'h2de == r_count_25_io_out ? io_r_734_b : _GEN_19573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19575 = 10'h2df == r_count_25_io_out ? io_r_735_b : _GEN_19574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19576 = 10'h2e0 == r_count_25_io_out ? io_r_736_b : _GEN_19575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19577 = 10'h2e1 == r_count_25_io_out ? io_r_737_b : _GEN_19576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19578 = 10'h2e2 == r_count_25_io_out ? io_r_738_b : _GEN_19577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19579 = 10'h2e3 == r_count_25_io_out ? io_r_739_b : _GEN_19578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19580 = 10'h2e4 == r_count_25_io_out ? io_r_740_b : _GEN_19579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19581 = 10'h2e5 == r_count_25_io_out ? io_r_741_b : _GEN_19580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19582 = 10'h2e6 == r_count_25_io_out ? io_r_742_b : _GEN_19581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19583 = 10'h2e7 == r_count_25_io_out ? io_r_743_b : _GEN_19582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19584 = 10'h2e8 == r_count_25_io_out ? io_r_744_b : _GEN_19583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19585 = 10'h2e9 == r_count_25_io_out ? io_r_745_b : _GEN_19584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19586 = 10'h2ea == r_count_25_io_out ? io_r_746_b : _GEN_19585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19587 = 10'h2eb == r_count_25_io_out ? io_r_747_b : _GEN_19586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19588 = 10'h2ec == r_count_25_io_out ? io_r_748_b : _GEN_19587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19591 = 10'h1 == r_count_26_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19592 = 10'h2 == r_count_26_io_out ? io_r_2_b : _GEN_19591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19593 = 10'h3 == r_count_26_io_out ? io_r_3_b : _GEN_19592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19594 = 10'h4 == r_count_26_io_out ? io_r_4_b : _GEN_19593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19595 = 10'h5 == r_count_26_io_out ? io_r_5_b : _GEN_19594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19596 = 10'h6 == r_count_26_io_out ? io_r_6_b : _GEN_19595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19597 = 10'h7 == r_count_26_io_out ? io_r_7_b : _GEN_19596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19598 = 10'h8 == r_count_26_io_out ? io_r_8_b : _GEN_19597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19599 = 10'h9 == r_count_26_io_out ? io_r_9_b : _GEN_19598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19600 = 10'ha == r_count_26_io_out ? io_r_10_b : _GEN_19599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19601 = 10'hb == r_count_26_io_out ? io_r_11_b : _GEN_19600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19602 = 10'hc == r_count_26_io_out ? io_r_12_b : _GEN_19601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19603 = 10'hd == r_count_26_io_out ? io_r_13_b : _GEN_19602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19604 = 10'he == r_count_26_io_out ? io_r_14_b : _GEN_19603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19605 = 10'hf == r_count_26_io_out ? io_r_15_b : _GEN_19604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19606 = 10'h10 == r_count_26_io_out ? io_r_16_b : _GEN_19605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19607 = 10'h11 == r_count_26_io_out ? io_r_17_b : _GEN_19606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19608 = 10'h12 == r_count_26_io_out ? io_r_18_b : _GEN_19607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19609 = 10'h13 == r_count_26_io_out ? io_r_19_b : _GEN_19608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19610 = 10'h14 == r_count_26_io_out ? io_r_20_b : _GEN_19609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19611 = 10'h15 == r_count_26_io_out ? io_r_21_b : _GEN_19610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19612 = 10'h16 == r_count_26_io_out ? io_r_22_b : _GEN_19611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19613 = 10'h17 == r_count_26_io_out ? io_r_23_b : _GEN_19612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19614 = 10'h18 == r_count_26_io_out ? io_r_24_b : _GEN_19613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19615 = 10'h19 == r_count_26_io_out ? io_r_25_b : _GEN_19614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19616 = 10'h1a == r_count_26_io_out ? io_r_26_b : _GEN_19615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19617 = 10'h1b == r_count_26_io_out ? io_r_27_b : _GEN_19616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19618 = 10'h1c == r_count_26_io_out ? io_r_28_b : _GEN_19617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19619 = 10'h1d == r_count_26_io_out ? io_r_29_b : _GEN_19618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19620 = 10'h1e == r_count_26_io_out ? io_r_30_b : _GEN_19619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19621 = 10'h1f == r_count_26_io_out ? io_r_31_b : _GEN_19620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19622 = 10'h20 == r_count_26_io_out ? io_r_32_b : _GEN_19621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19623 = 10'h21 == r_count_26_io_out ? io_r_33_b : _GEN_19622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19624 = 10'h22 == r_count_26_io_out ? io_r_34_b : _GEN_19623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19625 = 10'h23 == r_count_26_io_out ? io_r_35_b : _GEN_19624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19626 = 10'h24 == r_count_26_io_out ? io_r_36_b : _GEN_19625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19627 = 10'h25 == r_count_26_io_out ? io_r_37_b : _GEN_19626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19628 = 10'h26 == r_count_26_io_out ? io_r_38_b : _GEN_19627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19629 = 10'h27 == r_count_26_io_out ? io_r_39_b : _GEN_19628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19630 = 10'h28 == r_count_26_io_out ? io_r_40_b : _GEN_19629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19631 = 10'h29 == r_count_26_io_out ? io_r_41_b : _GEN_19630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19632 = 10'h2a == r_count_26_io_out ? io_r_42_b : _GEN_19631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19633 = 10'h2b == r_count_26_io_out ? io_r_43_b : _GEN_19632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19634 = 10'h2c == r_count_26_io_out ? io_r_44_b : _GEN_19633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19635 = 10'h2d == r_count_26_io_out ? io_r_45_b : _GEN_19634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19636 = 10'h2e == r_count_26_io_out ? io_r_46_b : _GEN_19635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19637 = 10'h2f == r_count_26_io_out ? io_r_47_b : _GEN_19636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19638 = 10'h30 == r_count_26_io_out ? io_r_48_b : _GEN_19637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19639 = 10'h31 == r_count_26_io_out ? io_r_49_b : _GEN_19638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19640 = 10'h32 == r_count_26_io_out ? io_r_50_b : _GEN_19639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19641 = 10'h33 == r_count_26_io_out ? io_r_51_b : _GEN_19640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19642 = 10'h34 == r_count_26_io_out ? io_r_52_b : _GEN_19641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19643 = 10'h35 == r_count_26_io_out ? io_r_53_b : _GEN_19642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19644 = 10'h36 == r_count_26_io_out ? io_r_54_b : _GEN_19643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19645 = 10'h37 == r_count_26_io_out ? io_r_55_b : _GEN_19644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19646 = 10'h38 == r_count_26_io_out ? io_r_56_b : _GEN_19645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19647 = 10'h39 == r_count_26_io_out ? io_r_57_b : _GEN_19646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19648 = 10'h3a == r_count_26_io_out ? io_r_58_b : _GEN_19647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19649 = 10'h3b == r_count_26_io_out ? io_r_59_b : _GEN_19648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19650 = 10'h3c == r_count_26_io_out ? io_r_60_b : _GEN_19649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19651 = 10'h3d == r_count_26_io_out ? io_r_61_b : _GEN_19650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19652 = 10'h3e == r_count_26_io_out ? io_r_62_b : _GEN_19651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19653 = 10'h3f == r_count_26_io_out ? io_r_63_b : _GEN_19652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19654 = 10'h40 == r_count_26_io_out ? io_r_64_b : _GEN_19653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19655 = 10'h41 == r_count_26_io_out ? io_r_65_b : _GEN_19654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19656 = 10'h42 == r_count_26_io_out ? io_r_66_b : _GEN_19655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19657 = 10'h43 == r_count_26_io_out ? io_r_67_b : _GEN_19656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19658 = 10'h44 == r_count_26_io_out ? io_r_68_b : _GEN_19657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19659 = 10'h45 == r_count_26_io_out ? io_r_69_b : _GEN_19658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19660 = 10'h46 == r_count_26_io_out ? io_r_70_b : _GEN_19659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19661 = 10'h47 == r_count_26_io_out ? io_r_71_b : _GEN_19660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19662 = 10'h48 == r_count_26_io_out ? io_r_72_b : _GEN_19661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19663 = 10'h49 == r_count_26_io_out ? io_r_73_b : _GEN_19662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19664 = 10'h4a == r_count_26_io_out ? io_r_74_b : _GEN_19663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19665 = 10'h4b == r_count_26_io_out ? io_r_75_b : _GEN_19664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19666 = 10'h4c == r_count_26_io_out ? io_r_76_b : _GEN_19665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19667 = 10'h4d == r_count_26_io_out ? io_r_77_b : _GEN_19666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19668 = 10'h4e == r_count_26_io_out ? io_r_78_b : _GEN_19667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19669 = 10'h4f == r_count_26_io_out ? io_r_79_b : _GEN_19668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19670 = 10'h50 == r_count_26_io_out ? io_r_80_b : _GEN_19669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19671 = 10'h51 == r_count_26_io_out ? io_r_81_b : _GEN_19670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19672 = 10'h52 == r_count_26_io_out ? io_r_82_b : _GEN_19671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19673 = 10'h53 == r_count_26_io_out ? io_r_83_b : _GEN_19672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19674 = 10'h54 == r_count_26_io_out ? io_r_84_b : _GEN_19673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19675 = 10'h55 == r_count_26_io_out ? io_r_85_b : _GEN_19674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19676 = 10'h56 == r_count_26_io_out ? io_r_86_b : _GEN_19675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19677 = 10'h57 == r_count_26_io_out ? io_r_87_b : _GEN_19676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19678 = 10'h58 == r_count_26_io_out ? io_r_88_b : _GEN_19677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19679 = 10'h59 == r_count_26_io_out ? io_r_89_b : _GEN_19678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19680 = 10'h5a == r_count_26_io_out ? io_r_90_b : _GEN_19679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19681 = 10'h5b == r_count_26_io_out ? io_r_91_b : _GEN_19680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19682 = 10'h5c == r_count_26_io_out ? io_r_92_b : _GEN_19681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19683 = 10'h5d == r_count_26_io_out ? io_r_93_b : _GEN_19682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19684 = 10'h5e == r_count_26_io_out ? io_r_94_b : _GEN_19683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19685 = 10'h5f == r_count_26_io_out ? io_r_95_b : _GEN_19684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19686 = 10'h60 == r_count_26_io_out ? io_r_96_b : _GEN_19685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19687 = 10'h61 == r_count_26_io_out ? io_r_97_b : _GEN_19686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19688 = 10'h62 == r_count_26_io_out ? io_r_98_b : _GEN_19687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19689 = 10'h63 == r_count_26_io_out ? io_r_99_b : _GEN_19688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19690 = 10'h64 == r_count_26_io_out ? io_r_100_b : _GEN_19689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19691 = 10'h65 == r_count_26_io_out ? io_r_101_b : _GEN_19690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19692 = 10'h66 == r_count_26_io_out ? io_r_102_b : _GEN_19691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19693 = 10'h67 == r_count_26_io_out ? io_r_103_b : _GEN_19692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19694 = 10'h68 == r_count_26_io_out ? io_r_104_b : _GEN_19693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19695 = 10'h69 == r_count_26_io_out ? io_r_105_b : _GEN_19694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19696 = 10'h6a == r_count_26_io_out ? io_r_106_b : _GEN_19695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19697 = 10'h6b == r_count_26_io_out ? io_r_107_b : _GEN_19696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19698 = 10'h6c == r_count_26_io_out ? io_r_108_b : _GEN_19697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19699 = 10'h6d == r_count_26_io_out ? io_r_109_b : _GEN_19698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19700 = 10'h6e == r_count_26_io_out ? io_r_110_b : _GEN_19699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19701 = 10'h6f == r_count_26_io_out ? io_r_111_b : _GEN_19700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19702 = 10'h70 == r_count_26_io_out ? io_r_112_b : _GEN_19701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19703 = 10'h71 == r_count_26_io_out ? io_r_113_b : _GEN_19702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19704 = 10'h72 == r_count_26_io_out ? io_r_114_b : _GEN_19703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19705 = 10'h73 == r_count_26_io_out ? io_r_115_b : _GEN_19704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19706 = 10'h74 == r_count_26_io_out ? io_r_116_b : _GEN_19705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19707 = 10'h75 == r_count_26_io_out ? io_r_117_b : _GEN_19706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19708 = 10'h76 == r_count_26_io_out ? io_r_118_b : _GEN_19707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19709 = 10'h77 == r_count_26_io_out ? io_r_119_b : _GEN_19708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19710 = 10'h78 == r_count_26_io_out ? io_r_120_b : _GEN_19709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19711 = 10'h79 == r_count_26_io_out ? io_r_121_b : _GEN_19710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19712 = 10'h7a == r_count_26_io_out ? io_r_122_b : _GEN_19711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19713 = 10'h7b == r_count_26_io_out ? io_r_123_b : _GEN_19712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19714 = 10'h7c == r_count_26_io_out ? io_r_124_b : _GEN_19713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19715 = 10'h7d == r_count_26_io_out ? io_r_125_b : _GEN_19714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19716 = 10'h7e == r_count_26_io_out ? io_r_126_b : _GEN_19715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19717 = 10'h7f == r_count_26_io_out ? io_r_127_b : _GEN_19716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19718 = 10'h80 == r_count_26_io_out ? io_r_128_b : _GEN_19717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19719 = 10'h81 == r_count_26_io_out ? io_r_129_b : _GEN_19718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19720 = 10'h82 == r_count_26_io_out ? io_r_130_b : _GEN_19719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19721 = 10'h83 == r_count_26_io_out ? io_r_131_b : _GEN_19720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19722 = 10'h84 == r_count_26_io_out ? io_r_132_b : _GEN_19721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19723 = 10'h85 == r_count_26_io_out ? io_r_133_b : _GEN_19722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19724 = 10'h86 == r_count_26_io_out ? io_r_134_b : _GEN_19723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19725 = 10'h87 == r_count_26_io_out ? io_r_135_b : _GEN_19724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19726 = 10'h88 == r_count_26_io_out ? io_r_136_b : _GEN_19725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19727 = 10'h89 == r_count_26_io_out ? io_r_137_b : _GEN_19726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19728 = 10'h8a == r_count_26_io_out ? io_r_138_b : _GEN_19727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19729 = 10'h8b == r_count_26_io_out ? io_r_139_b : _GEN_19728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19730 = 10'h8c == r_count_26_io_out ? io_r_140_b : _GEN_19729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19731 = 10'h8d == r_count_26_io_out ? io_r_141_b : _GEN_19730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19732 = 10'h8e == r_count_26_io_out ? io_r_142_b : _GEN_19731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19733 = 10'h8f == r_count_26_io_out ? io_r_143_b : _GEN_19732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19734 = 10'h90 == r_count_26_io_out ? io_r_144_b : _GEN_19733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19735 = 10'h91 == r_count_26_io_out ? io_r_145_b : _GEN_19734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19736 = 10'h92 == r_count_26_io_out ? io_r_146_b : _GEN_19735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19737 = 10'h93 == r_count_26_io_out ? io_r_147_b : _GEN_19736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19738 = 10'h94 == r_count_26_io_out ? io_r_148_b : _GEN_19737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19739 = 10'h95 == r_count_26_io_out ? io_r_149_b : _GEN_19738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19740 = 10'h96 == r_count_26_io_out ? io_r_150_b : _GEN_19739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19741 = 10'h97 == r_count_26_io_out ? io_r_151_b : _GEN_19740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19742 = 10'h98 == r_count_26_io_out ? io_r_152_b : _GEN_19741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19743 = 10'h99 == r_count_26_io_out ? io_r_153_b : _GEN_19742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19744 = 10'h9a == r_count_26_io_out ? io_r_154_b : _GEN_19743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19745 = 10'h9b == r_count_26_io_out ? io_r_155_b : _GEN_19744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19746 = 10'h9c == r_count_26_io_out ? io_r_156_b : _GEN_19745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19747 = 10'h9d == r_count_26_io_out ? io_r_157_b : _GEN_19746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19748 = 10'h9e == r_count_26_io_out ? io_r_158_b : _GEN_19747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19749 = 10'h9f == r_count_26_io_out ? io_r_159_b : _GEN_19748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19750 = 10'ha0 == r_count_26_io_out ? io_r_160_b : _GEN_19749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19751 = 10'ha1 == r_count_26_io_out ? io_r_161_b : _GEN_19750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19752 = 10'ha2 == r_count_26_io_out ? io_r_162_b : _GEN_19751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19753 = 10'ha3 == r_count_26_io_out ? io_r_163_b : _GEN_19752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19754 = 10'ha4 == r_count_26_io_out ? io_r_164_b : _GEN_19753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19755 = 10'ha5 == r_count_26_io_out ? io_r_165_b : _GEN_19754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19756 = 10'ha6 == r_count_26_io_out ? io_r_166_b : _GEN_19755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19757 = 10'ha7 == r_count_26_io_out ? io_r_167_b : _GEN_19756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19758 = 10'ha8 == r_count_26_io_out ? io_r_168_b : _GEN_19757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19759 = 10'ha9 == r_count_26_io_out ? io_r_169_b : _GEN_19758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19760 = 10'haa == r_count_26_io_out ? io_r_170_b : _GEN_19759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19761 = 10'hab == r_count_26_io_out ? io_r_171_b : _GEN_19760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19762 = 10'hac == r_count_26_io_out ? io_r_172_b : _GEN_19761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19763 = 10'had == r_count_26_io_out ? io_r_173_b : _GEN_19762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19764 = 10'hae == r_count_26_io_out ? io_r_174_b : _GEN_19763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19765 = 10'haf == r_count_26_io_out ? io_r_175_b : _GEN_19764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19766 = 10'hb0 == r_count_26_io_out ? io_r_176_b : _GEN_19765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19767 = 10'hb1 == r_count_26_io_out ? io_r_177_b : _GEN_19766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19768 = 10'hb2 == r_count_26_io_out ? io_r_178_b : _GEN_19767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19769 = 10'hb3 == r_count_26_io_out ? io_r_179_b : _GEN_19768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19770 = 10'hb4 == r_count_26_io_out ? io_r_180_b : _GEN_19769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19771 = 10'hb5 == r_count_26_io_out ? io_r_181_b : _GEN_19770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19772 = 10'hb6 == r_count_26_io_out ? io_r_182_b : _GEN_19771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19773 = 10'hb7 == r_count_26_io_out ? io_r_183_b : _GEN_19772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19774 = 10'hb8 == r_count_26_io_out ? io_r_184_b : _GEN_19773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19775 = 10'hb9 == r_count_26_io_out ? io_r_185_b : _GEN_19774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19776 = 10'hba == r_count_26_io_out ? io_r_186_b : _GEN_19775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19777 = 10'hbb == r_count_26_io_out ? io_r_187_b : _GEN_19776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19778 = 10'hbc == r_count_26_io_out ? io_r_188_b : _GEN_19777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19779 = 10'hbd == r_count_26_io_out ? io_r_189_b : _GEN_19778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19780 = 10'hbe == r_count_26_io_out ? io_r_190_b : _GEN_19779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19781 = 10'hbf == r_count_26_io_out ? io_r_191_b : _GEN_19780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19782 = 10'hc0 == r_count_26_io_out ? io_r_192_b : _GEN_19781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19783 = 10'hc1 == r_count_26_io_out ? io_r_193_b : _GEN_19782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19784 = 10'hc2 == r_count_26_io_out ? io_r_194_b : _GEN_19783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19785 = 10'hc3 == r_count_26_io_out ? io_r_195_b : _GEN_19784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19786 = 10'hc4 == r_count_26_io_out ? io_r_196_b : _GEN_19785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19787 = 10'hc5 == r_count_26_io_out ? io_r_197_b : _GEN_19786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19788 = 10'hc6 == r_count_26_io_out ? io_r_198_b : _GEN_19787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19789 = 10'hc7 == r_count_26_io_out ? io_r_199_b : _GEN_19788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19790 = 10'hc8 == r_count_26_io_out ? io_r_200_b : _GEN_19789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19791 = 10'hc9 == r_count_26_io_out ? io_r_201_b : _GEN_19790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19792 = 10'hca == r_count_26_io_out ? io_r_202_b : _GEN_19791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19793 = 10'hcb == r_count_26_io_out ? io_r_203_b : _GEN_19792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19794 = 10'hcc == r_count_26_io_out ? io_r_204_b : _GEN_19793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19795 = 10'hcd == r_count_26_io_out ? io_r_205_b : _GEN_19794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19796 = 10'hce == r_count_26_io_out ? io_r_206_b : _GEN_19795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19797 = 10'hcf == r_count_26_io_out ? io_r_207_b : _GEN_19796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19798 = 10'hd0 == r_count_26_io_out ? io_r_208_b : _GEN_19797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19799 = 10'hd1 == r_count_26_io_out ? io_r_209_b : _GEN_19798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19800 = 10'hd2 == r_count_26_io_out ? io_r_210_b : _GEN_19799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19801 = 10'hd3 == r_count_26_io_out ? io_r_211_b : _GEN_19800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19802 = 10'hd4 == r_count_26_io_out ? io_r_212_b : _GEN_19801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19803 = 10'hd5 == r_count_26_io_out ? io_r_213_b : _GEN_19802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19804 = 10'hd6 == r_count_26_io_out ? io_r_214_b : _GEN_19803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19805 = 10'hd7 == r_count_26_io_out ? io_r_215_b : _GEN_19804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19806 = 10'hd8 == r_count_26_io_out ? io_r_216_b : _GEN_19805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19807 = 10'hd9 == r_count_26_io_out ? io_r_217_b : _GEN_19806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19808 = 10'hda == r_count_26_io_out ? io_r_218_b : _GEN_19807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19809 = 10'hdb == r_count_26_io_out ? io_r_219_b : _GEN_19808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19810 = 10'hdc == r_count_26_io_out ? io_r_220_b : _GEN_19809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19811 = 10'hdd == r_count_26_io_out ? io_r_221_b : _GEN_19810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19812 = 10'hde == r_count_26_io_out ? io_r_222_b : _GEN_19811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19813 = 10'hdf == r_count_26_io_out ? io_r_223_b : _GEN_19812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19814 = 10'he0 == r_count_26_io_out ? io_r_224_b : _GEN_19813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19815 = 10'he1 == r_count_26_io_out ? io_r_225_b : _GEN_19814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19816 = 10'he2 == r_count_26_io_out ? io_r_226_b : _GEN_19815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19817 = 10'he3 == r_count_26_io_out ? io_r_227_b : _GEN_19816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19818 = 10'he4 == r_count_26_io_out ? io_r_228_b : _GEN_19817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19819 = 10'he5 == r_count_26_io_out ? io_r_229_b : _GEN_19818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19820 = 10'he6 == r_count_26_io_out ? io_r_230_b : _GEN_19819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19821 = 10'he7 == r_count_26_io_out ? io_r_231_b : _GEN_19820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19822 = 10'he8 == r_count_26_io_out ? io_r_232_b : _GEN_19821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19823 = 10'he9 == r_count_26_io_out ? io_r_233_b : _GEN_19822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19824 = 10'hea == r_count_26_io_out ? io_r_234_b : _GEN_19823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19825 = 10'heb == r_count_26_io_out ? io_r_235_b : _GEN_19824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19826 = 10'hec == r_count_26_io_out ? io_r_236_b : _GEN_19825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19827 = 10'hed == r_count_26_io_out ? io_r_237_b : _GEN_19826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19828 = 10'hee == r_count_26_io_out ? io_r_238_b : _GEN_19827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19829 = 10'hef == r_count_26_io_out ? io_r_239_b : _GEN_19828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19830 = 10'hf0 == r_count_26_io_out ? io_r_240_b : _GEN_19829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19831 = 10'hf1 == r_count_26_io_out ? io_r_241_b : _GEN_19830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19832 = 10'hf2 == r_count_26_io_out ? io_r_242_b : _GEN_19831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19833 = 10'hf3 == r_count_26_io_out ? io_r_243_b : _GEN_19832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19834 = 10'hf4 == r_count_26_io_out ? io_r_244_b : _GEN_19833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19835 = 10'hf5 == r_count_26_io_out ? io_r_245_b : _GEN_19834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19836 = 10'hf6 == r_count_26_io_out ? io_r_246_b : _GEN_19835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19837 = 10'hf7 == r_count_26_io_out ? io_r_247_b : _GEN_19836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19838 = 10'hf8 == r_count_26_io_out ? io_r_248_b : _GEN_19837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19839 = 10'hf9 == r_count_26_io_out ? io_r_249_b : _GEN_19838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19840 = 10'hfa == r_count_26_io_out ? io_r_250_b : _GEN_19839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19841 = 10'hfb == r_count_26_io_out ? io_r_251_b : _GEN_19840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19842 = 10'hfc == r_count_26_io_out ? io_r_252_b : _GEN_19841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19843 = 10'hfd == r_count_26_io_out ? io_r_253_b : _GEN_19842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19844 = 10'hfe == r_count_26_io_out ? io_r_254_b : _GEN_19843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19845 = 10'hff == r_count_26_io_out ? io_r_255_b : _GEN_19844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19846 = 10'h100 == r_count_26_io_out ? io_r_256_b : _GEN_19845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19847 = 10'h101 == r_count_26_io_out ? io_r_257_b : _GEN_19846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19848 = 10'h102 == r_count_26_io_out ? io_r_258_b : _GEN_19847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19849 = 10'h103 == r_count_26_io_out ? io_r_259_b : _GEN_19848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19850 = 10'h104 == r_count_26_io_out ? io_r_260_b : _GEN_19849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19851 = 10'h105 == r_count_26_io_out ? io_r_261_b : _GEN_19850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19852 = 10'h106 == r_count_26_io_out ? io_r_262_b : _GEN_19851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19853 = 10'h107 == r_count_26_io_out ? io_r_263_b : _GEN_19852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19854 = 10'h108 == r_count_26_io_out ? io_r_264_b : _GEN_19853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19855 = 10'h109 == r_count_26_io_out ? io_r_265_b : _GEN_19854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19856 = 10'h10a == r_count_26_io_out ? io_r_266_b : _GEN_19855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19857 = 10'h10b == r_count_26_io_out ? io_r_267_b : _GEN_19856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19858 = 10'h10c == r_count_26_io_out ? io_r_268_b : _GEN_19857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19859 = 10'h10d == r_count_26_io_out ? io_r_269_b : _GEN_19858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19860 = 10'h10e == r_count_26_io_out ? io_r_270_b : _GEN_19859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19861 = 10'h10f == r_count_26_io_out ? io_r_271_b : _GEN_19860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19862 = 10'h110 == r_count_26_io_out ? io_r_272_b : _GEN_19861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19863 = 10'h111 == r_count_26_io_out ? io_r_273_b : _GEN_19862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19864 = 10'h112 == r_count_26_io_out ? io_r_274_b : _GEN_19863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19865 = 10'h113 == r_count_26_io_out ? io_r_275_b : _GEN_19864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19866 = 10'h114 == r_count_26_io_out ? io_r_276_b : _GEN_19865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19867 = 10'h115 == r_count_26_io_out ? io_r_277_b : _GEN_19866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19868 = 10'h116 == r_count_26_io_out ? io_r_278_b : _GEN_19867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19869 = 10'h117 == r_count_26_io_out ? io_r_279_b : _GEN_19868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19870 = 10'h118 == r_count_26_io_out ? io_r_280_b : _GEN_19869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19871 = 10'h119 == r_count_26_io_out ? io_r_281_b : _GEN_19870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19872 = 10'h11a == r_count_26_io_out ? io_r_282_b : _GEN_19871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19873 = 10'h11b == r_count_26_io_out ? io_r_283_b : _GEN_19872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19874 = 10'h11c == r_count_26_io_out ? io_r_284_b : _GEN_19873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19875 = 10'h11d == r_count_26_io_out ? io_r_285_b : _GEN_19874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19876 = 10'h11e == r_count_26_io_out ? io_r_286_b : _GEN_19875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19877 = 10'h11f == r_count_26_io_out ? io_r_287_b : _GEN_19876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19878 = 10'h120 == r_count_26_io_out ? io_r_288_b : _GEN_19877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19879 = 10'h121 == r_count_26_io_out ? io_r_289_b : _GEN_19878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19880 = 10'h122 == r_count_26_io_out ? io_r_290_b : _GEN_19879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19881 = 10'h123 == r_count_26_io_out ? io_r_291_b : _GEN_19880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19882 = 10'h124 == r_count_26_io_out ? io_r_292_b : _GEN_19881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19883 = 10'h125 == r_count_26_io_out ? io_r_293_b : _GEN_19882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19884 = 10'h126 == r_count_26_io_out ? io_r_294_b : _GEN_19883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19885 = 10'h127 == r_count_26_io_out ? io_r_295_b : _GEN_19884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19886 = 10'h128 == r_count_26_io_out ? io_r_296_b : _GEN_19885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19887 = 10'h129 == r_count_26_io_out ? io_r_297_b : _GEN_19886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19888 = 10'h12a == r_count_26_io_out ? io_r_298_b : _GEN_19887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19889 = 10'h12b == r_count_26_io_out ? io_r_299_b : _GEN_19888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19890 = 10'h12c == r_count_26_io_out ? io_r_300_b : _GEN_19889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19891 = 10'h12d == r_count_26_io_out ? io_r_301_b : _GEN_19890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19892 = 10'h12e == r_count_26_io_out ? io_r_302_b : _GEN_19891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19893 = 10'h12f == r_count_26_io_out ? io_r_303_b : _GEN_19892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19894 = 10'h130 == r_count_26_io_out ? io_r_304_b : _GEN_19893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19895 = 10'h131 == r_count_26_io_out ? io_r_305_b : _GEN_19894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19896 = 10'h132 == r_count_26_io_out ? io_r_306_b : _GEN_19895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19897 = 10'h133 == r_count_26_io_out ? io_r_307_b : _GEN_19896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19898 = 10'h134 == r_count_26_io_out ? io_r_308_b : _GEN_19897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19899 = 10'h135 == r_count_26_io_out ? io_r_309_b : _GEN_19898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19900 = 10'h136 == r_count_26_io_out ? io_r_310_b : _GEN_19899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19901 = 10'h137 == r_count_26_io_out ? io_r_311_b : _GEN_19900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19902 = 10'h138 == r_count_26_io_out ? io_r_312_b : _GEN_19901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19903 = 10'h139 == r_count_26_io_out ? io_r_313_b : _GEN_19902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19904 = 10'h13a == r_count_26_io_out ? io_r_314_b : _GEN_19903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19905 = 10'h13b == r_count_26_io_out ? io_r_315_b : _GEN_19904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19906 = 10'h13c == r_count_26_io_out ? io_r_316_b : _GEN_19905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19907 = 10'h13d == r_count_26_io_out ? io_r_317_b : _GEN_19906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19908 = 10'h13e == r_count_26_io_out ? io_r_318_b : _GEN_19907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19909 = 10'h13f == r_count_26_io_out ? io_r_319_b : _GEN_19908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19910 = 10'h140 == r_count_26_io_out ? io_r_320_b : _GEN_19909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19911 = 10'h141 == r_count_26_io_out ? io_r_321_b : _GEN_19910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19912 = 10'h142 == r_count_26_io_out ? io_r_322_b : _GEN_19911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19913 = 10'h143 == r_count_26_io_out ? io_r_323_b : _GEN_19912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19914 = 10'h144 == r_count_26_io_out ? io_r_324_b : _GEN_19913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19915 = 10'h145 == r_count_26_io_out ? io_r_325_b : _GEN_19914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19916 = 10'h146 == r_count_26_io_out ? io_r_326_b : _GEN_19915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19917 = 10'h147 == r_count_26_io_out ? io_r_327_b : _GEN_19916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19918 = 10'h148 == r_count_26_io_out ? io_r_328_b : _GEN_19917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19919 = 10'h149 == r_count_26_io_out ? io_r_329_b : _GEN_19918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19920 = 10'h14a == r_count_26_io_out ? io_r_330_b : _GEN_19919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19921 = 10'h14b == r_count_26_io_out ? io_r_331_b : _GEN_19920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19922 = 10'h14c == r_count_26_io_out ? io_r_332_b : _GEN_19921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19923 = 10'h14d == r_count_26_io_out ? io_r_333_b : _GEN_19922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19924 = 10'h14e == r_count_26_io_out ? io_r_334_b : _GEN_19923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19925 = 10'h14f == r_count_26_io_out ? io_r_335_b : _GEN_19924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19926 = 10'h150 == r_count_26_io_out ? io_r_336_b : _GEN_19925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19927 = 10'h151 == r_count_26_io_out ? io_r_337_b : _GEN_19926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19928 = 10'h152 == r_count_26_io_out ? io_r_338_b : _GEN_19927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19929 = 10'h153 == r_count_26_io_out ? io_r_339_b : _GEN_19928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19930 = 10'h154 == r_count_26_io_out ? io_r_340_b : _GEN_19929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19931 = 10'h155 == r_count_26_io_out ? io_r_341_b : _GEN_19930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19932 = 10'h156 == r_count_26_io_out ? io_r_342_b : _GEN_19931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19933 = 10'h157 == r_count_26_io_out ? io_r_343_b : _GEN_19932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19934 = 10'h158 == r_count_26_io_out ? io_r_344_b : _GEN_19933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19935 = 10'h159 == r_count_26_io_out ? io_r_345_b : _GEN_19934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19936 = 10'h15a == r_count_26_io_out ? io_r_346_b : _GEN_19935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19937 = 10'h15b == r_count_26_io_out ? io_r_347_b : _GEN_19936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19938 = 10'h15c == r_count_26_io_out ? io_r_348_b : _GEN_19937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19939 = 10'h15d == r_count_26_io_out ? io_r_349_b : _GEN_19938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19940 = 10'h15e == r_count_26_io_out ? io_r_350_b : _GEN_19939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19941 = 10'h15f == r_count_26_io_out ? io_r_351_b : _GEN_19940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19942 = 10'h160 == r_count_26_io_out ? io_r_352_b : _GEN_19941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19943 = 10'h161 == r_count_26_io_out ? io_r_353_b : _GEN_19942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19944 = 10'h162 == r_count_26_io_out ? io_r_354_b : _GEN_19943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19945 = 10'h163 == r_count_26_io_out ? io_r_355_b : _GEN_19944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19946 = 10'h164 == r_count_26_io_out ? io_r_356_b : _GEN_19945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19947 = 10'h165 == r_count_26_io_out ? io_r_357_b : _GEN_19946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19948 = 10'h166 == r_count_26_io_out ? io_r_358_b : _GEN_19947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19949 = 10'h167 == r_count_26_io_out ? io_r_359_b : _GEN_19948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19950 = 10'h168 == r_count_26_io_out ? io_r_360_b : _GEN_19949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19951 = 10'h169 == r_count_26_io_out ? io_r_361_b : _GEN_19950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19952 = 10'h16a == r_count_26_io_out ? io_r_362_b : _GEN_19951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19953 = 10'h16b == r_count_26_io_out ? io_r_363_b : _GEN_19952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19954 = 10'h16c == r_count_26_io_out ? io_r_364_b : _GEN_19953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19955 = 10'h16d == r_count_26_io_out ? io_r_365_b : _GEN_19954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19956 = 10'h16e == r_count_26_io_out ? io_r_366_b : _GEN_19955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19957 = 10'h16f == r_count_26_io_out ? io_r_367_b : _GEN_19956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19958 = 10'h170 == r_count_26_io_out ? io_r_368_b : _GEN_19957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19959 = 10'h171 == r_count_26_io_out ? io_r_369_b : _GEN_19958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19960 = 10'h172 == r_count_26_io_out ? io_r_370_b : _GEN_19959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19961 = 10'h173 == r_count_26_io_out ? io_r_371_b : _GEN_19960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19962 = 10'h174 == r_count_26_io_out ? io_r_372_b : _GEN_19961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19963 = 10'h175 == r_count_26_io_out ? io_r_373_b : _GEN_19962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19964 = 10'h176 == r_count_26_io_out ? io_r_374_b : _GEN_19963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19965 = 10'h177 == r_count_26_io_out ? io_r_375_b : _GEN_19964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19966 = 10'h178 == r_count_26_io_out ? io_r_376_b : _GEN_19965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19967 = 10'h179 == r_count_26_io_out ? io_r_377_b : _GEN_19966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19968 = 10'h17a == r_count_26_io_out ? io_r_378_b : _GEN_19967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19969 = 10'h17b == r_count_26_io_out ? io_r_379_b : _GEN_19968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19970 = 10'h17c == r_count_26_io_out ? io_r_380_b : _GEN_19969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19971 = 10'h17d == r_count_26_io_out ? io_r_381_b : _GEN_19970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19972 = 10'h17e == r_count_26_io_out ? io_r_382_b : _GEN_19971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19973 = 10'h17f == r_count_26_io_out ? io_r_383_b : _GEN_19972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19974 = 10'h180 == r_count_26_io_out ? io_r_384_b : _GEN_19973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19975 = 10'h181 == r_count_26_io_out ? io_r_385_b : _GEN_19974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19976 = 10'h182 == r_count_26_io_out ? io_r_386_b : _GEN_19975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19977 = 10'h183 == r_count_26_io_out ? io_r_387_b : _GEN_19976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19978 = 10'h184 == r_count_26_io_out ? io_r_388_b : _GEN_19977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19979 = 10'h185 == r_count_26_io_out ? io_r_389_b : _GEN_19978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19980 = 10'h186 == r_count_26_io_out ? io_r_390_b : _GEN_19979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19981 = 10'h187 == r_count_26_io_out ? io_r_391_b : _GEN_19980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19982 = 10'h188 == r_count_26_io_out ? io_r_392_b : _GEN_19981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19983 = 10'h189 == r_count_26_io_out ? io_r_393_b : _GEN_19982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19984 = 10'h18a == r_count_26_io_out ? io_r_394_b : _GEN_19983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19985 = 10'h18b == r_count_26_io_out ? io_r_395_b : _GEN_19984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19986 = 10'h18c == r_count_26_io_out ? io_r_396_b : _GEN_19985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19987 = 10'h18d == r_count_26_io_out ? io_r_397_b : _GEN_19986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19988 = 10'h18e == r_count_26_io_out ? io_r_398_b : _GEN_19987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19989 = 10'h18f == r_count_26_io_out ? io_r_399_b : _GEN_19988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19990 = 10'h190 == r_count_26_io_out ? io_r_400_b : _GEN_19989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19991 = 10'h191 == r_count_26_io_out ? io_r_401_b : _GEN_19990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19992 = 10'h192 == r_count_26_io_out ? io_r_402_b : _GEN_19991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19993 = 10'h193 == r_count_26_io_out ? io_r_403_b : _GEN_19992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19994 = 10'h194 == r_count_26_io_out ? io_r_404_b : _GEN_19993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19995 = 10'h195 == r_count_26_io_out ? io_r_405_b : _GEN_19994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19996 = 10'h196 == r_count_26_io_out ? io_r_406_b : _GEN_19995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19997 = 10'h197 == r_count_26_io_out ? io_r_407_b : _GEN_19996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19998 = 10'h198 == r_count_26_io_out ? io_r_408_b : _GEN_19997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19999 = 10'h199 == r_count_26_io_out ? io_r_409_b : _GEN_19998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20000 = 10'h19a == r_count_26_io_out ? io_r_410_b : _GEN_19999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20001 = 10'h19b == r_count_26_io_out ? io_r_411_b : _GEN_20000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20002 = 10'h19c == r_count_26_io_out ? io_r_412_b : _GEN_20001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20003 = 10'h19d == r_count_26_io_out ? io_r_413_b : _GEN_20002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20004 = 10'h19e == r_count_26_io_out ? io_r_414_b : _GEN_20003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20005 = 10'h19f == r_count_26_io_out ? io_r_415_b : _GEN_20004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20006 = 10'h1a0 == r_count_26_io_out ? io_r_416_b : _GEN_20005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20007 = 10'h1a1 == r_count_26_io_out ? io_r_417_b : _GEN_20006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20008 = 10'h1a2 == r_count_26_io_out ? io_r_418_b : _GEN_20007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20009 = 10'h1a3 == r_count_26_io_out ? io_r_419_b : _GEN_20008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20010 = 10'h1a4 == r_count_26_io_out ? io_r_420_b : _GEN_20009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20011 = 10'h1a5 == r_count_26_io_out ? io_r_421_b : _GEN_20010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20012 = 10'h1a6 == r_count_26_io_out ? io_r_422_b : _GEN_20011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20013 = 10'h1a7 == r_count_26_io_out ? io_r_423_b : _GEN_20012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20014 = 10'h1a8 == r_count_26_io_out ? io_r_424_b : _GEN_20013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20015 = 10'h1a9 == r_count_26_io_out ? io_r_425_b : _GEN_20014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20016 = 10'h1aa == r_count_26_io_out ? io_r_426_b : _GEN_20015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20017 = 10'h1ab == r_count_26_io_out ? io_r_427_b : _GEN_20016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20018 = 10'h1ac == r_count_26_io_out ? io_r_428_b : _GEN_20017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20019 = 10'h1ad == r_count_26_io_out ? io_r_429_b : _GEN_20018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20020 = 10'h1ae == r_count_26_io_out ? io_r_430_b : _GEN_20019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20021 = 10'h1af == r_count_26_io_out ? io_r_431_b : _GEN_20020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20022 = 10'h1b0 == r_count_26_io_out ? io_r_432_b : _GEN_20021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20023 = 10'h1b1 == r_count_26_io_out ? io_r_433_b : _GEN_20022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20024 = 10'h1b2 == r_count_26_io_out ? io_r_434_b : _GEN_20023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20025 = 10'h1b3 == r_count_26_io_out ? io_r_435_b : _GEN_20024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20026 = 10'h1b4 == r_count_26_io_out ? io_r_436_b : _GEN_20025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20027 = 10'h1b5 == r_count_26_io_out ? io_r_437_b : _GEN_20026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20028 = 10'h1b6 == r_count_26_io_out ? io_r_438_b : _GEN_20027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20029 = 10'h1b7 == r_count_26_io_out ? io_r_439_b : _GEN_20028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20030 = 10'h1b8 == r_count_26_io_out ? io_r_440_b : _GEN_20029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20031 = 10'h1b9 == r_count_26_io_out ? io_r_441_b : _GEN_20030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20032 = 10'h1ba == r_count_26_io_out ? io_r_442_b : _GEN_20031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20033 = 10'h1bb == r_count_26_io_out ? io_r_443_b : _GEN_20032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20034 = 10'h1bc == r_count_26_io_out ? io_r_444_b : _GEN_20033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20035 = 10'h1bd == r_count_26_io_out ? io_r_445_b : _GEN_20034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20036 = 10'h1be == r_count_26_io_out ? io_r_446_b : _GEN_20035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20037 = 10'h1bf == r_count_26_io_out ? io_r_447_b : _GEN_20036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20038 = 10'h1c0 == r_count_26_io_out ? io_r_448_b : _GEN_20037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20039 = 10'h1c1 == r_count_26_io_out ? io_r_449_b : _GEN_20038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20040 = 10'h1c2 == r_count_26_io_out ? io_r_450_b : _GEN_20039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20041 = 10'h1c3 == r_count_26_io_out ? io_r_451_b : _GEN_20040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20042 = 10'h1c4 == r_count_26_io_out ? io_r_452_b : _GEN_20041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20043 = 10'h1c5 == r_count_26_io_out ? io_r_453_b : _GEN_20042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20044 = 10'h1c6 == r_count_26_io_out ? io_r_454_b : _GEN_20043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20045 = 10'h1c7 == r_count_26_io_out ? io_r_455_b : _GEN_20044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20046 = 10'h1c8 == r_count_26_io_out ? io_r_456_b : _GEN_20045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20047 = 10'h1c9 == r_count_26_io_out ? io_r_457_b : _GEN_20046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20048 = 10'h1ca == r_count_26_io_out ? io_r_458_b : _GEN_20047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20049 = 10'h1cb == r_count_26_io_out ? io_r_459_b : _GEN_20048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20050 = 10'h1cc == r_count_26_io_out ? io_r_460_b : _GEN_20049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20051 = 10'h1cd == r_count_26_io_out ? io_r_461_b : _GEN_20050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20052 = 10'h1ce == r_count_26_io_out ? io_r_462_b : _GEN_20051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20053 = 10'h1cf == r_count_26_io_out ? io_r_463_b : _GEN_20052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20054 = 10'h1d0 == r_count_26_io_out ? io_r_464_b : _GEN_20053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20055 = 10'h1d1 == r_count_26_io_out ? io_r_465_b : _GEN_20054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20056 = 10'h1d2 == r_count_26_io_out ? io_r_466_b : _GEN_20055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20057 = 10'h1d3 == r_count_26_io_out ? io_r_467_b : _GEN_20056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20058 = 10'h1d4 == r_count_26_io_out ? io_r_468_b : _GEN_20057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20059 = 10'h1d5 == r_count_26_io_out ? io_r_469_b : _GEN_20058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20060 = 10'h1d6 == r_count_26_io_out ? io_r_470_b : _GEN_20059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20061 = 10'h1d7 == r_count_26_io_out ? io_r_471_b : _GEN_20060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20062 = 10'h1d8 == r_count_26_io_out ? io_r_472_b : _GEN_20061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20063 = 10'h1d9 == r_count_26_io_out ? io_r_473_b : _GEN_20062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20064 = 10'h1da == r_count_26_io_out ? io_r_474_b : _GEN_20063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20065 = 10'h1db == r_count_26_io_out ? io_r_475_b : _GEN_20064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20066 = 10'h1dc == r_count_26_io_out ? io_r_476_b : _GEN_20065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20067 = 10'h1dd == r_count_26_io_out ? io_r_477_b : _GEN_20066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20068 = 10'h1de == r_count_26_io_out ? io_r_478_b : _GEN_20067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20069 = 10'h1df == r_count_26_io_out ? io_r_479_b : _GEN_20068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20070 = 10'h1e0 == r_count_26_io_out ? io_r_480_b : _GEN_20069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20071 = 10'h1e1 == r_count_26_io_out ? io_r_481_b : _GEN_20070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20072 = 10'h1e2 == r_count_26_io_out ? io_r_482_b : _GEN_20071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20073 = 10'h1e3 == r_count_26_io_out ? io_r_483_b : _GEN_20072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20074 = 10'h1e4 == r_count_26_io_out ? io_r_484_b : _GEN_20073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20075 = 10'h1e5 == r_count_26_io_out ? io_r_485_b : _GEN_20074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20076 = 10'h1e6 == r_count_26_io_out ? io_r_486_b : _GEN_20075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20077 = 10'h1e7 == r_count_26_io_out ? io_r_487_b : _GEN_20076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20078 = 10'h1e8 == r_count_26_io_out ? io_r_488_b : _GEN_20077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20079 = 10'h1e9 == r_count_26_io_out ? io_r_489_b : _GEN_20078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20080 = 10'h1ea == r_count_26_io_out ? io_r_490_b : _GEN_20079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20081 = 10'h1eb == r_count_26_io_out ? io_r_491_b : _GEN_20080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20082 = 10'h1ec == r_count_26_io_out ? io_r_492_b : _GEN_20081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20083 = 10'h1ed == r_count_26_io_out ? io_r_493_b : _GEN_20082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20084 = 10'h1ee == r_count_26_io_out ? io_r_494_b : _GEN_20083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20085 = 10'h1ef == r_count_26_io_out ? io_r_495_b : _GEN_20084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20086 = 10'h1f0 == r_count_26_io_out ? io_r_496_b : _GEN_20085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20087 = 10'h1f1 == r_count_26_io_out ? io_r_497_b : _GEN_20086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20088 = 10'h1f2 == r_count_26_io_out ? io_r_498_b : _GEN_20087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20089 = 10'h1f3 == r_count_26_io_out ? io_r_499_b : _GEN_20088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20090 = 10'h1f4 == r_count_26_io_out ? io_r_500_b : _GEN_20089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20091 = 10'h1f5 == r_count_26_io_out ? io_r_501_b : _GEN_20090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20092 = 10'h1f6 == r_count_26_io_out ? io_r_502_b : _GEN_20091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20093 = 10'h1f7 == r_count_26_io_out ? io_r_503_b : _GEN_20092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20094 = 10'h1f8 == r_count_26_io_out ? io_r_504_b : _GEN_20093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20095 = 10'h1f9 == r_count_26_io_out ? io_r_505_b : _GEN_20094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20096 = 10'h1fa == r_count_26_io_out ? io_r_506_b : _GEN_20095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20097 = 10'h1fb == r_count_26_io_out ? io_r_507_b : _GEN_20096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20098 = 10'h1fc == r_count_26_io_out ? io_r_508_b : _GEN_20097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20099 = 10'h1fd == r_count_26_io_out ? io_r_509_b : _GEN_20098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20100 = 10'h1fe == r_count_26_io_out ? io_r_510_b : _GEN_20099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20101 = 10'h1ff == r_count_26_io_out ? io_r_511_b : _GEN_20100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20102 = 10'h200 == r_count_26_io_out ? io_r_512_b : _GEN_20101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20103 = 10'h201 == r_count_26_io_out ? io_r_513_b : _GEN_20102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20104 = 10'h202 == r_count_26_io_out ? io_r_514_b : _GEN_20103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20105 = 10'h203 == r_count_26_io_out ? io_r_515_b : _GEN_20104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20106 = 10'h204 == r_count_26_io_out ? io_r_516_b : _GEN_20105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20107 = 10'h205 == r_count_26_io_out ? io_r_517_b : _GEN_20106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20108 = 10'h206 == r_count_26_io_out ? io_r_518_b : _GEN_20107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20109 = 10'h207 == r_count_26_io_out ? io_r_519_b : _GEN_20108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20110 = 10'h208 == r_count_26_io_out ? io_r_520_b : _GEN_20109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20111 = 10'h209 == r_count_26_io_out ? io_r_521_b : _GEN_20110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20112 = 10'h20a == r_count_26_io_out ? io_r_522_b : _GEN_20111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20113 = 10'h20b == r_count_26_io_out ? io_r_523_b : _GEN_20112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20114 = 10'h20c == r_count_26_io_out ? io_r_524_b : _GEN_20113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20115 = 10'h20d == r_count_26_io_out ? io_r_525_b : _GEN_20114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20116 = 10'h20e == r_count_26_io_out ? io_r_526_b : _GEN_20115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20117 = 10'h20f == r_count_26_io_out ? io_r_527_b : _GEN_20116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20118 = 10'h210 == r_count_26_io_out ? io_r_528_b : _GEN_20117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20119 = 10'h211 == r_count_26_io_out ? io_r_529_b : _GEN_20118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20120 = 10'h212 == r_count_26_io_out ? io_r_530_b : _GEN_20119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20121 = 10'h213 == r_count_26_io_out ? io_r_531_b : _GEN_20120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20122 = 10'h214 == r_count_26_io_out ? io_r_532_b : _GEN_20121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20123 = 10'h215 == r_count_26_io_out ? io_r_533_b : _GEN_20122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20124 = 10'h216 == r_count_26_io_out ? io_r_534_b : _GEN_20123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20125 = 10'h217 == r_count_26_io_out ? io_r_535_b : _GEN_20124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20126 = 10'h218 == r_count_26_io_out ? io_r_536_b : _GEN_20125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20127 = 10'h219 == r_count_26_io_out ? io_r_537_b : _GEN_20126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20128 = 10'h21a == r_count_26_io_out ? io_r_538_b : _GEN_20127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20129 = 10'h21b == r_count_26_io_out ? io_r_539_b : _GEN_20128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20130 = 10'h21c == r_count_26_io_out ? io_r_540_b : _GEN_20129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20131 = 10'h21d == r_count_26_io_out ? io_r_541_b : _GEN_20130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20132 = 10'h21e == r_count_26_io_out ? io_r_542_b : _GEN_20131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20133 = 10'h21f == r_count_26_io_out ? io_r_543_b : _GEN_20132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20134 = 10'h220 == r_count_26_io_out ? io_r_544_b : _GEN_20133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20135 = 10'h221 == r_count_26_io_out ? io_r_545_b : _GEN_20134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20136 = 10'h222 == r_count_26_io_out ? io_r_546_b : _GEN_20135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20137 = 10'h223 == r_count_26_io_out ? io_r_547_b : _GEN_20136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20138 = 10'h224 == r_count_26_io_out ? io_r_548_b : _GEN_20137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20139 = 10'h225 == r_count_26_io_out ? io_r_549_b : _GEN_20138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20140 = 10'h226 == r_count_26_io_out ? io_r_550_b : _GEN_20139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20141 = 10'h227 == r_count_26_io_out ? io_r_551_b : _GEN_20140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20142 = 10'h228 == r_count_26_io_out ? io_r_552_b : _GEN_20141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20143 = 10'h229 == r_count_26_io_out ? io_r_553_b : _GEN_20142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20144 = 10'h22a == r_count_26_io_out ? io_r_554_b : _GEN_20143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20145 = 10'h22b == r_count_26_io_out ? io_r_555_b : _GEN_20144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20146 = 10'h22c == r_count_26_io_out ? io_r_556_b : _GEN_20145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20147 = 10'h22d == r_count_26_io_out ? io_r_557_b : _GEN_20146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20148 = 10'h22e == r_count_26_io_out ? io_r_558_b : _GEN_20147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20149 = 10'h22f == r_count_26_io_out ? io_r_559_b : _GEN_20148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20150 = 10'h230 == r_count_26_io_out ? io_r_560_b : _GEN_20149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20151 = 10'h231 == r_count_26_io_out ? io_r_561_b : _GEN_20150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20152 = 10'h232 == r_count_26_io_out ? io_r_562_b : _GEN_20151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20153 = 10'h233 == r_count_26_io_out ? io_r_563_b : _GEN_20152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20154 = 10'h234 == r_count_26_io_out ? io_r_564_b : _GEN_20153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20155 = 10'h235 == r_count_26_io_out ? io_r_565_b : _GEN_20154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20156 = 10'h236 == r_count_26_io_out ? io_r_566_b : _GEN_20155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20157 = 10'h237 == r_count_26_io_out ? io_r_567_b : _GEN_20156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20158 = 10'h238 == r_count_26_io_out ? io_r_568_b : _GEN_20157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20159 = 10'h239 == r_count_26_io_out ? io_r_569_b : _GEN_20158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20160 = 10'h23a == r_count_26_io_out ? io_r_570_b : _GEN_20159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20161 = 10'h23b == r_count_26_io_out ? io_r_571_b : _GEN_20160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20162 = 10'h23c == r_count_26_io_out ? io_r_572_b : _GEN_20161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20163 = 10'h23d == r_count_26_io_out ? io_r_573_b : _GEN_20162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20164 = 10'h23e == r_count_26_io_out ? io_r_574_b : _GEN_20163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20165 = 10'h23f == r_count_26_io_out ? io_r_575_b : _GEN_20164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20166 = 10'h240 == r_count_26_io_out ? io_r_576_b : _GEN_20165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20167 = 10'h241 == r_count_26_io_out ? io_r_577_b : _GEN_20166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20168 = 10'h242 == r_count_26_io_out ? io_r_578_b : _GEN_20167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20169 = 10'h243 == r_count_26_io_out ? io_r_579_b : _GEN_20168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20170 = 10'h244 == r_count_26_io_out ? io_r_580_b : _GEN_20169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20171 = 10'h245 == r_count_26_io_out ? io_r_581_b : _GEN_20170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20172 = 10'h246 == r_count_26_io_out ? io_r_582_b : _GEN_20171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20173 = 10'h247 == r_count_26_io_out ? io_r_583_b : _GEN_20172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20174 = 10'h248 == r_count_26_io_out ? io_r_584_b : _GEN_20173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20175 = 10'h249 == r_count_26_io_out ? io_r_585_b : _GEN_20174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20176 = 10'h24a == r_count_26_io_out ? io_r_586_b : _GEN_20175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20177 = 10'h24b == r_count_26_io_out ? io_r_587_b : _GEN_20176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20178 = 10'h24c == r_count_26_io_out ? io_r_588_b : _GEN_20177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20179 = 10'h24d == r_count_26_io_out ? io_r_589_b : _GEN_20178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20180 = 10'h24e == r_count_26_io_out ? io_r_590_b : _GEN_20179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20181 = 10'h24f == r_count_26_io_out ? io_r_591_b : _GEN_20180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20182 = 10'h250 == r_count_26_io_out ? io_r_592_b : _GEN_20181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20183 = 10'h251 == r_count_26_io_out ? io_r_593_b : _GEN_20182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20184 = 10'h252 == r_count_26_io_out ? io_r_594_b : _GEN_20183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20185 = 10'h253 == r_count_26_io_out ? io_r_595_b : _GEN_20184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20186 = 10'h254 == r_count_26_io_out ? io_r_596_b : _GEN_20185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20187 = 10'h255 == r_count_26_io_out ? io_r_597_b : _GEN_20186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20188 = 10'h256 == r_count_26_io_out ? io_r_598_b : _GEN_20187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20189 = 10'h257 == r_count_26_io_out ? io_r_599_b : _GEN_20188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20190 = 10'h258 == r_count_26_io_out ? io_r_600_b : _GEN_20189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20191 = 10'h259 == r_count_26_io_out ? io_r_601_b : _GEN_20190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20192 = 10'h25a == r_count_26_io_out ? io_r_602_b : _GEN_20191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20193 = 10'h25b == r_count_26_io_out ? io_r_603_b : _GEN_20192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20194 = 10'h25c == r_count_26_io_out ? io_r_604_b : _GEN_20193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20195 = 10'h25d == r_count_26_io_out ? io_r_605_b : _GEN_20194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20196 = 10'h25e == r_count_26_io_out ? io_r_606_b : _GEN_20195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20197 = 10'h25f == r_count_26_io_out ? io_r_607_b : _GEN_20196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20198 = 10'h260 == r_count_26_io_out ? io_r_608_b : _GEN_20197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20199 = 10'h261 == r_count_26_io_out ? io_r_609_b : _GEN_20198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20200 = 10'h262 == r_count_26_io_out ? io_r_610_b : _GEN_20199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20201 = 10'h263 == r_count_26_io_out ? io_r_611_b : _GEN_20200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20202 = 10'h264 == r_count_26_io_out ? io_r_612_b : _GEN_20201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20203 = 10'h265 == r_count_26_io_out ? io_r_613_b : _GEN_20202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20204 = 10'h266 == r_count_26_io_out ? io_r_614_b : _GEN_20203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20205 = 10'h267 == r_count_26_io_out ? io_r_615_b : _GEN_20204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20206 = 10'h268 == r_count_26_io_out ? io_r_616_b : _GEN_20205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20207 = 10'h269 == r_count_26_io_out ? io_r_617_b : _GEN_20206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20208 = 10'h26a == r_count_26_io_out ? io_r_618_b : _GEN_20207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20209 = 10'h26b == r_count_26_io_out ? io_r_619_b : _GEN_20208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20210 = 10'h26c == r_count_26_io_out ? io_r_620_b : _GEN_20209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20211 = 10'h26d == r_count_26_io_out ? io_r_621_b : _GEN_20210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20212 = 10'h26e == r_count_26_io_out ? io_r_622_b : _GEN_20211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20213 = 10'h26f == r_count_26_io_out ? io_r_623_b : _GEN_20212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20214 = 10'h270 == r_count_26_io_out ? io_r_624_b : _GEN_20213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20215 = 10'h271 == r_count_26_io_out ? io_r_625_b : _GEN_20214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20216 = 10'h272 == r_count_26_io_out ? io_r_626_b : _GEN_20215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20217 = 10'h273 == r_count_26_io_out ? io_r_627_b : _GEN_20216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20218 = 10'h274 == r_count_26_io_out ? io_r_628_b : _GEN_20217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20219 = 10'h275 == r_count_26_io_out ? io_r_629_b : _GEN_20218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20220 = 10'h276 == r_count_26_io_out ? io_r_630_b : _GEN_20219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20221 = 10'h277 == r_count_26_io_out ? io_r_631_b : _GEN_20220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20222 = 10'h278 == r_count_26_io_out ? io_r_632_b : _GEN_20221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20223 = 10'h279 == r_count_26_io_out ? io_r_633_b : _GEN_20222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20224 = 10'h27a == r_count_26_io_out ? io_r_634_b : _GEN_20223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20225 = 10'h27b == r_count_26_io_out ? io_r_635_b : _GEN_20224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20226 = 10'h27c == r_count_26_io_out ? io_r_636_b : _GEN_20225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20227 = 10'h27d == r_count_26_io_out ? io_r_637_b : _GEN_20226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20228 = 10'h27e == r_count_26_io_out ? io_r_638_b : _GEN_20227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20229 = 10'h27f == r_count_26_io_out ? io_r_639_b : _GEN_20228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20230 = 10'h280 == r_count_26_io_out ? io_r_640_b : _GEN_20229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20231 = 10'h281 == r_count_26_io_out ? io_r_641_b : _GEN_20230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20232 = 10'h282 == r_count_26_io_out ? io_r_642_b : _GEN_20231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20233 = 10'h283 == r_count_26_io_out ? io_r_643_b : _GEN_20232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20234 = 10'h284 == r_count_26_io_out ? io_r_644_b : _GEN_20233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20235 = 10'h285 == r_count_26_io_out ? io_r_645_b : _GEN_20234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20236 = 10'h286 == r_count_26_io_out ? io_r_646_b : _GEN_20235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20237 = 10'h287 == r_count_26_io_out ? io_r_647_b : _GEN_20236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20238 = 10'h288 == r_count_26_io_out ? io_r_648_b : _GEN_20237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20239 = 10'h289 == r_count_26_io_out ? io_r_649_b : _GEN_20238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20240 = 10'h28a == r_count_26_io_out ? io_r_650_b : _GEN_20239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20241 = 10'h28b == r_count_26_io_out ? io_r_651_b : _GEN_20240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20242 = 10'h28c == r_count_26_io_out ? io_r_652_b : _GEN_20241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20243 = 10'h28d == r_count_26_io_out ? io_r_653_b : _GEN_20242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20244 = 10'h28e == r_count_26_io_out ? io_r_654_b : _GEN_20243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20245 = 10'h28f == r_count_26_io_out ? io_r_655_b : _GEN_20244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20246 = 10'h290 == r_count_26_io_out ? io_r_656_b : _GEN_20245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20247 = 10'h291 == r_count_26_io_out ? io_r_657_b : _GEN_20246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20248 = 10'h292 == r_count_26_io_out ? io_r_658_b : _GEN_20247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20249 = 10'h293 == r_count_26_io_out ? io_r_659_b : _GEN_20248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20250 = 10'h294 == r_count_26_io_out ? io_r_660_b : _GEN_20249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20251 = 10'h295 == r_count_26_io_out ? io_r_661_b : _GEN_20250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20252 = 10'h296 == r_count_26_io_out ? io_r_662_b : _GEN_20251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20253 = 10'h297 == r_count_26_io_out ? io_r_663_b : _GEN_20252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20254 = 10'h298 == r_count_26_io_out ? io_r_664_b : _GEN_20253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20255 = 10'h299 == r_count_26_io_out ? io_r_665_b : _GEN_20254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20256 = 10'h29a == r_count_26_io_out ? io_r_666_b : _GEN_20255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20257 = 10'h29b == r_count_26_io_out ? io_r_667_b : _GEN_20256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20258 = 10'h29c == r_count_26_io_out ? io_r_668_b : _GEN_20257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20259 = 10'h29d == r_count_26_io_out ? io_r_669_b : _GEN_20258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20260 = 10'h29e == r_count_26_io_out ? io_r_670_b : _GEN_20259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20261 = 10'h29f == r_count_26_io_out ? io_r_671_b : _GEN_20260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20262 = 10'h2a0 == r_count_26_io_out ? io_r_672_b : _GEN_20261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20263 = 10'h2a1 == r_count_26_io_out ? io_r_673_b : _GEN_20262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20264 = 10'h2a2 == r_count_26_io_out ? io_r_674_b : _GEN_20263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20265 = 10'h2a3 == r_count_26_io_out ? io_r_675_b : _GEN_20264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20266 = 10'h2a4 == r_count_26_io_out ? io_r_676_b : _GEN_20265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20267 = 10'h2a5 == r_count_26_io_out ? io_r_677_b : _GEN_20266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20268 = 10'h2a6 == r_count_26_io_out ? io_r_678_b : _GEN_20267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20269 = 10'h2a7 == r_count_26_io_out ? io_r_679_b : _GEN_20268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20270 = 10'h2a8 == r_count_26_io_out ? io_r_680_b : _GEN_20269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20271 = 10'h2a9 == r_count_26_io_out ? io_r_681_b : _GEN_20270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20272 = 10'h2aa == r_count_26_io_out ? io_r_682_b : _GEN_20271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20273 = 10'h2ab == r_count_26_io_out ? io_r_683_b : _GEN_20272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20274 = 10'h2ac == r_count_26_io_out ? io_r_684_b : _GEN_20273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20275 = 10'h2ad == r_count_26_io_out ? io_r_685_b : _GEN_20274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20276 = 10'h2ae == r_count_26_io_out ? io_r_686_b : _GEN_20275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20277 = 10'h2af == r_count_26_io_out ? io_r_687_b : _GEN_20276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20278 = 10'h2b0 == r_count_26_io_out ? io_r_688_b : _GEN_20277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20279 = 10'h2b1 == r_count_26_io_out ? io_r_689_b : _GEN_20278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20280 = 10'h2b2 == r_count_26_io_out ? io_r_690_b : _GEN_20279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20281 = 10'h2b3 == r_count_26_io_out ? io_r_691_b : _GEN_20280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20282 = 10'h2b4 == r_count_26_io_out ? io_r_692_b : _GEN_20281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20283 = 10'h2b5 == r_count_26_io_out ? io_r_693_b : _GEN_20282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20284 = 10'h2b6 == r_count_26_io_out ? io_r_694_b : _GEN_20283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20285 = 10'h2b7 == r_count_26_io_out ? io_r_695_b : _GEN_20284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20286 = 10'h2b8 == r_count_26_io_out ? io_r_696_b : _GEN_20285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20287 = 10'h2b9 == r_count_26_io_out ? io_r_697_b : _GEN_20286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20288 = 10'h2ba == r_count_26_io_out ? io_r_698_b : _GEN_20287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20289 = 10'h2bb == r_count_26_io_out ? io_r_699_b : _GEN_20288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20290 = 10'h2bc == r_count_26_io_out ? io_r_700_b : _GEN_20289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20291 = 10'h2bd == r_count_26_io_out ? io_r_701_b : _GEN_20290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20292 = 10'h2be == r_count_26_io_out ? io_r_702_b : _GEN_20291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20293 = 10'h2bf == r_count_26_io_out ? io_r_703_b : _GEN_20292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20294 = 10'h2c0 == r_count_26_io_out ? io_r_704_b : _GEN_20293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20295 = 10'h2c1 == r_count_26_io_out ? io_r_705_b : _GEN_20294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20296 = 10'h2c2 == r_count_26_io_out ? io_r_706_b : _GEN_20295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20297 = 10'h2c3 == r_count_26_io_out ? io_r_707_b : _GEN_20296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20298 = 10'h2c4 == r_count_26_io_out ? io_r_708_b : _GEN_20297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20299 = 10'h2c5 == r_count_26_io_out ? io_r_709_b : _GEN_20298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20300 = 10'h2c6 == r_count_26_io_out ? io_r_710_b : _GEN_20299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20301 = 10'h2c7 == r_count_26_io_out ? io_r_711_b : _GEN_20300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20302 = 10'h2c8 == r_count_26_io_out ? io_r_712_b : _GEN_20301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20303 = 10'h2c9 == r_count_26_io_out ? io_r_713_b : _GEN_20302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20304 = 10'h2ca == r_count_26_io_out ? io_r_714_b : _GEN_20303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20305 = 10'h2cb == r_count_26_io_out ? io_r_715_b : _GEN_20304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20306 = 10'h2cc == r_count_26_io_out ? io_r_716_b : _GEN_20305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20307 = 10'h2cd == r_count_26_io_out ? io_r_717_b : _GEN_20306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20308 = 10'h2ce == r_count_26_io_out ? io_r_718_b : _GEN_20307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20309 = 10'h2cf == r_count_26_io_out ? io_r_719_b : _GEN_20308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20310 = 10'h2d0 == r_count_26_io_out ? io_r_720_b : _GEN_20309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20311 = 10'h2d1 == r_count_26_io_out ? io_r_721_b : _GEN_20310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20312 = 10'h2d2 == r_count_26_io_out ? io_r_722_b : _GEN_20311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20313 = 10'h2d3 == r_count_26_io_out ? io_r_723_b : _GEN_20312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20314 = 10'h2d4 == r_count_26_io_out ? io_r_724_b : _GEN_20313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20315 = 10'h2d5 == r_count_26_io_out ? io_r_725_b : _GEN_20314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20316 = 10'h2d6 == r_count_26_io_out ? io_r_726_b : _GEN_20315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20317 = 10'h2d7 == r_count_26_io_out ? io_r_727_b : _GEN_20316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20318 = 10'h2d8 == r_count_26_io_out ? io_r_728_b : _GEN_20317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20319 = 10'h2d9 == r_count_26_io_out ? io_r_729_b : _GEN_20318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20320 = 10'h2da == r_count_26_io_out ? io_r_730_b : _GEN_20319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20321 = 10'h2db == r_count_26_io_out ? io_r_731_b : _GEN_20320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20322 = 10'h2dc == r_count_26_io_out ? io_r_732_b : _GEN_20321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20323 = 10'h2dd == r_count_26_io_out ? io_r_733_b : _GEN_20322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20324 = 10'h2de == r_count_26_io_out ? io_r_734_b : _GEN_20323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20325 = 10'h2df == r_count_26_io_out ? io_r_735_b : _GEN_20324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20326 = 10'h2e0 == r_count_26_io_out ? io_r_736_b : _GEN_20325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20327 = 10'h2e1 == r_count_26_io_out ? io_r_737_b : _GEN_20326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20328 = 10'h2e2 == r_count_26_io_out ? io_r_738_b : _GEN_20327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20329 = 10'h2e3 == r_count_26_io_out ? io_r_739_b : _GEN_20328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20330 = 10'h2e4 == r_count_26_io_out ? io_r_740_b : _GEN_20329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20331 = 10'h2e5 == r_count_26_io_out ? io_r_741_b : _GEN_20330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20332 = 10'h2e6 == r_count_26_io_out ? io_r_742_b : _GEN_20331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20333 = 10'h2e7 == r_count_26_io_out ? io_r_743_b : _GEN_20332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20334 = 10'h2e8 == r_count_26_io_out ? io_r_744_b : _GEN_20333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20335 = 10'h2e9 == r_count_26_io_out ? io_r_745_b : _GEN_20334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20336 = 10'h2ea == r_count_26_io_out ? io_r_746_b : _GEN_20335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20337 = 10'h2eb == r_count_26_io_out ? io_r_747_b : _GEN_20336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20338 = 10'h2ec == r_count_26_io_out ? io_r_748_b : _GEN_20337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20341 = 10'h1 == r_count_27_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20342 = 10'h2 == r_count_27_io_out ? io_r_2_b : _GEN_20341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20343 = 10'h3 == r_count_27_io_out ? io_r_3_b : _GEN_20342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20344 = 10'h4 == r_count_27_io_out ? io_r_4_b : _GEN_20343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20345 = 10'h5 == r_count_27_io_out ? io_r_5_b : _GEN_20344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20346 = 10'h6 == r_count_27_io_out ? io_r_6_b : _GEN_20345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20347 = 10'h7 == r_count_27_io_out ? io_r_7_b : _GEN_20346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20348 = 10'h8 == r_count_27_io_out ? io_r_8_b : _GEN_20347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20349 = 10'h9 == r_count_27_io_out ? io_r_9_b : _GEN_20348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20350 = 10'ha == r_count_27_io_out ? io_r_10_b : _GEN_20349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20351 = 10'hb == r_count_27_io_out ? io_r_11_b : _GEN_20350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20352 = 10'hc == r_count_27_io_out ? io_r_12_b : _GEN_20351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20353 = 10'hd == r_count_27_io_out ? io_r_13_b : _GEN_20352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20354 = 10'he == r_count_27_io_out ? io_r_14_b : _GEN_20353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20355 = 10'hf == r_count_27_io_out ? io_r_15_b : _GEN_20354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20356 = 10'h10 == r_count_27_io_out ? io_r_16_b : _GEN_20355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20357 = 10'h11 == r_count_27_io_out ? io_r_17_b : _GEN_20356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20358 = 10'h12 == r_count_27_io_out ? io_r_18_b : _GEN_20357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20359 = 10'h13 == r_count_27_io_out ? io_r_19_b : _GEN_20358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20360 = 10'h14 == r_count_27_io_out ? io_r_20_b : _GEN_20359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20361 = 10'h15 == r_count_27_io_out ? io_r_21_b : _GEN_20360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20362 = 10'h16 == r_count_27_io_out ? io_r_22_b : _GEN_20361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20363 = 10'h17 == r_count_27_io_out ? io_r_23_b : _GEN_20362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20364 = 10'h18 == r_count_27_io_out ? io_r_24_b : _GEN_20363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20365 = 10'h19 == r_count_27_io_out ? io_r_25_b : _GEN_20364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20366 = 10'h1a == r_count_27_io_out ? io_r_26_b : _GEN_20365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20367 = 10'h1b == r_count_27_io_out ? io_r_27_b : _GEN_20366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20368 = 10'h1c == r_count_27_io_out ? io_r_28_b : _GEN_20367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20369 = 10'h1d == r_count_27_io_out ? io_r_29_b : _GEN_20368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20370 = 10'h1e == r_count_27_io_out ? io_r_30_b : _GEN_20369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20371 = 10'h1f == r_count_27_io_out ? io_r_31_b : _GEN_20370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20372 = 10'h20 == r_count_27_io_out ? io_r_32_b : _GEN_20371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20373 = 10'h21 == r_count_27_io_out ? io_r_33_b : _GEN_20372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20374 = 10'h22 == r_count_27_io_out ? io_r_34_b : _GEN_20373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20375 = 10'h23 == r_count_27_io_out ? io_r_35_b : _GEN_20374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20376 = 10'h24 == r_count_27_io_out ? io_r_36_b : _GEN_20375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20377 = 10'h25 == r_count_27_io_out ? io_r_37_b : _GEN_20376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20378 = 10'h26 == r_count_27_io_out ? io_r_38_b : _GEN_20377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20379 = 10'h27 == r_count_27_io_out ? io_r_39_b : _GEN_20378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20380 = 10'h28 == r_count_27_io_out ? io_r_40_b : _GEN_20379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20381 = 10'h29 == r_count_27_io_out ? io_r_41_b : _GEN_20380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20382 = 10'h2a == r_count_27_io_out ? io_r_42_b : _GEN_20381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20383 = 10'h2b == r_count_27_io_out ? io_r_43_b : _GEN_20382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20384 = 10'h2c == r_count_27_io_out ? io_r_44_b : _GEN_20383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20385 = 10'h2d == r_count_27_io_out ? io_r_45_b : _GEN_20384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20386 = 10'h2e == r_count_27_io_out ? io_r_46_b : _GEN_20385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20387 = 10'h2f == r_count_27_io_out ? io_r_47_b : _GEN_20386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20388 = 10'h30 == r_count_27_io_out ? io_r_48_b : _GEN_20387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20389 = 10'h31 == r_count_27_io_out ? io_r_49_b : _GEN_20388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20390 = 10'h32 == r_count_27_io_out ? io_r_50_b : _GEN_20389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20391 = 10'h33 == r_count_27_io_out ? io_r_51_b : _GEN_20390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20392 = 10'h34 == r_count_27_io_out ? io_r_52_b : _GEN_20391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20393 = 10'h35 == r_count_27_io_out ? io_r_53_b : _GEN_20392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20394 = 10'h36 == r_count_27_io_out ? io_r_54_b : _GEN_20393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20395 = 10'h37 == r_count_27_io_out ? io_r_55_b : _GEN_20394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20396 = 10'h38 == r_count_27_io_out ? io_r_56_b : _GEN_20395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20397 = 10'h39 == r_count_27_io_out ? io_r_57_b : _GEN_20396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20398 = 10'h3a == r_count_27_io_out ? io_r_58_b : _GEN_20397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20399 = 10'h3b == r_count_27_io_out ? io_r_59_b : _GEN_20398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20400 = 10'h3c == r_count_27_io_out ? io_r_60_b : _GEN_20399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20401 = 10'h3d == r_count_27_io_out ? io_r_61_b : _GEN_20400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20402 = 10'h3e == r_count_27_io_out ? io_r_62_b : _GEN_20401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20403 = 10'h3f == r_count_27_io_out ? io_r_63_b : _GEN_20402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20404 = 10'h40 == r_count_27_io_out ? io_r_64_b : _GEN_20403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20405 = 10'h41 == r_count_27_io_out ? io_r_65_b : _GEN_20404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20406 = 10'h42 == r_count_27_io_out ? io_r_66_b : _GEN_20405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20407 = 10'h43 == r_count_27_io_out ? io_r_67_b : _GEN_20406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20408 = 10'h44 == r_count_27_io_out ? io_r_68_b : _GEN_20407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20409 = 10'h45 == r_count_27_io_out ? io_r_69_b : _GEN_20408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20410 = 10'h46 == r_count_27_io_out ? io_r_70_b : _GEN_20409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20411 = 10'h47 == r_count_27_io_out ? io_r_71_b : _GEN_20410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20412 = 10'h48 == r_count_27_io_out ? io_r_72_b : _GEN_20411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20413 = 10'h49 == r_count_27_io_out ? io_r_73_b : _GEN_20412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20414 = 10'h4a == r_count_27_io_out ? io_r_74_b : _GEN_20413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20415 = 10'h4b == r_count_27_io_out ? io_r_75_b : _GEN_20414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20416 = 10'h4c == r_count_27_io_out ? io_r_76_b : _GEN_20415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20417 = 10'h4d == r_count_27_io_out ? io_r_77_b : _GEN_20416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20418 = 10'h4e == r_count_27_io_out ? io_r_78_b : _GEN_20417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20419 = 10'h4f == r_count_27_io_out ? io_r_79_b : _GEN_20418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20420 = 10'h50 == r_count_27_io_out ? io_r_80_b : _GEN_20419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20421 = 10'h51 == r_count_27_io_out ? io_r_81_b : _GEN_20420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20422 = 10'h52 == r_count_27_io_out ? io_r_82_b : _GEN_20421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20423 = 10'h53 == r_count_27_io_out ? io_r_83_b : _GEN_20422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20424 = 10'h54 == r_count_27_io_out ? io_r_84_b : _GEN_20423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20425 = 10'h55 == r_count_27_io_out ? io_r_85_b : _GEN_20424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20426 = 10'h56 == r_count_27_io_out ? io_r_86_b : _GEN_20425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20427 = 10'h57 == r_count_27_io_out ? io_r_87_b : _GEN_20426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20428 = 10'h58 == r_count_27_io_out ? io_r_88_b : _GEN_20427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20429 = 10'h59 == r_count_27_io_out ? io_r_89_b : _GEN_20428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20430 = 10'h5a == r_count_27_io_out ? io_r_90_b : _GEN_20429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20431 = 10'h5b == r_count_27_io_out ? io_r_91_b : _GEN_20430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20432 = 10'h5c == r_count_27_io_out ? io_r_92_b : _GEN_20431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20433 = 10'h5d == r_count_27_io_out ? io_r_93_b : _GEN_20432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20434 = 10'h5e == r_count_27_io_out ? io_r_94_b : _GEN_20433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20435 = 10'h5f == r_count_27_io_out ? io_r_95_b : _GEN_20434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20436 = 10'h60 == r_count_27_io_out ? io_r_96_b : _GEN_20435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20437 = 10'h61 == r_count_27_io_out ? io_r_97_b : _GEN_20436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20438 = 10'h62 == r_count_27_io_out ? io_r_98_b : _GEN_20437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20439 = 10'h63 == r_count_27_io_out ? io_r_99_b : _GEN_20438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20440 = 10'h64 == r_count_27_io_out ? io_r_100_b : _GEN_20439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20441 = 10'h65 == r_count_27_io_out ? io_r_101_b : _GEN_20440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20442 = 10'h66 == r_count_27_io_out ? io_r_102_b : _GEN_20441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20443 = 10'h67 == r_count_27_io_out ? io_r_103_b : _GEN_20442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20444 = 10'h68 == r_count_27_io_out ? io_r_104_b : _GEN_20443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20445 = 10'h69 == r_count_27_io_out ? io_r_105_b : _GEN_20444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20446 = 10'h6a == r_count_27_io_out ? io_r_106_b : _GEN_20445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20447 = 10'h6b == r_count_27_io_out ? io_r_107_b : _GEN_20446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20448 = 10'h6c == r_count_27_io_out ? io_r_108_b : _GEN_20447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20449 = 10'h6d == r_count_27_io_out ? io_r_109_b : _GEN_20448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20450 = 10'h6e == r_count_27_io_out ? io_r_110_b : _GEN_20449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20451 = 10'h6f == r_count_27_io_out ? io_r_111_b : _GEN_20450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20452 = 10'h70 == r_count_27_io_out ? io_r_112_b : _GEN_20451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20453 = 10'h71 == r_count_27_io_out ? io_r_113_b : _GEN_20452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20454 = 10'h72 == r_count_27_io_out ? io_r_114_b : _GEN_20453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20455 = 10'h73 == r_count_27_io_out ? io_r_115_b : _GEN_20454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20456 = 10'h74 == r_count_27_io_out ? io_r_116_b : _GEN_20455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20457 = 10'h75 == r_count_27_io_out ? io_r_117_b : _GEN_20456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20458 = 10'h76 == r_count_27_io_out ? io_r_118_b : _GEN_20457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20459 = 10'h77 == r_count_27_io_out ? io_r_119_b : _GEN_20458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20460 = 10'h78 == r_count_27_io_out ? io_r_120_b : _GEN_20459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20461 = 10'h79 == r_count_27_io_out ? io_r_121_b : _GEN_20460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20462 = 10'h7a == r_count_27_io_out ? io_r_122_b : _GEN_20461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20463 = 10'h7b == r_count_27_io_out ? io_r_123_b : _GEN_20462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20464 = 10'h7c == r_count_27_io_out ? io_r_124_b : _GEN_20463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20465 = 10'h7d == r_count_27_io_out ? io_r_125_b : _GEN_20464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20466 = 10'h7e == r_count_27_io_out ? io_r_126_b : _GEN_20465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20467 = 10'h7f == r_count_27_io_out ? io_r_127_b : _GEN_20466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20468 = 10'h80 == r_count_27_io_out ? io_r_128_b : _GEN_20467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20469 = 10'h81 == r_count_27_io_out ? io_r_129_b : _GEN_20468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20470 = 10'h82 == r_count_27_io_out ? io_r_130_b : _GEN_20469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20471 = 10'h83 == r_count_27_io_out ? io_r_131_b : _GEN_20470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20472 = 10'h84 == r_count_27_io_out ? io_r_132_b : _GEN_20471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20473 = 10'h85 == r_count_27_io_out ? io_r_133_b : _GEN_20472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20474 = 10'h86 == r_count_27_io_out ? io_r_134_b : _GEN_20473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20475 = 10'h87 == r_count_27_io_out ? io_r_135_b : _GEN_20474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20476 = 10'h88 == r_count_27_io_out ? io_r_136_b : _GEN_20475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20477 = 10'h89 == r_count_27_io_out ? io_r_137_b : _GEN_20476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20478 = 10'h8a == r_count_27_io_out ? io_r_138_b : _GEN_20477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20479 = 10'h8b == r_count_27_io_out ? io_r_139_b : _GEN_20478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20480 = 10'h8c == r_count_27_io_out ? io_r_140_b : _GEN_20479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20481 = 10'h8d == r_count_27_io_out ? io_r_141_b : _GEN_20480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20482 = 10'h8e == r_count_27_io_out ? io_r_142_b : _GEN_20481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20483 = 10'h8f == r_count_27_io_out ? io_r_143_b : _GEN_20482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20484 = 10'h90 == r_count_27_io_out ? io_r_144_b : _GEN_20483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20485 = 10'h91 == r_count_27_io_out ? io_r_145_b : _GEN_20484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20486 = 10'h92 == r_count_27_io_out ? io_r_146_b : _GEN_20485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20487 = 10'h93 == r_count_27_io_out ? io_r_147_b : _GEN_20486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20488 = 10'h94 == r_count_27_io_out ? io_r_148_b : _GEN_20487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20489 = 10'h95 == r_count_27_io_out ? io_r_149_b : _GEN_20488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20490 = 10'h96 == r_count_27_io_out ? io_r_150_b : _GEN_20489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20491 = 10'h97 == r_count_27_io_out ? io_r_151_b : _GEN_20490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20492 = 10'h98 == r_count_27_io_out ? io_r_152_b : _GEN_20491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20493 = 10'h99 == r_count_27_io_out ? io_r_153_b : _GEN_20492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20494 = 10'h9a == r_count_27_io_out ? io_r_154_b : _GEN_20493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20495 = 10'h9b == r_count_27_io_out ? io_r_155_b : _GEN_20494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20496 = 10'h9c == r_count_27_io_out ? io_r_156_b : _GEN_20495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20497 = 10'h9d == r_count_27_io_out ? io_r_157_b : _GEN_20496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20498 = 10'h9e == r_count_27_io_out ? io_r_158_b : _GEN_20497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20499 = 10'h9f == r_count_27_io_out ? io_r_159_b : _GEN_20498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20500 = 10'ha0 == r_count_27_io_out ? io_r_160_b : _GEN_20499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20501 = 10'ha1 == r_count_27_io_out ? io_r_161_b : _GEN_20500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20502 = 10'ha2 == r_count_27_io_out ? io_r_162_b : _GEN_20501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20503 = 10'ha3 == r_count_27_io_out ? io_r_163_b : _GEN_20502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20504 = 10'ha4 == r_count_27_io_out ? io_r_164_b : _GEN_20503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20505 = 10'ha5 == r_count_27_io_out ? io_r_165_b : _GEN_20504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20506 = 10'ha6 == r_count_27_io_out ? io_r_166_b : _GEN_20505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20507 = 10'ha7 == r_count_27_io_out ? io_r_167_b : _GEN_20506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20508 = 10'ha8 == r_count_27_io_out ? io_r_168_b : _GEN_20507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20509 = 10'ha9 == r_count_27_io_out ? io_r_169_b : _GEN_20508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20510 = 10'haa == r_count_27_io_out ? io_r_170_b : _GEN_20509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20511 = 10'hab == r_count_27_io_out ? io_r_171_b : _GEN_20510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20512 = 10'hac == r_count_27_io_out ? io_r_172_b : _GEN_20511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20513 = 10'had == r_count_27_io_out ? io_r_173_b : _GEN_20512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20514 = 10'hae == r_count_27_io_out ? io_r_174_b : _GEN_20513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20515 = 10'haf == r_count_27_io_out ? io_r_175_b : _GEN_20514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20516 = 10'hb0 == r_count_27_io_out ? io_r_176_b : _GEN_20515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20517 = 10'hb1 == r_count_27_io_out ? io_r_177_b : _GEN_20516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20518 = 10'hb2 == r_count_27_io_out ? io_r_178_b : _GEN_20517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20519 = 10'hb3 == r_count_27_io_out ? io_r_179_b : _GEN_20518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20520 = 10'hb4 == r_count_27_io_out ? io_r_180_b : _GEN_20519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20521 = 10'hb5 == r_count_27_io_out ? io_r_181_b : _GEN_20520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20522 = 10'hb6 == r_count_27_io_out ? io_r_182_b : _GEN_20521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20523 = 10'hb7 == r_count_27_io_out ? io_r_183_b : _GEN_20522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20524 = 10'hb8 == r_count_27_io_out ? io_r_184_b : _GEN_20523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20525 = 10'hb9 == r_count_27_io_out ? io_r_185_b : _GEN_20524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20526 = 10'hba == r_count_27_io_out ? io_r_186_b : _GEN_20525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20527 = 10'hbb == r_count_27_io_out ? io_r_187_b : _GEN_20526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20528 = 10'hbc == r_count_27_io_out ? io_r_188_b : _GEN_20527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20529 = 10'hbd == r_count_27_io_out ? io_r_189_b : _GEN_20528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20530 = 10'hbe == r_count_27_io_out ? io_r_190_b : _GEN_20529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20531 = 10'hbf == r_count_27_io_out ? io_r_191_b : _GEN_20530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20532 = 10'hc0 == r_count_27_io_out ? io_r_192_b : _GEN_20531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20533 = 10'hc1 == r_count_27_io_out ? io_r_193_b : _GEN_20532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20534 = 10'hc2 == r_count_27_io_out ? io_r_194_b : _GEN_20533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20535 = 10'hc3 == r_count_27_io_out ? io_r_195_b : _GEN_20534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20536 = 10'hc4 == r_count_27_io_out ? io_r_196_b : _GEN_20535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20537 = 10'hc5 == r_count_27_io_out ? io_r_197_b : _GEN_20536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20538 = 10'hc6 == r_count_27_io_out ? io_r_198_b : _GEN_20537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20539 = 10'hc7 == r_count_27_io_out ? io_r_199_b : _GEN_20538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20540 = 10'hc8 == r_count_27_io_out ? io_r_200_b : _GEN_20539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20541 = 10'hc9 == r_count_27_io_out ? io_r_201_b : _GEN_20540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20542 = 10'hca == r_count_27_io_out ? io_r_202_b : _GEN_20541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20543 = 10'hcb == r_count_27_io_out ? io_r_203_b : _GEN_20542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20544 = 10'hcc == r_count_27_io_out ? io_r_204_b : _GEN_20543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20545 = 10'hcd == r_count_27_io_out ? io_r_205_b : _GEN_20544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20546 = 10'hce == r_count_27_io_out ? io_r_206_b : _GEN_20545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20547 = 10'hcf == r_count_27_io_out ? io_r_207_b : _GEN_20546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20548 = 10'hd0 == r_count_27_io_out ? io_r_208_b : _GEN_20547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20549 = 10'hd1 == r_count_27_io_out ? io_r_209_b : _GEN_20548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20550 = 10'hd2 == r_count_27_io_out ? io_r_210_b : _GEN_20549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20551 = 10'hd3 == r_count_27_io_out ? io_r_211_b : _GEN_20550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20552 = 10'hd4 == r_count_27_io_out ? io_r_212_b : _GEN_20551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20553 = 10'hd5 == r_count_27_io_out ? io_r_213_b : _GEN_20552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20554 = 10'hd6 == r_count_27_io_out ? io_r_214_b : _GEN_20553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20555 = 10'hd7 == r_count_27_io_out ? io_r_215_b : _GEN_20554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20556 = 10'hd8 == r_count_27_io_out ? io_r_216_b : _GEN_20555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20557 = 10'hd9 == r_count_27_io_out ? io_r_217_b : _GEN_20556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20558 = 10'hda == r_count_27_io_out ? io_r_218_b : _GEN_20557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20559 = 10'hdb == r_count_27_io_out ? io_r_219_b : _GEN_20558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20560 = 10'hdc == r_count_27_io_out ? io_r_220_b : _GEN_20559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20561 = 10'hdd == r_count_27_io_out ? io_r_221_b : _GEN_20560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20562 = 10'hde == r_count_27_io_out ? io_r_222_b : _GEN_20561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20563 = 10'hdf == r_count_27_io_out ? io_r_223_b : _GEN_20562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20564 = 10'he0 == r_count_27_io_out ? io_r_224_b : _GEN_20563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20565 = 10'he1 == r_count_27_io_out ? io_r_225_b : _GEN_20564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20566 = 10'he2 == r_count_27_io_out ? io_r_226_b : _GEN_20565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20567 = 10'he3 == r_count_27_io_out ? io_r_227_b : _GEN_20566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20568 = 10'he4 == r_count_27_io_out ? io_r_228_b : _GEN_20567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20569 = 10'he5 == r_count_27_io_out ? io_r_229_b : _GEN_20568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20570 = 10'he6 == r_count_27_io_out ? io_r_230_b : _GEN_20569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20571 = 10'he7 == r_count_27_io_out ? io_r_231_b : _GEN_20570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20572 = 10'he8 == r_count_27_io_out ? io_r_232_b : _GEN_20571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20573 = 10'he9 == r_count_27_io_out ? io_r_233_b : _GEN_20572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20574 = 10'hea == r_count_27_io_out ? io_r_234_b : _GEN_20573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20575 = 10'heb == r_count_27_io_out ? io_r_235_b : _GEN_20574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20576 = 10'hec == r_count_27_io_out ? io_r_236_b : _GEN_20575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20577 = 10'hed == r_count_27_io_out ? io_r_237_b : _GEN_20576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20578 = 10'hee == r_count_27_io_out ? io_r_238_b : _GEN_20577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20579 = 10'hef == r_count_27_io_out ? io_r_239_b : _GEN_20578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20580 = 10'hf0 == r_count_27_io_out ? io_r_240_b : _GEN_20579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20581 = 10'hf1 == r_count_27_io_out ? io_r_241_b : _GEN_20580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20582 = 10'hf2 == r_count_27_io_out ? io_r_242_b : _GEN_20581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20583 = 10'hf3 == r_count_27_io_out ? io_r_243_b : _GEN_20582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20584 = 10'hf4 == r_count_27_io_out ? io_r_244_b : _GEN_20583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20585 = 10'hf5 == r_count_27_io_out ? io_r_245_b : _GEN_20584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20586 = 10'hf6 == r_count_27_io_out ? io_r_246_b : _GEN_20585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20587 = 10'hf7 == r_count_27_io_out ? io_r_247_b : _GEN_20586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20588 = 10'hf8 == r_count_27_io_out ? io_r_248_b : _GEN_20587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20589 = 10'hf9 == r_count_27_io_out ? io_r_249_b : _GEN_20588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20590 = 10'hfa == r_count_27_io_out ? io_r_250_b : _GEN_20589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20591 = 10'hfb == r_count_27_io_out ? io_r_251_b : _GEN_20590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20592 = 10'hfc == r_count_27_io_out ? io_r_252_b : _GEN_20591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20593 = 10'hfd == r_count_27_io_out ? io_r_253_b : _GEN_20592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20594 = 10'hfe == r_count_27_io_out ? io_r_254_b : _GEN_20593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20595 = 10'hff == r_count_27_io_out ? io_r_255_b : _GEN_20594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20596 = 10'h100 == r_count_27_io_out ? io_r_256_b : _GEN_20595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20597 = 10'h101 == r_count_27_io_out ? io_r_257_b : _GEN_20596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20598 = 10'h102 == r_count_27_io_out ? io_r_258_b : _GEN_20597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20599 = 10'h103 == r_count_27_io_out ? io_r_259_b : _GEN_20598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20600 = 10'h104 == r_count_27_io_out ? io_r_260_b : _GEN_20599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20601 = 10'h105 == r_count_27_io_out ? io_r_261_b : _GEN_20600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20602 = 10'h106 == r_count_27_io_out ? io_r_262_b : _GEN_20601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20603 = 10'h107 == r_count_27_io_out ? io_r_263_b : _GEN_20602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20604 = 10'h108 == r_count_27_io_out ? io_r_264_b : _GEN_20603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20605 = 10'h109 == r_count_27_io_out ? io_r_265_b : _GEN_20604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20606 = 10'h10a == r_count_27_io_out ? io_r_266_b : _GEN_20605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20607 = 10'h10b == r_count_27_io_out ? io_r_267_b : _GEN_20606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20608 = 10'h10c == r_count_27_io_out ? io_r_268_b : _GEN_20607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20609 = 10'h10d == r_count_27_io_out ? io_r_269_b : _GEN_20608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20610 = 10'h10e == r_count_27_io_out ? io_r_270_b : _GEN_20609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20611 = 10'h10f == r_count_27_io_out ? io_r_271_b : _GEN_20610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20612 = 10'h110 == r_count_27_io_out ? io_r_272_b : _GEN_20611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20613 = 10'h111 == r_count_27_io_out ? io_r_273_b : _GEN_20612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20614 = 10'h112 == r_count_27_io_out ? io_r_274_b : _GEN_20613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20615 = 10'h113 == r_count_27_io_out ? io_r_275_b : _GEN_20614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20616 = 10'h114 == r_count_27_io_out ? io_r_276_b : _GEN_20615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20617 = 10'h115 == r_count_27_io_out ? io_r_277_b : _GEN_20616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20618 = 10'h116 == r_count_27_io_out ? io_r_278_b : _GEN_20617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20619 = 10'h117 == r_count_27_io_out ? io_r_279_b : _GEN_20618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20620 = 10'h118 == r_count_27_io_out ? io_r_280_b : _GEN_20619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20621 = 10'h119 == r_count_27_io_out ? io_r_281_b : _GEN_20620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20622 = 10'h11a == r_count_27_io_out ? io_r_282_b : _GEN_20621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20623 = 10'h11b == r_count_27_io_out ? io_r_283_b : _GEN_20622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20624 = 10'h11c == r_count_27_io_out ? io_r_284_b : _GEN_20623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20625 = 10'h11d == r_count_27_io_out ? io_r_285_b : _GEN_20624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20626 = 10'h11e == r_count_27_io_out ? io_r_286_b : _GEN_20625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20627 = 10'h11f == r_count_27_io_out ? io_r_287_b : _GEN_20626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20628 = 10'h120 == r_count_27_io_out ? io_r_288_b : _GEN_20627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20629 = 10'h121 == r_count_27_io_out ? io_r_289_b : _GEN_20628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20630 = 10'h122 == r_count_27_io_out ? io_r_290_b : _GEN_20629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20631 = 10'h123 == r_count_27_io_out ? io_r_291_b : _GEN_20630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20632 = 10'h124 == r_count_27_io_out ? io_r_292_b : _GEN_20631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20633 = 10'h125 == r_count_27_io_out ? io_r_293_b : _GEN_20632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20634 = 10'h126 == r_count_27_io_out ? io_r_294_b : _GEN_20633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20635 = 10'h127 == r_count_27_io_out ? io_r_295_b : _GEN_20634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20636 = 10'h128 == r_count_27_io_out ? io_r_296_b : _GEN_20635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20637 = 10'h129 == r_count_27_io_out ? io_r_297_b : _GEN_20636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20638 = 10'h12a == r_count_27_io_out ? io_r_298_b : _GEN_20637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20639 = 10'h12b == r_count_27_io_out ? io_r_299_b : _GEN_20638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20640 = 10'h12c == r_count_27_io_out ? io_r_300_b : _GEN_20639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20641 = 10'h12d == r_count_27_io_out ? io_r_301_b : _GEN_20640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20642 = 10'h12e == r_count_27_io_out ? io_r_302_b : _GEN_20641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20643 = 10'h12f == r_count_27_io_out ? io_r_303_b : _GEN_20642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20644 = 10'h130 == r_count_27_io_out ? io_r_304_b : _GEN_20643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20645 = 10'h131 == r_count_27_io_out ? io_r_305_b : _GEN_20644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20646 = 10'h132 == r_count_27_io_out ? io_r_306_b : _GEN_20645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20647 = 10'h133 == r_count_27_io_out ? io_r_307_b : _GEN_20646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20648 = 10'h134 == r_count_27_io_out ? io_r_308_b : _GEN_20647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20649 = 10'h135 == r_count_27_io_out ? io_r_309_b : _GEN_20648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20650 = 10'h136 == r_count_27_io_out ? io_r_310_b : _GEN_20649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20651 = 10'h137 == r_count_27_io_out ? io_r_311_b : _GEN_20650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20652 = 10'h138 == r_count_27_io_out ? io_r_312_b : _GEN_20651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20653 = 10'h139 == r_count_27_io_out ? io_r_313_b : _GEN_20652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20654 = 10'h13a == r_count_27_io_out ? io_r_314_b : _GEN_20653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20655 = 10'h13b == r_count_27_io_out ? io_r_315_b : _GEN_20654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20656 = 10'h13c == r_count_27_io_out ? io_r_316_b : _GEN_20655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20657 = 10'h13d == r_count_27_io_out ? io_r_317_b : _GEN_20656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20658 = 10'h13e == r_count_27_io_out ? io_r_318_b : _GEN_20657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20659 = 10'h13f == r_count_27_io_out ? io_r_319_b : _GEN_20658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20660 = 10'h140 == r_count_27_io_out ? io_r_320_b : _GEN_20659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20661 = 10'h141 == r_count_27_io_out ? io_r_321_b : _GEN_20660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20662 = 10'h142 == r_count_27_io_out ? io_r_322_b : _GEN_20661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20663 = 10'h143 == r_count_27_io_out ? io_r_323_b : _GEN_20662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20664 = 10'h144 == r_count_27_io_out ? io_r_324_b : _GEN_20663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20665 = 10'h145 == r_count_27_io_out ? io_r_325_b : _GEN_20664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20666 = 10'h146 == r_count_27_io_out ? io_r_326_b : _GEN_20665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20667 = 10'h147 == r_count_27_io_out ? io_r_327_b : _GEN_20666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20668 = 10'h148 == r_count_27_io_out ? io_r_328_b : _GEN_20667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20669 = 10'h149 == r_count_27_io_out ? io_r_329_b : _GEN_20668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20670 = 10'h14a == r_count_27_io_out ? io_r_330_b : _GEN_20669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20671 = 10'h14b == r_count_27_io_out ? io_r_331_b : _GEN_20670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20672 = 10'h14c == r_count_27_io_out ? io_r_332_b : _GEN_20671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20673 = 10'h14d == r_count_27_io_out ? io_r_333_b : _GEN_20672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20674 = 10'h14e == r_count_27_io_out ? io_r_334_b : _GEN_20673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20675 = 10'h14f == r_count_27_io_out ? io_r_335_b : _GEN_20674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20676 = 10'h150 == r_count_27_io_out ? io_r_336_b : _GEN_20675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20677 = 10'h151 == r_count_27_io_out ? io_r_337_b : _GEN_20676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20678 = 10'h152 == r_count_27_io_out ? io_r_338_b : _GEN_20677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20679 = 10'h153 == r_count_27_io_out ? io_r_339_b : _GEN_20678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20680 = 10'h154 == r_count_27_io_out ? io_r_340_b : _GEN_20679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20681 = 10'h155 == r_count_27_io_out ? io_r_341_b : _GEN_20680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20682 = 10'h156 == r_count_27_io_out ? io_r_342_b : _GEN_20681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20683 = 10'h157 == r_count_27_io_out ? io_r_343_b : _GEN_20682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20684 = 10'h158 == r_count_27_io_out ? io_r_344_b : _GEN_20683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20685 = 10'h159 == r_count_27_io_out ? io_r_345_b : _GEN_20684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20686 = 10'h15a == r_count_27_io_out ? io_r_346_b : _GEN_20685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20687 = 10'h15b == r_count_27_io_out ? io_r_347_b : _GEN_20686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20688 = 10'h15c == r_count_27_io_out ? io_r_348_b : _GEN_20687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20689 = 10'h15d == r_count_27_io_out ? io_r_349_b : _GEN_20688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20690 = 10'h15e == r_count_27_io_out ? io_r_350_b : _GEN_20689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20691 = 10'h15f == r_count_27_io_out ? io_r_351_b : _GEN_20690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20692 = 10'h160 == r_count_27_io_out ? io_r_352_b : _GEN_20691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20693 = 10'h161 == r_count_27_io_out ? io_r_353_b : _GEN_20692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20694 = 10'h162 == r_count_27_io_out ? io_r_354_b : _GEN_20693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20695 = 10'h163 == r_count_27_io_out ? io_r_355_b : _GEN_20694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20696 = 10'h164 == r_count_27_io_out ? io_r_356_b : _GEN_20695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20697 = 10'h165 == r_count_27_io_out ? io_r_357_b : _GEN_20696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20698 = 10'h166 == r_count_27_io_out ? io_r_358_b : _GEN_20697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20699 = 10'h167 == r_count_27_io_out ? io_r_359_b : _GEN_20698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20700 = 10'h168 == r_count_27_io_out ? io_r_360_b : _GEN_20699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20701 = 10'h169 == r_count_27_io_out ? io_r_361_b : _GEN_20700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20702 = 10'h16a == r_count_27_io_out ? io_r_362_b : _GEN_20701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20703 = 10'h16b == r_count_27_io_out ? io_r_363_b : _GEN_20702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20704 = 10'h16c == r_count_27_io_out ? io_r_364_b : _GEN_20703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20705 = 10'h16d == r_count_27_io_out ? io_r_365_b : _GEN_20704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20706 = 10'h16e == r_count_27_io_out ? io_r_366_b : _GEN_20705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20707 = 10'h16f == r_count_27_io_out ? io_r_367_b : _GEN_20706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20708 = 10'h170 == r_count_27_io_out ? io_r_368_b : _GEN_20707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20709 = 10'h171 == r_count_27_io_out ? io_r_369_b : _GEN_20708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20710 = 10'h172 == r_count_27_io_out ? io_r_370_b : _GEN_20709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20711 = 10'h173 == r_count_27_io_out ? io_r_371_b : _GEN_20710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20712 = 10'h174 == r_count_27_io_out ? io_r_372_b : _GEN_20711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20713 = 10'h175 == r_count_27_io_out ? io_r_373_b : _GEN_20712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20714 = 10'h176 == r_count_27_io_out ? io_r_374_b : _GEN_20713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20715 = 10'h177 == r_count_27_io_out ? io_r_375_b : _GEN_20714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20716 = 10'h178 == r_count_27_io_out ? io_r_376_b : _GEN_20715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20717 = 10'h179 == r_count_27_io_out ? io_r_377_b : _GEN_20716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20718 = 10'h17a == r_count_27_io_out ? io_r_378_b : _GEN_20717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20719 = 10'h17b == r_count_27_io_out ? io_r_379_b : _GEN_20718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20720 = 10'h17c == r_count_27_io_out ? io_r_380_b : _GEN_20719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20721 = 10'h17d == r_count_27_io_out ? io_r_381_b : _GEN_20720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20722 = 10'h17e == r_count_27_io_out ? io_r_382_b : _GEN_20721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20723 = 10'h17f == r_count_27_io_out ? io_r_383_b : _GEN_20722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20724 = 10'h180 == r_count_27_io_out ? io_r_384_b : _GEN_20723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20725 = 10'h181 == r_count_27_io_out ? io_r_385_b : _GEN_20724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20726 = 10'h182 == r_count_27_io_out ? io_r_386_b : _GEN_20725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20727 = 10'h183 == r_count_27_io_out ? io_r_387_b : _GEN_20726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20728 = 10'h184 == r_count_27_io_out ? io_r_388_b : _GEN_20727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20729 = 10'h185 == r_count_27_io_out ? io_r_389_b : _GEN_20728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20730 = 10'h186 == r_count_27_io_out ? io_r_390_b : _GEN_20729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20731 = 10'h187 == r_count_27_io_out ? io_r_391_b : _GEN_20730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20732 = 10'h188 == r_count_27_io_out ? io_r_392_b : _GEN_20731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20733 = 10'h189 == r_count_27_io_out ? io_r_393_b : _GEN_20732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20734 = 10'h18a == r_count_27_io_out ? io_r_394_b : _GEN_20733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20735 = 10'h18b == r_count_27_io_out ? io_r_395_b : _GEN_20734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20736 = 10'h18c == r_count_27_io_out ? io_r_396_b : _GEN_20735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20737 = 10'h18d == r_count_27_io_out ? io_r_397_b : _GEN_20736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20738 = 10'h18e == r_count_27_io_out ? io_r_398_b : _GEN_20737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20739 = 10'h18f == r_count_27_io_out ? io_r_399_b : _GEN_20738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20740 = 10'h190 == r_count_27_io_out ? io_r_400_b : _GEN_20739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20741 = 10'h191 == r_count_27_io_out ? io_r_401_b : _GEN_20740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20742 = 10'h192 == r_count_27_io_out ? io_r_402_b : _GEN_20741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20743 = 10'h193 == r_count_27_io_out ? io_r_403_b : _GEN_20742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20744 = 10'h194 == r_count_27_io_out ? io_r_404_b : _GEN_20743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20745 = 10'h195 == r_count_27_io_out ? io_r_405_b : _GEN_20744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20746 = 10'h196 == r_count_27_io_out ? io_r_406_b : _GEN_20745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20747 = 10'h197 == r_count_27_io_out ? io_r_407_b : _GEN_20746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20748 = 10'h198 == r_count_27_io_out ? io_r_408_b : _GEN_20747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20749 = 10'h199 == r_count_27_io_out ? io_r_409_b : _GEN_20748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20750 = 10'h19a == r_count_27_io_out ? io_r_410_b : _GEN_20749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20751 = 10'h19b == r_count_27_io_out ? io_r_411_b : _GEN_20750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20752 = 10'h19c == r_count_27_io_out ? io_r_412_b : _GEN_20751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20753 = 10'h19d == r_count_27_io_out ? io_r_413_b : _GEN_20752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20754 = 10'h19e == r_count_27_io_out ? io_r_414_b : _GEN_20753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20755 = 10'h19f == r_count_27_io_out ? io_r_415_b : _GEN_20754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20756 = 10'h1a0 == r_count_27_io_out ? io_r_416_b : _GEN_20755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20757 = 10'h1a1 == r_count_27_io_out ? io_r_417_b : _GEN_20756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20758 = 10'h1a2 == r_count_27_io_out ? io_r_418_b : _GEN_20757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20759 = 10'h1a3 == r_count_27_io_out ? io_r_419_b : _GEN_20758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20760 = 10'h1a4 == r_count_27_io_out ? io_r_420_b : _GEN_20759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20761 = 10'h1a5 == r_count_27_io_out ? io_r_421_b : _GEN_20760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20762 = 10'h1a6 == r_count_27_io_out ? io_r_422_b : _GEN_20761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20763 = 10'h1a7 == r_count_27_io_out ? io_r_423_b : _GEN_20762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20764 = 10'h1a8 == r_count_27_io_out ? io_r_424_b : _GEN_20763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20765 = 10'h1a9 == r_count_27_io_out ? io_r_425_b : _GEN_20764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20766 = 10'h1aa == r_count_27_io_out ? io_r_426_b : _GEN_20765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20767 = 10'h1ab == r_count_27_io_out ? io_r_427_b : _GEN_20766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20768 = 10'h1ac == r_count_27_io_out ? io_r_428_b : _GEN_20767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20769 = 10'h1ad == r_count_27_io_out ? io_r_429_b : _GEN_20768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20770 = 10'h1ae == r_count_27_io_out ? io_r_430_b : _GEN_20769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20771 = 10'h1af == r_count_27_io_out ? io_r_431_b : _GEN_20770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20772 = 10'h1b0 == r_count_27_io_out ? io_r_432_b : _GEN_20771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20773 = 10'h1b1 == r_count_27_io_out ? io_r_433_b : _GEN_20772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20774 = 10'h1b2 == r_count_27_io_out ? io_r_434_b : _GEN_20773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20775 = 10'h1b3 == r_count_27_io_out ? io_r_435_b : _GEN_20774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20776 = 10'h1b4 == r_count_27_io_out ? io_r_436_b : _GEN_20775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20777 = 10'h1b5 == r_count_27_io_out ? io_r_437_b : _GEN_20776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20778 = 10'h1b6 == r_count_27_io_out ? io_r_438_b : _GEN_20777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20779 = 10'h1b7 == r_count_27_io_out ? io_r_439_b : _GEN_20778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20780 = 10'h1b8 == r_count_27_io_out ? io_r_440_b : _GEN_20779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20781 = 10'h1b9 == r_count_27_io_out ? io_r_441_b : _GEN_20780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20782 = 10'h1ba == r_count_27_io_out ? io_r_442_b : _GEN_20781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20783 = 10'h1bb == r_count_27_io_out ? io_r_443_b : _GEN_20782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20784 = 10'h1bc == r_count_27_io_out ? io_r_444_b : _GEN_20783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20785 = 10'h1bd == r_count_27_io_out ? io_r_445_b : _GEN_20784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20786 = 10'h1be == r_count_27_io_out ? io_r_446_b : _GEN_20785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20787 = 10'h1bf == r_count_27_io_out ? io_r_447_b : _GEN_20786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20788 = 10'h1c0 == r_count_27_io_out ? io_r_448_b : _GEN_20787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20789 = 10'h1c1 == r_count_27_io_out ? io_r_449_b : _GEN_20788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20790 = 10'h1c2 == r_count_27_io_out ? io_r_450_b : _GEN_20789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20791 = 10'h1c3 == r_count_27_io_out ? io_r_451_b : _GEN_20790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20792 = 10'h1c4 == r_count_27_io_out ? io_r_452_b : _GEN_20791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20793 = 10'h1c5 == r_count_27_io_out ? io_r_453_b : _GEN_20792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20794 = 10'h1c6 == r_count_27_io_out ? io_r_454_b : _GEN_20793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20795 = 10'h1c7 == r_count_27_io_out ? io_r_455_b : _GEN_20794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20796 = 10'h1c8 == r_count_27_io_out ? io_r_456_b : _GEN_20795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20797 = 10'h1c9 == r_count_27_io_out ? io_r_457_b : _GEN_20796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20798 = 10'h1ca == r_count_27_io_out ? io_r_458_b : _GEN_20797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20799 = 10'h1cb == r_count_27_io_out ? io_r_459_b : _GEN_20798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20800 = 10'h1cc == r_count_27_io_out ? io_r_460_b : _GEN_20799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20801 = 10'h1cd == r_count_27_io_out ? io_r_461_b : _GEN_20800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20802 = 10'h1ce == r_count_27_io_out ? io_r_462_b : _GEN_20801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20803 = 10'h1cf == r_count_27_io_out ? io_r_463_b : _GEN_20802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20804 = 10'h1d0 == r_count_27_io_out ? io_r_464_b : _GEN_20803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20805 = 10'h1d1 == r_count_27_io_out ? io_r_465_b : _GEN_20804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20806 = 10'h1d2 == r_count_27_io_out ? io_r_466_b : _GEN_20805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20807 = 10'h1d3 == r_count_27_io_out ? io_r_467_b : _GEN_20806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20808 = 10'h1d4 == r_count_27_io_out ? io_r_468_b : _GEN_20807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20809 = 10'h1d5 == r_count_27_io_out ? io_r_469_b : _GEN_20808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20810 = 10'h1d6 == r_count_27_io_out ? io_r_470_b : _GEN_20809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20811 = 10'h1d7 == r_count_27_io_out ? io_r_471_b : _GEN_20810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20812 = 10'h1d8 == r_count_27_io_out ? io_r_472_b : _GEN_20811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20813 = 10'h1d9 == r_count_27_io_out ? io_r_473_b : _GEN_20812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20814 = 10'h1da == r_count_27_io_out ? io_r_474_b : _GEN_20813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20815 = 10'h1db == r_count_27_io_out ? io_r_475_b : _GEN_20814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20816 = 10'h1dc == r_count_27_io_out ? io_r_476_b : _GEN_20815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20817 = 10'h1dd == r_count_27_io_out ? io_r_477_b : _GEN_20816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20818 = 10'h1de == r_count_27_io_out ? io_r_478_b : _GEN_20817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20819 = 10'h1df == r_count_27_io_out ? io_r_479_b : _GEN_20818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20820 = 10'h1e0 == r_count_27_io_out ? io_r_480_b : _GEN_20819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20821 = 10'h1e1 == r_count_27_io_out ? io_r_481_b : _GEN_20820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20822 = 10'h1e2 == r_count_27_io_out ? io_r_482_b : _GEN_20821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20823 = 10'h1e3 == r_count_27_io_out ? io_r_483_b : _GEN_20822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20824 = 10'h1e4 == r_count_27_io_out ? io_r_484_b : _GEN_20823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20825 = 10'h1e5 == r_count_27_io_out ? io_r_485_b : _GEN_20824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20826 = 10'h1e6 == r_count_27_io_out ? io_r_486_b : _GEN_20825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20827 = 10'h1e7 == r_count_27_io_out ? io_r_487_b : _GEN_20826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20828 = 10'h1e8 == r_count_27_io_out ? io_r_488_b : _GEN_20827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20829 = 10'h1e9 == r_count_27_io_out ? io_r_489_b : _GEN_20828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20830 = 10'h1ea == r_count_27_io_out ? io_r_490_b : _GEN_20829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20831 = 10'h1eb == r_count_27_io_out ? io_r_491_b : _GEN_20830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20832 = 10'h1ec == r_count_27_io_out ? io_r_492_b : _GEN_20831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20833 = 10'h1ed == r_count_27_io_out ? io_r_493_b : _GEN_20832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20834 = 10'h1ee == r_count_27_io_out ? io_r_494_b : _GEN_20833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20835 = 10'h1ef == r_count_27_io_out ? io_r_495_b : _GEN_20834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20836 = 10'h1f0 == r_count_27_io_out ? io_r_496_b : _GEN_20835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20837 = 10'h1f1 == r_count_27_io_out ? io_r_497_b : _GEN_20836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20838 = 10'h1f2 == r_count_27_io_out ? io_r_498_b : _GEN_20837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20839 = 10'h1f3 == r_count_27_io_out ? io_r_499_b : _GEN_20838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20840 = 10'h1f4 == r_count_27_io_out ? io_r_500_b : _GEN_20839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20841 = 10'h1f5 == r_count_27_io_out ? io_r_501_b : _GEN_20840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20842 = 10'h1f6 == r_count_27_io_out ? io_r_502_b : _GEN_20841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20843 = 10'h1f7 == r_count_27_io_out ? io_r_503_b : _GEN_20842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20844 = 10'h1f8 == r_count_27_io_out ? io_r_504_b : _GEN_20843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20845 = 10'h1f9 == r_count_27_io_out ? io_r_505_b : _GEN_20844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20846 = 10'h1fa == r_count_27_io_out ? io_r_506_b : _GEN_20845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20847 = 10'h1fb == r_count_27_io_out ? io_r_507_b : _GEN_20846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20848 = 10'h1fc == r_count_27_io_out ? io_r_508_b : _GEN_20847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20849 = 10'h1fd == r_count_27_io_out ? io_r_509_b : _GEN_20848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20850 = 10'h1fe == r_count_27_io_out ? io_r_510_b : _GEN_20849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20851 = 10'h1ff == r_count_27_io_out ? io_r_511_b : _GEN_20850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20852 = 10'h200 == r_count_27_io_out ? io_r_512_b : _GEN_20851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20853 = 10'h201 == r_count_27_io_out ? io_r_513_b : _GEN_20852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20854 = 10'h202 == r_count_27_io_out ? io_r_514_b : _GEN_20853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20855 = 10'h203 == r_count_27_io_out ? io_r_515_b : _GEN_20854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20856 = 10'h204 == r_count_27_io_out ? io_r_516_b : _GEN_20855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20857 = 10'h205 == r_count_27_io_out ? io_r_517_b : _GEN_20856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20858 = 10'h206 == r_count_27_io_out ? io_r_518_b : _GEN_20857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20859 = 10'h207 == r_count_27_io_out ? io_r_519_b : _GEN_20858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20860 = 10'h208 == r_count_27_io_out ? io_r_520_b : _GEN_20859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20861 = 10'h209 == r_count_27_io_out ? io_r_521_b : _GEN_20860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20862 = 10'h20a == r_count_27_io_out ? io_r_522_b : _GEN_20861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20863 = 10'h20b == r_count_27_io_out ? io_r_523_b : _GEN_20862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20864 = 10'h20c == r_count_27_io_out ? io_r_524_b : _GEN_20863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20865 = 10'h20d == r_count_27_io_out ? io_r_525_b : _GEN_20864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20866 = 10'h20e == r_count_27_io_out ? io_r_526_b : _GEN_20865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20867 = 10'h20f == r_count_27_io_out ? io_r_527_b : _GEN_20866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20868 = 10'h210 == r_count_27_io_out ? io_r_528_b : _GEN_20867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20869 = 10'h211 == r_count_27_io_out ? io_r_529_b : _GEN_20868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20870 = 10'h212 == r_count_27_io_out ? io_r_530_b : _GEN_20869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20871 = 10'h213 == r_count_27_io_out ? io_r_531_b : _GEN_20870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20872 = 10'h214 == r_count_27_io_out ? io_r_532_b : _GEN_20871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20873 = 10'h215 == r_count_27_io_out ? io_r_533_b : _GEN_20872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20874 = 10'h216 == r_count_27_io_out ? io_r_534_b : _GEN_20873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20875 = 10'h217 == r_count_27_io_out ? io_r_535_b : _GEN_20874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20876 = 10'h218 == r_count_27_io_out ? io_r_536_b : _GEN_20875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20877 = 10'h219 == r_count_27_io_out ? io_r_537_b : _GEN_20876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20878 = 10'h21a == r_count_27_io_out ? io_r_538_b : _GEN_20877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20879 = 10'h21b == r_count_27_io_out ? io_r_539_b : _GEN_20878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20880 = 10'h21c == r_count_27_io_out ? io_r_540_b : _GEN_20879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20881 = 10'h21d == r_count_27_io_out ? io_r_541_b : _GEN_20880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20882 = 10'h21e == r_count_27_io_out ? io_r_542_b : _GEN_20881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20883 = 10'h21f == r_count_27_io_out ? io_r_543_b : _GEN_20882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20884 = 10'h220 == r_count_27_io_out ? io_r_544_b : _GEN_20883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20885 = 10'h221 == r_count_27_io_out ? io_r_545_b : _GEN_20884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20886 = 10'h222 == r_count_27_io_out ? io_r_546_b : _GEN_20885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20887 = 10'h223 == r_count_27_io_out ? io_r_547_b : _GEN_20886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20888 = 10'h224 == r_count_27_io_out ? io_r_548_b : _GEN_20887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20889 = 10'h225 == r_count_27_io_out ? io_r_549_b : _GEN_20888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20890 = 10'h226 == r_count_27_io_out ? io_r_550_b : _GEN_20889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20891 = 10'h227 == r_count_27_io_out ? io_r_551_b : _GEN_20890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20892 = 10'h228 == r_count_27_io_out ? io_r_552_b : _GEN_20891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20893 = 10'h229 == r_count_27_io_out ? io_r_553_b : _GEN_20892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20894 = 10'h22a == r_count_27_io_out ? io_r_554_b : _GEN_20893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20895 = 10'h22b == r_count_27_io_out ? io_r_555_b : _GEN_20894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20896 = 10'h22c == r_count_27_io_out ? io_r_556_b : _GEN_20895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20897 = 10'h22d == r_count_27_io_out ? io_r_557_b : _GEN_20896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20898 = 10'h22e == r_count_27_io_out ? io_r_558_b : _GEN_20897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20899 = 10'h22f == r_count_27_io_out ? io_r_559_b : _GEN_20898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20900 = 10'h230 == r_count_27_io_out ? io_r_560_b : _GEN_20899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20901 = 10'h231 == r_count_27_io_out ? io_r_561_b : _GEN_20900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20902 = 10'h232 == r_count_27_io_out ? io_r_562_b : _GEN_20901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20903 = 10'h233 == r_count_27_io_out ? io_r_563_b : _GEN_20902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20904 = 10'h234 == r_count_27_io_out ? io_r_564_b : _GEN_20903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20905 = 10'h235 == r_count_27_io_out ? io_r_565_b : _GEN_20904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20906 = 10'h236 == r_count_27_io_out ? io_r_566_b : _GEN_20905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20907 = 10'h237 == r_count_27_io_out ? io_r_567_b : _GEN_20906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20908 = 10'h238 == r_count_27_io_out ? io_r_568_b : _GEN_20907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20909 = 10'h239 == r_count_27_io_out ? io_r_569_b : _GEN_20908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20910 = 10'h23a == r_count_27_io_out ? io_r_570_b : _GEN_20909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20911 = 10'h23b == r_count_27_io_out ? io_r_571_b : _GEN_20910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20912 = 10'h23c == r_count_27_io_out ? io_r_572_b : _GEN_20911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20913 = 10'h23d == r_count_27_io_out ? io_r_573_b : _GEN_20912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20914 = 10'h23e == r_count_27_io_out ? io_r_574_b : _GEN_20913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20915 = 10'h23f == r_count_27_io_out ? io_r_575_b : _GEN_20914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20916 = 10'h240 == r_count_27_io_out ? io_r_576_b : _GEN_20915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20917 = 10'h241 == r_count_27_io_out ? io_r_577_b : _GEN_20916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20918 = 10'h242 == r_count_27_io_out ? io_r_578_b : _GEN_20917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20919 = 10'h243 == r_count_27_io_out ? io_r_579_b : _GEN_20918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20920 = 10'h244 == r_count_27_io_out ? io_r_580_b : _GEN_20919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20921 = 10'h245 == r_count_27_io_out ? io_r_581_b : _GEN_20920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20922 = 10'h246 == r_count_27_io_out ? io_r_582_b : _GEN_20921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20923 = 10'h247 == r_count_27_io_out ? io_r_583_b : _GEN_20922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20924 = 10'h248 == r_count_27_io_out ? io_r_584_b : _GEN_20923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20925 = 10'h249 == r_count_27_io_out ? io_r_585_b : _GEN_20924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20926 = 10'h24a == r_count_27_io_out ? io_r_586_b : _GEN_20925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20927 = 10'h24b == r_count_27_io_out ? io_r_587_b : _GEN_20926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20928 = 10'h24c == r_count_27_io_out ? io_r_588_b : _GEN_20927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20929 = 10'h24d == r_count_27_io_out ? io_r_589_b : _GEN_20928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20930 = 10'h24e == r_count_27_io_out ? io_r_590_b : _GEN_20929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20931 = 10'h24f == r_count_27_io_out ? io_r_591_b : _GEN_20930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20932 = 10'h250 == r_count_27_io_out ? io_r_592_b : _GEN_20931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20933 = 10'h251 == r_count_27_io_out ? io_r_593_b : _GEN_20932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20934 = 10'h252 == r_count_27_io_out ? io_r_594_b : _GEN_20933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20935 = 10'h253 == r_count_27_io_out ? io_r_595_b : _GEN_20934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20936 = 10'h254 == r_count_27_io_out ? io_r_596_b : _GEN_20935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20937 = 10'h255 == r_count_27_io_out ? io_r_597_b : _GEN_20936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20938 = 10'h256 == r_count_27_io_out ? io_r_598_b : _GEN_20937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20939 = 10'h257 == r_count_27_io_out ? io_r_599_b : _GEN_20938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20940 = 10'h258 == r_count_27_io_out ? io_r_600_b : _GEN_20939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20941 = 10'h259 == r_count_27_io_out ? io_r_601_b : _GEN_20940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20942 = 10'h25a == r_count_27_io_out ? io_r_602_b : _GEN_20941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20943 = 10'h25b == r_count_27_io_out ? io_r_603_b : _GEN_20942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20944 = 10'h25c == r_count_27_io_out ? io_r_604_b : _GEN_20943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20945 = 10'h25d == r_count_27_io_out ? io_r_605_b : _GEN_20944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20946 = 10'h25e == r_count_27_io_out ? io_r_606_b : _GEN_20945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20947 = 10'h25f == r_count_27_io_out ? io_r_607_b : _GEN_20946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20948 = 10'h260 == r_count_27_io_out ? io_r_608_b : _GEN_20947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20949 = 10'h261 == r_count_27_io_out ? io_r_609_b : _GEN_20948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20950 = 10'h262 == r_count_27_io_out ? io_r_610_b : _GEN_20949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20951 = 10'h263 == r_count_27_io_out ? io_r_611_b : _GEN_20950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20952 = 10'h264 == r_count_27_io_out ? io_r_612_b : _GEN_20951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20953 = 10'h265 == r_count_27_io_out ? io_r_613_b : _GEN_20952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20954 = 10'h266 == r_count_27_io_out ? io_r_614_b : _GEN_20953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20955 = 10'h267 == r_count_27_io_out ? io_r_615_b : _GEN_20954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20956 = 10'h268 == r_count_27_io_out ? io_r_616_b : _GEN_20955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20957 = 10'h269 == r_count_27_io_out ? io_r_617_b : _GEN_20956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20958 = 10'h26a == r_count_27_io_out ? io_r_618_b : _GEN_20957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20959 = 10'h26b == r_count_27_io_out ? io_r_619_b : _GEN_20958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20960 = 10'h26c == r_count_27_io_out ? io_r_620_b : _GEN_20959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20961 = 10'h26d == r_count_27_io_out ? io_r_621_b : _GEN_20960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20962 = 10'h26e == r_count_27_io_out ? io_r_622_b : _GEN_20961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20963 = 10'h26f == r_count_27_io_out ? io_r_623_b : _GEN_20962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20964 = 10'h270 == r_count_27_io_out ? io_r_624_b : _GEN_20963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20965 = 10'h271 == r_count_27_io_out ? io_r_625_b : _GEN_20964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20966 = 10'h272 == r_count_27_io_out ? io_r_626_b : _GEN_20965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20967 = 10'h273 == r_count_27_io_out ? io_r_627_b : _GEN_20966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20968 = 10'h274 == r_count_27_io_out ? io_r_628_b : _GEN_20967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20969 = 10'h275 == r_count_27_io_out ? io_r_629_b : _GEN_20968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20970 = 10'h276 == r_count_27_io_out ? io_r_630_b : _GEN_20969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20971 = 10'h277 == r_count_27_io_out ? io_r_631_b : _GEN_20970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20972 = 10'h278 == r_count_27_io_out ? io_r_632_b : _GEN_20971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20973 = 10'h279 == r_count_27_io_out ? io_r_633_b : _GEN_20972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20974 = 10'h27a == r_count_27_io_out ? io_r_634_b : _GEN_20973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20975 = 10'h27b == r_count_27_io_out ? io_r_635_b : _GEN_20974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20976 = 10'h27c == r_count_27_io_out ? io_r_636_b : _GEN_20975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20977 = 10'h27d == r_count_27_io_out ? io_r_637_b : _GEN_20976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20978 = 10'h27e == r_count_27_io_out ? io_r_638_b : _GEN_20977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20979 = 10'h27f == r_count_27_io_out ? io_r_639_b : _GEN_20978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20980 = 10'h280 == r_count_27_io_out ? io_r_640_b : _GEN_20979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20981 = 10'h281 == r_count_27_io_out ? io_r_641_b : _GEN_20980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20982 = 10'h282 == r_count_27_io_out ? io_r_642_b : _GEN_20981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20983 = 10'h283 == r_count_27_io_out ? io_r_643_b : _GEN_20982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20984 = 10'h284 == r_count_27_io_out ? io_r_644_b : _GEN_20983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20985 = 10'h285 == r_count_27_io_out ? io_r_645_b : _GEN_20984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20986 = 10'h286 == r_count_27_io_out ? io_r_646_b : _GEN_20985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20987 = 10'h287 == r_count_27_io_out ? io_r_647_b : _GEN_20986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20988 = 10'h288 == r_count_27_io_out ? io_r_648_b : _GEN_20987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20989 = 10'h289 == r_count_27_io_out ? io_r_649_b : _GEN_20988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20990 = 10'h28a == r_count_27_io_out ? io_r_650_b : _GEN_20989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20991 = 10'h28b == r_count_27_io_out ? io_r_651_b : _GEN_20990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20992 = 10'h28c == r_count_27_io_out ? io_r_652_b : _GEN_20991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20993 = 10'h28d == r_count_27_io_out ? io_r_653_b : _GEN_20992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20994 = 10'h28e == r_count_27_io_out ? io_r_654_b : _GEN_20993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20995 = 10'h28f == r_count_27_io_out ? io_r_655_b : _GEN_20994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20996 = 10'h290 == r_count_27_io_out ? io_r_656_b : _GEN_20995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20997 = 10'h291 == r_count_27_io_out ? io_r_657_b : _GEN_20996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20998 = 10'h292 == r_count_27_io_out ? io_r_658_b : _GEN_20997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20999 = 10'h293 == r_count_27_io_out ? io_r_659_b : _GEN_20998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21000 = 10'h294 == r_count_27_io_out ? io_r_660_b : _GEN_20999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21001 = 10'h295 == r_count_27_io_out ? io_r_661_b : _GEN_21000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21002 = 10'h296 == r_count_27_io_out ? io_r_662_b : _GEN_21001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21003 = 10'h297 == r_count_27_io_out ? io_r_663_b : _GEN_21002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21004 = 10'h298 == r_count_27_io_out ? io_r_664_b : _GEN_21003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21005 = 10'h299 == r_count_27_io_out ? io_r_665_b : _GEN_21004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21006 = 10'h29a == r_count_27_io_out ? io_r_666_b : _GEN_21005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21007 = 10'h29b == r_count_27_io_out ? io_r_667_b : _GEN_21006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21008 = 10'h29c == r_count_27_io_out ? io_r_668_b : _GEN_21007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21009 = 10'h29d == r_count_27_io_out ? io_r_669_b : _GEN_21008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21010 = 10'h29e == r_count_27_io_out ? io_r_670_b : _GEN_21009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21011 = 10'h29f == r_count_27_io_out ? io_r_671_b : _GEN_21010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21012 = 10'h2a0 == r_count_27_io_out ? io_r_672_b : _GEN_21011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21013 = 10'h2a1 == r_count_27_io_out ? io_r_673_b : _GEN_21012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21014 = 10'h2a2 == r_count_27_io_out ? io_r_674_b : _GEN_21013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21015 = 10'h2a3 == r_count_27_io_out ? io_r_675_b : _GEN_21014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21016 = 10'h2a4 == r_count_27_io_out ? io_r_676_b : _GEN_21015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21017 = 10'h2a5 == r_count_27_io_out ? io_r_677_b : _GEN_21016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21018 = 10'h2a6 == r_count_27_io_out ? io_r_678_b : _GEN_21017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21019 = 10'h2a7 == r_count_27_io_out ? io_r_679_b : _GEN_21018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21020 = 10'h2a8 == r_count_27_io_out ? io_r_680_b : _GEN_21019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21021 = 10'h2a9 == r_count_27_io_out ? io_r_681_b : _GEN_21020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21022 = 10'h2aa == r_count_27_io_out ? io_r_682_b : _GEN_21021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21023 = 10'h2ab == r_count_27_io_out ? io_r_683_b : _GEN_21022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21024 = 10'h2ac == r_count_27_io_out ? io_r_684_b : _GEN_21023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21025 = 10'h2ad == r_count_27_io_out ? io_r_685_b : _GEN_21024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21026 = 10'h2ae == r_count_27_io_out ? io_r_686_b : _GEN_21025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21027 = 10'h2af == r_count_27_io_out ? io_r_687_b : _GEN_21026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21028 = 10'h2b0 == r_count_27_io_out ? io_r_688_b : _GEN_21027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21029 = 10'h2b1 == r_count_27_io_out ? io_r_689_b : _GEN_21028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21030 = 10'h2b2 == r_count_27_io_out ? io_r_690_b : _GEN_21029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21031 = 10'h2b3 == r_count_27_io_out ? io_r_691_b : _GEN_21030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21032 = 10'h2b4 == r_count_27_io_out ? io_r_692_b : _GEN_21031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21033 = 10'h2b5 == r_count_27_io_out ? io_r_693_b : _GEN_21032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21034 = 10'h2b6 == r_count_27_io_out ? io_r_694_b : _GEN_21033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21035 = 10'h2b7 == r_count_27_io_out ? io_r_695_b : _GEN_21034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21036 = 10'h2b8 == r_count_27_io_out ? io_r_696_b : _GEN_21035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21037 = 10'h2b9 == r_count_27_io_out ? io_r_697_b : _GEN_21036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21038 = 10'h2ba == r_count_27_io_out ? io_r_698_b : _GEN_21037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21039 = 10'h2bb == r_count_27_io_out ? io_r_699_b : _GEN_21038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21040 = 10'h2bc == r_count_27_io_out ? io_r_700_b : _GEN_21039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21041 = 10'h2bd == r_count_27_io_out ? io_r_701_b : _GEN_21040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21042 = 10'h2be == r_count_27_io_out ? io_r_702_b : _GEN_21041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21043 = 10'h2bf == r_count_27_io_out ? io_r_703_b : _GEN_21042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21044 = 10'h2c0 == r_count_27_io_out ? io_r_704_b : _GEN_21043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21045 = 10'h2c1 == r_count_27_io_out ? io_r_705_b : _GEN_21044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21046 = 10'h2c2 == r_count_27_io_out ? io_r_706_b : _GEN_21045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21047 = 10'h2c3 == r_count_27_io_out ? io_r_707_b : _GEN_21046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21048 = 10'h2c4 == r_count_27_io_out ? io_r_708_b : _GEN_21047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21049 = 10'h2c5 == r_count_27_io_out ? io_r_709_b : _GEN_21048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21050 = 10'h2c6 == r_count_27_io_out ? io_r_710_b : _GEN_21049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21051 = 10'h2c7 == r_count_27_io_out ? io_r_711_b : _GEN_21050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21052 = 10'h2c8 == r_count_27_io_out ? io_r_712_b : _GEN_21051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21053 = 10'h2c9 == r_count_27_io_out ? io_r_713_b : _GEN_21052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21054 = 10'h2ca == r_count_27_io_out ? io_r_714_b : _GEN_21053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21055 = 10'h2cb == r_count_27_io_out ? io_r_715_b : _GEN_21054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21056 = 10'h2cc == r_count_27_io_out ? io_r_716_b : _GEN_21055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21057 = 10'h2cd == r_count_27_io_out ? io_r_717_b : _GEN_21056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21058 = 10'h2ce == r_count_27_io_out ? io_r_718_b : _GEN_21057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21059 = 10'h2cf == r_count_27_io_out ? io_r_719_b : _GEN_21058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21060 = 10'h2d0 == r_count_27_io_out ? io_r_720_b : _GEN_21059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21061 = 10'h2d1 == r_count_27_io_out ? io_r_721_b : _GEN_21060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21062 = 10'h2d2 == r_count_27_io_out ? io_r_722_b : _GEN_21061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21063 = 10'h2d3 == r_count_27_io_out ? io_r_723_b : _GEN_21062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21064 = 10'h2d4 == r_count_27_io_out ? io_r_724_b : _GEN_21063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21065 = 10'h2d5 == r_count_27_io_out ? io_r_725_b : _GEN_21064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21066 = 10'h2d6 == r_count_27_io_out ? io_r_726_b : _GEN_21065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21067 = 10'h2d7 == r_count_27_io_out ? io_r_727_b : _GEN_21066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21068 = 10'h2d8 == r_count_27_io_out ? io_r_728_b : _GEN_21067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21069 = 10'h2d9 == r_count_27_io_out ? io_r_729_b : _GEN_21068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21070 = 10'h2da == r_count_27_io_out ? io_r_730_b : _GEN_21069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21071 = 10'h2db == r_count_27_io_out ? io_r_731_b : _GEN_21070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21072 = 10'h2dc == r_count_27_io_out ? io_r_732_b : _GEN_21071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21073 = 10'h2dd == r_count_27_io_out ? io_r_733_b : _GEN_21072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21074 = 10'h2de == r_count_27_io_out ? io_r_734_b : _GEN_21073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21075 = 10'h2df == r_count_27_io_out ? io_r_735_b : _GEN_21074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21076 = 10'h2e0 == r_count_27_io_out ? io_r_736_b : _GEN_21075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21077 = 10'h2e1 == r_count_27_io_out ? io_r_737_b : _GEN_21076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21078 = 10'h2e2 == r_count_27_io_out ? io_r_738_b : _GEN_21077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21079 = 10'h2e3 == r_count_27_io_out ? io_r_739_b : _GEN_21078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21080 = 10'h2e4 == r_count_27_io_out ? io_r_740_b : _GEN_21079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21081 = 10'h2e5 == r_count_27_io_out ? io_r_741_b : _GEN_21080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21082 = 10'h2e6 == r_count_27_io_out ? io_r_742_b : _GEN_21081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21083 = 10'h2e7 == r_count_27_io_out ? io_r_743_b : _GEN_21082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21084 = 10'h2e8 == r_count_27_io_out ? io_r_744_b : _GEN_21083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21085 = 10'h2e9 == r_count_27_io_out ? io_r_745_b : _GEN_21084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21086 = 10'h2ea == r_count_27_io_out ? io_r_746_b : _GEN_21085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21087 = 10'h2eb == r_count_27_io_out ? io_r_747_b : _GEN_21086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21088 = 10'h2ec == r_count_27_io_out ? io_r_748_b : _GEN_21087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21091 = 10'h1 == r_count_28_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21092 = 10'h2 == r_count_28_io_out ? io_r_2_b : _GEN_21091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21093 = 10'h3 == r_count_28_io_out ? io_r_3_b : _GEN_21092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21094 = 10'h4 == r_count_28_io_out ? io_r_4_b : _GEN_21093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21095 = 10'h5 == r_count_28_io_out ? io_r_5_b : _GEN_21094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21096 = 10'h6 == r_count_28_io_out ? io_r_6_b : _GEN_21095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21097 = 10'h7 == r_count_28_io_out ? io_r_7_b : _GEN_21096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21098 = 10'h8 == r_count_28_io_out ? io_r_8_b : _GEN_21097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21099 = 10'h9 == r_count_28_io_out ? io_r_9_b : _GEN_21098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21100 = 10'ha == r_count_28_io_out ? io_r_10_b : _GEN_21099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21101 = 10'hb == r_count_28_io_out ? io_r_11_b : _GEN_21100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21102 = 10'hc == r_count_28_io_out ? io_r_12_b : _GEN_21101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21103 = 10'hd == r_count_28_io_out ? io_r_13_b : _GEN_21102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21104 = 10'he == r_count_28_io_out ? io_r_14_b : _GEN_21103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21105 = 10'hf == r_count_28_io_out ? io_r_15_b : _GEN_21104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21106 = 10'h10 == r_count_28_io_out ? io_r_16_b : _GEN_21105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21107 = 10'h11 == r_count_28_io_out ? io_r_17_b : _GEN_21106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21108 = 10'h12 == r_count_28_io_out ? io_r_18_b : _GEN_21107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21109 = 10'h13 == r_count_28_io_out ? io_r_19_b : _GEN_21108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21110 = 10'h14 == r_count_28_io_out ? io_r_20_b : _GEN_21109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21111 = 10'h15 == r_count_28_io_out ? io_r_21_b : _GEN_21110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21112 = 10'h16 == r_count_28_io_out ? io_r_22_b : _GEN_21111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21113 = 10'h17 == r_count_28_io_out ? io_r_23_b : _GEN_21112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21114 = 10'h18 == r_count_28_io_out ? io_r_24_b : _GEN_21113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21115 = 10'h19 == r_count_28_io_out ? io_r_25_b : _GEN_21114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21116 = 10'h1a == r_count_28_io_out ? io_r_26_b : _GEN_21115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21117 = 10'h1b == r_count_28_io_out ? io_r_27_b : _GEN_21116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21118 = 10'h1c == r_count_28_io_out ? io_r_28_b : _GEN_21117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21119 = 10'h1d == r_count_28_io_out ? io_r_29_b : _GEN_21118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21120 = 10'h1e == r_count_28_io_out ? io_r_30_b : _GEN_21119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21121 = 10'h1f == r_count_28_io_out ? io_r_31_b : _GEN_21120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21122 = 10'h20 == r_count_28_io_out ? io_r_32_b : _GEN_21121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21123 = 10'h21 == r_count_28_io_out ? io_r_33_b : _GEN_21122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21124 = 10'h22 == r_count_28_io_out ? io_r_34_b : _GEN_21123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21125 = 10'h23 == r_count_28_io_out ? io_r_35_b : _GEN_21124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21126 = 10'h24 == r_count_28_io_out ? io_r_36_b : _GEN_21125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21127 = 10'h25 == r_count_28_io_out ? io_r_37_b : _GEN_21126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21128 = 10'h26 == r_count_28_io_out ? io_r_38_b : _GEN_21127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21129 = 10'h27 == r_count_28_io_out ? io_r_39_b : _GEN_21128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21130 = 10'h28 == r_count_28_io_out ? io_r_40_b : _GEN_21129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21131 = 10'h29 == r_count_28_io_out ? io_r_41_b : _GEN_21130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21132 = 10'h2a == r_count_28_io_out ? io_r_42_b : _GEN_21131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21133 = 10'h2b == r_count_28_io_out ? io_r_43_b : _GEN_21132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21134 = 10'h2c == r_count_28_io_out ? io_r_44_b : _GEN_21133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21135 = 10'h2d == r_count_28_io_out ? io_r_45_b : _GEN_21134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21136 = 10'h2e == r_count_28_io_out ? io_r_46_b : _GEN_21135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21137 = 10'h2f == r_count_28_io_out ? io_r_47_b : _GEN_21136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21138 = 10'h30 == r_count_28_io_out ? io_r_48_b : _GEN_21137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21139 = 10'h31 == r_count_28_io_out ? io_r_49_b : _GEN_21138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21140 = 10'h32 == r_count_28_io_out ? io_r_50_b : _GEN_21139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21141 = 10'h33 == r_count_28_io_out ? io_r_51_b : _GEN_21140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21142 = 10'h34 == r_count_28_io_out ? io_r_52_b : _GEN_21141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21143 = 10'h35 == r_count_28_io_out ? io_r_53_b : _GEN_21142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21144 = 10'h36 == r_count_28_io_out ? io_r_54_b : _GEN_21143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21145 = 10'h37 == r_count_28_io_out ? io_r_55_b : _GEN_21144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21146 = 10'h38 == r_count_28_io_out ? io_r_56_b : _GEN_21145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21147 = 10'h39 == r_count_28_io_out ? io_r_57_b : _GEN_21146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21148 = 10'h3a == r_count_28_io_out ? io_r_58_b : _GEN_21147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21149 = 10'h3b == r_count_28_io_out ? io_r_59_b : _GEN_21148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21150 = 10'h3c == r_count_28_io_out ? io_r_60_b : _GEN_21149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21151 = 10'h3d == r_count_28_io_out ? io_r_61_b : _GEN_21150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21152 = 10'h3e == r_count_28_io_out ? io_r_62_b : _GEN_21151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21153 = 10'h3f == r_count_28_io_out ? io_r_63_b : _GEN_21152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21154 = 10'h40 == r_count_28_io_out ? io_r_64_b : _GEN_21153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21155 = 10'h41 == r_count_28_io_out ? io_r_65_b : _GEN_21154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21156 = 10'h42 == r_count_28_io_out ? io_r_66_b : _GEN_21155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21157 = 10'h43 == r_count_28_io_out ? io_r_67_b : _GEN_21156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21158 = 10'h44 == r_count_28_io_out ? io_r_68_b : _GEN_21157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21159 = 10'h45 == r_count_28_io_out ? io_r_69_b : _GEN_21158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21160 = 10'h46 == r_count_28_io_out ? io_r_70_b : _GEN_21159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21161 = 10'h47 == r_count_28_io_out ? io_r_71_b : _GEN_21160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21162 = 10'h48 == r_count_28_io_out ? io_r_72_b : _GEN_21161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21163 = 10'h49 == r_count_28_io_out ? io_r_73_b : _GEN_21162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21164 = 10'h4a == r_count_28_io_out ? io_r_74_b : _GEN_21163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21165 = 10'h4b == r_count_28_io_out ? io_r_75_b : _GEN_21164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21166 = 10'h4c == r_count_28_io_out ? io_r_76_b : _GEN_21165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21167 = 10'h4d == r_count_28_io_out ? io_r_77_b : _GEN_21166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21168 = 10'h4e == r_count_28_io_out ? io_r_78_b : _GEN_21167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21169 = 10'h4f == r_count_28_io_out ? io_r_79_b : _GEN_21168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21170 = 10'h50 == r_count_28_io_out ? io_r_80_b : _GEN_21169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21171 = 10'h51 == r_count_28_io_out ? io_r_81_b : _GEN_21170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21172 = 10'h52 == r_count_28_io_out ? io_r_82_b : _GEN_21171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21173 = 10'h53 == r_count_28_io_out ? io_r_83_b : _GEN_21172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21174 = 10'h54 == r_count_28_io_out ? io_r_84_b : _GEN_21173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21175 = 10'h55 == r_count_28_io_out ? io_r_85_b : _GEN_21174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21176 = 10'h56 == r_count_28_io_out ? io_r_86_b : _GEN_21175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21177 = 10'h57 == r_count_28_io_out ? io_r_87_b : _GEN_21176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21178 = 10'h58 == r_count_28_io_out ? io_r_88_b : _GEN_21177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21179 = 10'h59 == r_count_28_io_out ? io_r_89_b : _GEN_21178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21180 = 10'h5a == r_count_28_io_out ? io_r_90_b : _GEN_21179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21181 = 10'h5b == r_count_28_io_out ? io_r_91_b : _GEN_21180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21182 = 10'h5c == r_count_28_io_out ? io_r_92_b : _GEN_21181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21183 = 10'h5d == r_count_28_io_out ? io_r_93_b : _GEN_21182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21184 = 10'h5e == r_count_28_io_out ? io_r_94_b : _GEN_21183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21185 = 10'h5f == r_count_28_io_out ? io_r_95_b : _GEN_21184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21186 = 10'h60 == r_count_28_io_out ? io_r_96_b : _GEN_21185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21187 = 10'h61 == r_count_28_io_out ? io_r_97_b : _GEN_21186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21188 = 10'h62 == r_count_28_io_out ? io_r_98_b : _GEN_21187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21189 = 10'h63 == r_count_28_io_out ? io_r_99_b : _GEN_21188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21190 = 10'h64 == r_count_28_io_out ? io_r_100_b : _GEN_21189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21191 = 10'h65 == r_count_28_io_out ? io_r_101_b : _GEN_21190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21192 = 10'h66 == r_count_28_io_out ? io_r_102_b : _GEN_21191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21193 = 10'h67 == r_count_28_io_out ? io_r_103_b : _GEN_21192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21194 = 10'h68 == r_count_28_io_out ? io_r_104_b : _GEN_21193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21195 = 10'h69 == r_count_28_io_out ? io_r_105_b : _GEN_21194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21196 = 10'h6a == r_count_28_io_out ? io_r_106_b : _GEN_21195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21197 = 10'h6b == r_count_28_io_out ? io_r_107_b : _GEN_21196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21198 = 10'h6c == r_count_28_io_out ? io_r_108_b : _GEN_21197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21199 = 10'h6d == r_count_28_io_out ? io_r_109_b : _GEN_21198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21200 = 10'h6e == r_count_28_io_out ? io_r_110_b : _GEN_21199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21201 = 10'h6f == r_count_28_io_out ? io_r_111_b : _GEN_21200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21202 = 10'h70 == r_count_28_io_out ? io_r_112_b : _GEN_21201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21203 = 10'h71 == r_count_28_io_out ? io_r_113_b : _GEN_21202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21204 = 10'h72 == r_count_28_io_out ? io_r_114_b : _GEN_21203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21205 = 10'h73 == r_count_28_io_out ? io_r_115_b : _GEN_21204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21206 = 10'h74 == r_count_28_io_out ? io_r_116_b : _GEN_21205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21207 = 10'h75 == r_count_28_io_out ? io_r_117_b : _GEN_21206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21208 = 10'h76 == r_count_28_io_out ? io_r_118_b : _GEN_21207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21209 = 10'h77 == r_count_28_io_out ? io_r_119_b : _GEN_21208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21210 = 10'h78 == r_count_28_io_out ? io_r_120_b : _GEN_21209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21211 = 10'h79 == r_count_28_io_out ? io_r_121_b : _GEN_21210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21212 = 10'h7a == r_count_28_io_out ? io_r_122_b : _GEN_21211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21213 = 10'h7b == r_count_28_io_out ? io_r_123_b : _GEN_21212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21214 = 10'h7c == r_count_28_io_out ? io_r_124_b : _GEN_21213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21215 = 10'h7d == r_count_28_io_out ? io_r_125_b : _GEN_21214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21216 = 10'h7e == r_count_28_io_out ? io_r_126_b : _GEN_21215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21217 = 10'h7f == r_count_28_io_out ? io_r_127_b : _GEN_21216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21218 = 10'h80 == r_count_28_io_out ? io_r_128_b : _GEN_21217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21219 = 10'h81 == r_count_28_io_out ? io_r_129_b : _GEN_21218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21220 = 10'h82 == r_count_28_io_out ? io_r_130_b : _GEN_21219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21221 = 10'h83 == r_count_28_io_out ? io_r_131_b : _GEN_21220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21222 = 10'h84 == r_count_28_io_out ? io_r_132_b : _GEN_21221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21223 = 10'h85 == r_count_28_io_out ? io_r_133_b : _GEN_21222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21224 = 10'h86 == r_count_28_io_out ? io_r_134_b : _GEN_21223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21225 = 10'h87 == r_count_28_io_out ? io_r_135_b : _GEN_21224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21226 = 10'h88 == r_count_28_io_out ? io_r_136_b : _GEN_21225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21227 = 10'h89 == r_count_28_io_out ? io_r_137_b : _GEN_21226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21228 = 10'h8a == r_count_28_io_out ? io_r_138_b : _GEN_21227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21229 = 10'h8b == r_count_28_io_out ? io_r_139_b : _GEN_21228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21230 = 10'h8c == r_count_28_io_out ? io_r_140_b : _GEN_21229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21231 = 10'h8d == r_count_28_io_out ? io_r_141_b : _GEN_21230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21232 = 10'h8e == r_count_28_io_out ? io_r_142_b : _GEN_21231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21233 = 10'h8f == r_count_28_io_out ? io_r_143_b : _GEN_21232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21234 = 10'h90 == r_count_28_io_out ? io_r_144_b : _GEN_21233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21235 = 10'h91 == r_count_28_io_out ? io_r_145_b : _GEN_21234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21236 = 10'h92 == r_count_28_io_out ? io_r_146_b : _GEN_21235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21237 = 10'h93 == r_count_28_io_out ? io_r_147_b : _GEN_21236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21238 = 10'h94 == r_count_28_io_out ? io_r_148_b : _GEN_21237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21239 = 10'h95 == r_count_28_io_out ? io_r_149_b : _GEN_21238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21240 = 10'h96 == r_count_28_io_out ? io_r_150_b : _GEN_21239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21241 = 10'h97 == r_count_28_io_out ? io_r_151_b : _GEN_21240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21242 = 10'h98 == r_count_28_io_out ? io_r_152_b : _GEN_21241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21243 = 10'h99 == r_count_28_io_out ? io_r_153_b : _GEN_21242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21244 = 10'h9a == r_count_28_io_out ? io_r_154_b : _GEN_21243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21245 = 10'h9b == r_count_28_io_out ? io_r_155_b : _GEN_21244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21246 = 10'h9c == r_count_28_io_out ? io_r_156_b : _GEN_21245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21247 = 10'h9d == r_count_28_io_out ? io_r_157_b : _GEN_21246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21248 = 10'h9e == r_count_28_io_out ? io_r_158_b : _GEN_21247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21249 = 10'h9f == r_count_28_io_out ? io_r_159_b : _GEN_21248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21250 = 10'ha0 == r_count_28_io_out ? io_r_160_b : _GEN_21249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21251 = 10'ha1 == r_count_28_io_out ? io_r_161_b : _GEN_21250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21252 = 10'ha2 == r_count_28_io_out ? io_r_162_b : _GEN_21251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21253 = 10'ha3 == r_count_28_io_out ? io_r_163_b : _GEN_21252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21254 = 10'ha4 == r_count_28_io_out ? io_r_164_b : _GEN_21253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21255 = 10'ha5 == r_count_28_io_out ? io_r_165_b : _GEN_21254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21256 = 10'ha6 == r_count_28_io_out ? io_r_166_b : _GEN_21255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21257 = 10'ha7 == r_count_28_io_out ? io_r_167_b : _GEN_21256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21258 = 10'ha8 == r_count_28_io_out ? io_r_168_b : _GEN_21257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21259 = 10'ha9 == r_count_28_io_out ? io_r_169_b : _GEN_21258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21260 = 10'haa == r_count_28_io_out ? io_r_170_b : _GEN_21259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21261 = 10'hab == r_count_28_io_out ? io_r_171_b : _GEN_21260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21262 = 10'hac == r_count_28_io_out ? io_r_172_b : _GEN_21261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21263 = 10'had == r_count_28_io_out ? io_r_173_b : _GEN_21262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21264 = 10'hae == r_count_28_io_out ? io_r_174_b : _GEN_21263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21265 = 10'haf == r_count_28_io_out ? io_r_175_b : _GEN_21264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21266 = 10'hb0 == r_count_28_io_out ? io_r_176_b : _GEN_21265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21267 = 10'hb1 == r_count_28_io_out ? io_r_177_b : _GEN_21266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21268 = 10'hb2 == r_count_28_io_out ? io_r_178_b : _GEN_21267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21269 = 10'hb3 == r_count_28_io_out ? io_r_179_b : _GEN_21268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21270 = 10'hb4 == r_count_28_io_out ? io_r_180_b : _GEN_21269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21271 = 10'hb5 == r_count_28_io_out ? io_r_181_b : _GEN_21270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21272 = 10'hb6 == r_count_28_io_out ? io_r_182_b : _GEN_21271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21273 = 10'hb7 == r_count_28_io_out ? io_r_183_b : _GEN_21272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21274 = 10'hb8 == r_count_28_io_out ? io_r_184_b : _GEN_21273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21275 = 10'hb9 == r_count_28_io_out ? io_r_185_b : _GEN_21274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21276 = 10'hba == r_count_28_io_out ? io_r_186_b : _GEN_21275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21277 = 10'hbb == r_count_28_io_out ? io_r_187_b : _GEN_21276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21278 = 10'hbc == r_count_28_io_out ? io_r_188_b : _GEN_21277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21279 = 10'hbd == r_count_28_io_out ? io_r_189_b : _GEN_21278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21280 = 10'hbe == r_count_28_io_out ? io_r_190_b : _GEN_21279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21281 = 10'hbf == r_count_28_io_out ? io_r_191_b : _GEN_21280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21282 = 10'hc0 == r_count_28_io_out ? io_r_192_b : _GEN_21281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21283 = 10'hc1 == r_count_28_io_out ? io_r_193_b : _GEN_21282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21284 = 10'hc2 == r_count_28_io_out ? io_r_194_b : _GEN_21283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21285 = 10'hc3 == r_count_28_io_out ? io_r_195_b : _GEN_21284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21286 = 10'hc4 == r_count_28_io_out ? io_r_196_b : _GEN_21285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21287 = 10'hc5 == r_count_28_io_out ? io_r_197_b : _GEN_21286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21288 = 10'hc6 == r_count_28_io_out ? io_r_198_b : _GEN_21287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21289 = 10'hc7 == r_count_28_io_out ? io_r_199_b : _GEN_21288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21290 = 10'hc8 == r_count_28_io_out ? io_r_200_b : _GEN_21289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21291 = 10'hc9 == r_count_28_io_out ? io_r_201_b : _GEN_21290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21292 = 10'hca == r_count_28_io_out ? io_r_202_b : _GEN_21291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21293 = 10'hcb == r_count_28_io_out ? io_r_203_b : _GEN_21292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21294 = 10'hcc == r_count_28_io_out ? io_r_204_b : _GEN_21293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21295 = 10'hcd == r_count_28_io_out ? io_r_205_b : _GEN_21294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21296 = 10'hce == r_count_28_io_out ? io_r_206_b : _GEN_21295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21297 = 10'hcf == r_count_28_io_out ? io_r_207_b : _GEN_21296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21298 = 10'hd0 == r_count_28_io_out ? io_r_208_b : _GEN_21297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21299 = 10'hd1 == r_count_28_io_out ? io_r_209_b : _GEN_21298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21300 = 10'hd2 == r_count_28_io_out ? io_r_210_b : _GEN_21299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21301 = 10'hd3 == r_count_28_io_out ? io_r_211_b : _GEN_21300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21302 = 10'hd4 == r_count_28_io_out ? io_r_212_b : _GEN_21301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21303 = 10'hd5 == r_count_28_io_out ? io_r_213_b : _GEN_21302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21304 = 10'hd6 == r_count_28_io_out ? io_r_214_b : _GEN_21303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21305 = 10'hd7 == r_count_28_io_out ? io_r_215_b : _GEN_21304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21306 = 10'hd8 == r_count_28_io_out ? io_r_216_b : _GEN_21305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21307 = 10'hd9 == r_count_28_io_out ? io_r_217_b : _GEN_21306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21308 = 10'hda == r_count_28_io_out ? io_r_218_b : _GEN_21307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21309 = 10'hdb == r_count_28_io_out ? io_r_219_b : _GEN_21308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21310 = 10'hdc == r_count_28_io_out ? io_r_220_b : _GEN_21309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21311 = 10'hdd == r_count_28_io_out ? io_r_221_b : _GEN_21310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21312 = 10'hde == r_count_28_io_out ? io_r_222_b : _GEN_21311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21313 = 10'hdf == r_count_28_io_out ? io_r_223_b : _GEN_21312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21314 = 10'he0 == r_count_28_io_out ? io_r_224_b : _GEN_21313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21315 = 10'he1 == r_count_28_io_out ? io_r_225_b : _GEN_21314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21316 = 10'he2 == r_count_28_io_out ? io_r_226_b : _GEN_21315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21317 = 10'he3 == r_count_28_io_out ? io_r_227_b : _GEN_21316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21318 = 10'he4 == r_count_28_io_out ? io_r_228_b : _GEN_21317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21319 = 10'he5 == r_count_28_io_out ? io_r_229_b : _GEN_21318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21320 = 10'he6 == r_count_28_io_out ? io_r_230_b : _GEN_21319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21321 = 10'he7 == r_count_28_io_out ? io_r_231_b : _GEN_21320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21322 = 10'he8 == r_count_28_io_out ? io_r_232_b : _GEN_21321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21323 = 10'he9 == r_count_28_io_out ? io_r_233_b : _GEN_21322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21324 = 10'hea == r_count_28_io_out ? io_r_234_b : _GEN_21323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21325 = 10'heb == r_count_28_io_out ? io_r_235_b : _GEN_21324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21326 = 10'hec == r_count_28_io_out ? io_r_236_b : _GEN_21325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21327 = 10'hed == r_count_28_io_out ? io_r_237_b : _GEN_21326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21328 = 10'hee == r_count_28_io_out ? io_r_238_b : _GEN_21327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21329 = 10'hef == r_count_28_io_out ? io_r_239_b : _GEN_21328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21330 = 10'hf0 == r_count_28_io_out ? io_r_240_b : _GEN_21329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21331 = 10'hf1 == r_count_28_io_out ? io_r_241_b : _GEN_21330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21332 = 10'hf2 == r_count_28_io_out ? io_r_242_b : _GEN_21331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21333 = 10'hf3 == r_count_28_io_out ? io_r_243_b : _GEN_21332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21334 = 10'hf4 == r_count_28_io_out ? io_r_244_b : _GEN_21333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21335 = 10'hf5 == r_count_28_io_out ? io_r_245_b : _GEN_21334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21336 = 10'hf6 == r_count_28_io_out ? io_r_246_b : _GEN_21335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21337 = 10'hf7 == r_count_28_io_out ? io_r_247_b : _GEN_21336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21338 = 10'hf8 == r_count_28_io_out ? io_r_248_b : _GEN_21337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21339 = 10'hf9 == r_count_28_io_out ? io_r_249_b : _GEN_21338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21340 = 10'hfa == r_count_28_io_out ? io_r_250_b : _GEN_21339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21341 = 10'hfb == r_count_28_io_out ? io_r_251_b : _GEN_21340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21342 = 10'hfc == r_count_28_io_out ? io_r_252_b : _GEN_21341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21343 = 10'hfd == r_count_28_io_out ? io_r_253_b : _GEN_21342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21344 = 10'hfe == r_count_28_io_out ? io_r_254_b : _GEN_21343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21345 = 10'hff == r_count_28_io_out ? io_r_255_b : _GEN_21344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21346 = 10'h100 == r_count_28_io_out ? io_r_256_b : _GEN_21345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21347 = 10'h101 == r_count_28_io_out ? io_r_257_b : _GEN_21346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21348 = 10'h102 == r_count_28_io_out ? io_r_258_b : _GEN_21347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21349 = 10'h103 == r_count_28_io_out ? io_r_259_b : _GEN_21348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21350 = 10'h104 == r_count_28_io_out ? io_r_260_b : _GEN_21349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21351 = 10'h105 == r_count_28_io_out ? io_r_261_b : _GEN_21350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21352 = 10'h106 == r_count_28_io_out ? io_r_262_b : _GEN_21351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21353 = 10'h107 == r_count_28_io_out ? io_r_263_b : _GEN_21352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21354 = 10'h108 == r_count_28_io_out ? io_r_264_b : _GEN_21353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21355 = 10'h109 == r_count_28_io_out ? io_r_265_b : _GEN_21354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21356 = 10'h10a == r_count_28_io_out ? io_r_266_b : _GEN_21355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21357 = 10'h10b == r_count_28_io_out ? io_r_267_b : _GEN_21356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21358 = 10'h10c == r_count_28_io_out ? io_r_268_b : _GEN_21357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21359 = 10'h10d == r_count_28_io_out ? io_r_269_b : _GEN_21358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21360 = 10'h10e == r_count_28_io_out ? io_r_270_b : _GEN_21359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21361 = 10'h10f == r_count_28_io_out ? io_r_271_b : _GEN_21360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21362 = 10'h110 == r_count_28_io_out ? io_r_272_b : _GEN_21361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21363 = 10'h111 == r_count_28_io_out ? io_r_273_b : _GEN_21362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21364 = 10'h112 == r_count_28_io_out ? io_r_274_b : _GEN_21363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21365 = 10'h113 == r_count_28_io_out ? io_r_275_b : _GEN_21364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21366 = 10'h114 == r_count_28_io_out ? io_r_276_b : _GEN_21365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21367 = 10'h115 == r_count_28_io_out ? io_r_277_b : _GEN_21366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21368 = 10'h116 == r_count_28_io_out ? io_r_278_b : _GEN_21367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21369 = 10'h117 == r_count_28_io_out ? io_r_279_b : _GEN_21368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21370 = 10'h118 == r_count_28_io_out ? io_r_280_b : _GEN_21369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21371 = 10'h119 == r_count_28_io_out ? io_r_281_b : _GEN_21370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21372 = 10'h11a == r_count_28_io_out ? io_r_282_b : _GEN_21371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21373 = 10'h11b == r_count_28_io_out ? io_r_283_b : _GEN_21372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21374 = 10'h11c == r_count_28_io_out ? io_r_284_b : _GEN_21373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21375 = 10'h11d == r_count_28_io_out ? io_r_285_b : _GEN_21374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21376 = 10'h11e == r_count_28_io_out ? io_r_286_b : _GEN_21375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21377 = 10'h11f == r_count_28_io_out ? io_r_287_b : _GEN_21376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21378 = 10'h120 == r_count_28_io_out ? io_r_288_b : _GEN_21377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21379 = 10'h121 == r_count_28_io_out ? io_r_289_b : _GEN_21378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21380 = 10'h122 == r_count_28_io_out ? io_r_290_b : _GEN_21379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21381 = 10'h123 == r_count_28_io_out ? io_r_291_b : _GEN_21380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21382 = 10'h124 == r_count_28_io_out ? io_r_292_b : _GEN_21381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21383 = 10'h125 == r_count_28_io_out ? io_r_293_b : _GEN_21382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21384 = 10'h126 == r_count_28_io_out ? io_r_294_b : _GEN_21383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21385 = 10'h127 == r_count_28_io_out ? io_r_295_b : _GEN_21384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21386 = 10'h128 == r_count_28_io_out ? io_r_296_b : _GEN_21385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21387 = 10'h129 == r_count_28_io_out ? io_r_297_b : _GEN_21386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21388 = 10'h12a == r_count_28_io_out ? io_r_298_b : _GEN_21387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21389 = 10'h12b == r_count_28_io_out ? io_r_299_b : _GEN_21388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21390 = 10'h12c == r_count_28_io_out ? io_r_300_b : _GEN_21389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21391 = 10'h12d == r_count_28_io_out ? io_r_301_b : _GEN_21390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21392 = 10'h12e == r_count_28_io_out ? io_r_302_b : _GEN_21391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21393 = 10'h12f == r_count_28_io_out ? io_r_303_b : _GEN_21392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21394 = 10'h130 == r_count_28_io_out ? io_r_304_b : _GEN_21393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21395 = 10'h131 == r_count_28_io_out ? io_r_305_b : _GEN_21394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21396 = 10'h132 == r_count_28_io_out ? io_r_306_b : _GEN_21395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21397 = 10'h133 == r_count_28_io_out ? io_r_307_b : _GEN_21396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21398 = 10'h134 == r_count_28_io_out ? io_r_308_b : _GEN_21397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21399 = 10'h135 == r_count_28_io_out ? io_r_309_b : _GEN_21398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21400 = 10'h136 == r_count_28_io_out ? io_r_310_b : _GEN_21399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21401 = 10'h137 == r_count_28_io_out ? io_r_311_b : _GEN_21400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21402 = 10'h138 == r_count_28_io_out ? io_r_312_b : _GEN_21401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21403 = 10'h139 == r_count_28_io_out ? io_r_313_b : _GEN_21402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21404 = 10'h13a == r_count_28_io_out ? io_r_314_b : _GEN_21403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21405 = 10'h13b == r_count_28_io_out ? io_r_315_b : _GEN_21404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21406 = 10'h13c == r_count_28_io_out ? io_r_316_b : _GEN_21405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21407 = 10'h13d == r_count_28_io_out ? io_r_317_b : _GEN_21406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21408 = 10'h13e == r_count_28_io_out ? io_r_318_b : _GEN_21407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21409 = 10'h13f == r_count_28_io_out ? io_r_319_b : _GEN_21408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21410 = 10'h140 == r_count_28_io_out ? io_r_320_b : _GEN_21409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21411 = 10'h141 == r_count_28_io_out ? io_r_321_b : _GEN_21410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21412 = 10'h142 == r_count_28_io_out ? io_r_322_b : _GEN_21411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21413 = 10'h143 == r_count_28_io_out ? io_r_323_b : _GEN_21412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21414 = 10'h144 == r_count_28_io_out ? io_r_324_b : _GEN_21413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21415 = 10'h145 == r_count_28_io_out ? io_r_325_b : _GEN_21414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21416 = 10'h146 == r_count_28_io_out ? io_r_326_b : _GEN_21415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21417 = 10'h147 == r_count_28_io_out ? io_r_327_b : _GEN_21416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21418 = 10'h148 == r_count_28_io_out ? io_r_328_b : _GEN_21417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21419 = 10'h149 == r_count_28_io_out ? io_r_329_b : _GEN_21418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21420 = 10'h14a == r_count_28_io_out ? io_r_330_b : _GEN_21419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21421 = 10'h14b == r_count_28_io_out ? io_r_331_b : _GEN_21420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21422 = 10'h14c == r_count_28_io_out ? io_r_332_b : _GEN_21421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21423 = 10'h14d == r_count_28_io_out ? io_r_333_b : _GEN_21422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21424 = 10'h14e == r_count_28_io_out ? io_r_334_b : _GEN_21423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21425 = 10'h14f == r_count_28_io_out ? io_r_335_b : _GEN_21424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21426 = 10'h150 == r_count_28_io_out ? io_r_336_b : _GEN_21425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21427 = 10'h151 == r_count_28_io_out ? io_r_337_b : _GEN_21426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21428 = 10'h152 == r_count_28_io_out ? io_r_338_b : _GEN_21427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21429 = 10'h153 == r_count_28_io_out ? io_r_339_b : _GEN_21428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21430 = 10'h154 == r_count_28_io_out ? io_r_340_b : _GEN_21429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21431 = 10'h155 == r_count_28_io_out ? io_r_341_b : _GEN_21430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21432 = 10'h156 == r_count_28_io_out ? io_r_342_b : _GEN_21431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21433 = 10'h157 == r_count_28_io_out ? io_r_343_b : _GEN_21432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21434 = 10'h158 == r_count_28_io_out ? io_r_344_b : _GEN_21433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21435 = 10'h159 == r_count_28_io_out ? io_r_345_b : _GEN_21434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21436 = 10'h15a == r_count_28_io_out ? io_r_346_b : _GEN_21435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21437 = 10'h15b == r_count_28_io_out ? io_r_347_b : _GEN_21436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21438 = 10'h15c == r_count_28_io_out ? io_r_348_b : _GEN_21437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21439 = 10'h15d == r_count_28_io_out ? io_r_349_b : _GEN_21438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21440 = 10'h15e == r_count_28_io_out ? io_r_350_b : _GEN_21439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21441 = 10'h15f == r_count_28_io_out ? io_r_351_b : _GEN_21440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21442 = 10'h160 == r_count_28_io_out ? io_r_352_b : _GEN_21441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21443 = 10'h161 == r_count_28_io_out ? io_r_353_b : _GEN_21442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21444 = 10'h162 == r_count_28_io_out ? io_r_354_b : _GEN_21443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21445 = 10'h163 == r_count_28_io_out ? io_r_355_b : _GEN_21444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21446 = 10'h164 == r_count_28_io_out ? io_r_356_b : _GEN_21445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21447 = 10'h165 == r_count_28_io_out ? io_r_357_b : _GEN_21446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21448 = 10'h166 == r_count_28_io_out ? io_r_358_b : _GEN_21447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21449 = 10'h167 == r_count_28_io_out ? io_r_359_b : _GEN_21448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21450 = 10'h168 == r_count_28_io_out ? io_r_360_b : _GEN_21449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21451 = 10'h169 == r_count_28_io_out ? io_r_361_b : _GEN_21450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21452 = 10'h16a == r_count_28_io_out ? io_r_362_b : _GEN_21451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21453 = 10'h16b == r_count_28_io_out ? io_r_363_b : _GEN_21452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21454 = 10'h16c == r_count_28_io_out ? io_r_364_b : _GEN_21453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21455 = 10'h16d == r_count_28_io_out ? io_r_365_b : _GEN_21454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21456 = 10'h16e == r_count_28_io_out ? io_r_366_b : _GEN_21455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21457 = 10'h16f == r_count_28_io_out ? io_r_367_b : _GEN_21456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21458 = 10'h170 == r_count_28_io_out ? io_r_368_b : _GEN_21457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21459 = 10'h171 == r_count_28_io_out ? io_r_369_b : _GEN_21458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21460 = 10'h172 == r_count_28_io_out ? io_r_370_b : _GEN_21459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21461 = 10'h173 == r_count_28_io_out ? io_r_371_b : _GEN_21460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21462 = 10'h174 == r_count_28_io_out ? io_r_372_b : _GEN_21461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21463 = 10'h175 == r_count_28_io_out ? io_r_373_b : _GEN_21462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21464 = 10'h176 == r_count_28_io_out ? io_r_374_b : _GEN_21463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21465 = 10'h177 == r_count_28_io_out ? io_r_375_b : _GEN_21464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21466 = 10'h178 == r_count_28_io_out ? io_r_376_b : _GEN_21465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21467 = 10'h179 == r_count_28_io_out ? io_r_377_b : _GEN_21466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21468 = 10'h17a == r_count_28_io_out ? io_r_378_b : _GEN_21467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21469 = 10'h17b == r_count_28_io_out ? io_r_379_b : _GEN_21468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21470 = 10'h17c == r_count_28_io_out ? io_r_380_b : _GEN_21469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21471 = 10'h17d == r_count_28_io_out ? io_r_381_b : _GEN_21470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21472 = 10'h17e == r_count_28_io_out ? io_r_382_b : _GEN_21471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21473 = 10'h17f == r_count_28_io_out ? io_r_383_b : _GEN_21472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21474 = 10'h180 == r_count_28_io_out ? io_r_384_b : _GEN_21473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21475 = 10'h181 == r_count_28_io_out ? io_r_385_b : _GEN_21474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21476 = 10'h182 == r_count_28_io_out ? io_r_386_b : _GEN_21475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21477 = 10'h183 == r_count_28_io_out ? io_r_387_b : _GEN_21476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21478 = 10'h184 == r_count_28_io_out ? io_r_388_b : _GEN_21477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21479 = 10'h185 == r_count_28_io_out ? io_r_389_b : _GEN_21478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21480 = 10'h186 == r_count_28_io_out ? io_r_390_b : _GEN_21479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21481 = 10'h187 == r_count_28_io_out ? io_r_391_b : _GEN_21480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21482 = 10'h188 == r_count_28_io_out ? io_r_392_b : _GEN_21481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21483 = 10'h189 == r_count_28_io_out ? io_r_393_b : _GEN_21482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21484 = 10'h18a == r_count_28_io_out ? io_r_394_b : _GEN_21483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21485 = 10'h18b == r_count_28_io_out ? io_r_395_b : _GEN_21484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21486 = 10'h18c == r_count_28_io_out ? io_r_396_b : _GEN_21485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21487 = 10'h18d == r_count_28_io_out ? io_r_397_b : _GEN_21486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21488 = 10'h18e == r_count_28_io_out ? io_r_398_b : _GEN_21487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21489 = 10'h18f == r_count_28_io_out ? io_r_399_b : _GEN_21488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21490 = 10'h190 == r_count_28_io_out ? io_r_400_b : _GEN_21489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21491 = 10'h191 == r_count_28_io_out ? io_r_401_b : _GEN_21490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21492 = 10'h192 == r_count_28_io_out ? io_r_402_b : _GEN_21491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21493 = 10'h193 == r_count_28_io_out ? io_r_403_b : _GEN_21492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21494 = 10'h194 == r_count_28_io_out ? io_r_404_b : _GEN_21493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21495 = 10'h195 == r_count_28_io_out ? io_r_405_b : _GEN_21494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21496 = 10'h196 == r_count_28_io_out ? io_r_406_b : _GEN_21495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21497 = 10'h197 == r_count_28_io_out ? io_r_407_b : _GEN_21496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21498 = 10'h198 == r_count_28_io_out ? io_r_408_b : _GEN_21497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21499 = 10'h199 == r_count_28_io_out ? io_r_409_b : _GEN_21498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21500 = 10'h19a == r_count_28_io_out ? io_r_410_b : _GEN_21499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21501 = 10'h19b == r_count_28_io_out ? io_r_411_b : _GEN_21500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21502 = 10'h19c == r_count_28_io_out ? io_r_412_b : _GEN_21501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21503 = 10'h19d == r_count_28_io_out ? io_r_413_b : _GEN_21502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21504 = 10'h19e == r_count_28_io_out ? io_r_414_b : _GEN_21503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21505 = 10'h19f == r_count_28_io_out ? io_r_415_b : _GEN_21504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21506 = 10'h1a0 == r_count_28_io_out ? io_r_416_b : _GEN_21505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21507 = 10'h1a1 == r_count_28_io_out ? io_r_417_b : _GEN_21506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21508 = 10'h1a2 == r_count_28_io_out ? io_r_418_b : _GEN_21507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21509 = 10'h1a3 == r_count_28_io_out ? io_r_419_b : _GEN_21508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21510 = 10'h1a4 == r_count_28_io_out ? io_r_420_b : _GEN_21509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21511 = 10'h1a5 == r_count_28_io_out ? io_r_421_b : _GEN_21510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21512 = 10'h1a6 == r_count_28_io_out ? io_r_422_b : _GEN_21511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21513 = 10'h1a7 == r_count_28_io_out ? io_r_423_b : _GEN_21512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21514 = 10'h1a8 == r_count_28_io_out ? io_r_424_b : _GEN_21513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21515 = 10'h1a9 == r_count_28_io_out ? io_r_425_b : _GEN_21514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21516 = 10'h1aa == r_count_28_io_out ? io_r_426_b : _GEN_21515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21517 = 10'h1ab == r_count_28_io_out ? io_r_427_b : _GEN_21516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21518 = 10'h1ac == r_count_28_io_out ? io_r_428_b : _GEN_21517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21519 = 10'h1ad == r_count_28_io_out ? io_r_429_b : _GEN_21518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21520 = 10'h1ae == r_count_28_io_out ? io_r_430_b : _GEN_21519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21521 = 10'h1af == r_count_28_io_out ? io_r_431_b : _GEN_21520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21522 = 10'h1b0 == r_count_28_io_out ? io_r_432_b : _GEN_21521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21523 = 10'h1b1 == r_count_28_io_out ? io_r_433_b : _GEN_21522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21524 = 10'h1b2 == r_count_28_io_out ? io_r_434_b : _GEN_21523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21525 = 10'h1b3 == r_count_28_io_out ? io_r_435_b : _GEN_21524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21526 = 10'h1b4 == r_count_28_io_out ? io_r_436_b : _GEN_21525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21527 = 10'h1b5 == r_count_28_io_out ? io_r_437_b : _GEN_21526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21528 = 10'h1b6 == r_count_28_io_out ? io_r_438_b : _GEN_21527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21529 = 10'h1b7 == r_count_28_io_out ? io_r_439_b : _GEN_21528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21530 = 10'h1b8 == r_count_28_io_out ? io_r_440_b : _GEN_21529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21531 = 10'h1b9 == r_count_28_io_out ? io_r_441_b : _GEN_21530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21532 = 10'h1ba == r_count_28_io_out ? io_r_442_b : _GEN_21531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21533 = 10'h1bb == r_count_28_io_out ? io_r_443_b : _GEN_21532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21534 = 10'h1bc == r_count_28_io_out ? io_r_444_b : _GEN_21533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21535 = 10'h1bd == r_count_28_io_out ? io_r_445_b : _GEN_21534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21536 = 10'h1be == r_count_28_io_out ? io_r_446_b : _GEN_21535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21537 = 10'h1bf == r_count_28_io_out ? io_r_447_b : _GEN_21536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21538 = 10'h1c0 == r_count_28_io_out ? io_r_448_b : _GEN_21537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21539 = 10'h1c1 == r_count_28_io_out ? io_r_449_b : _GEN_21538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21540 = 10'h1c2 == r_count_28_io_out ? io_r_450_b : _GEN_21539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21541 = 10'h1c3 == r_count_28_io_out ? io_r_451_b : _GEN_21540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21542 = 10'h1c4 == r_count_28_io_out ? io_r_452_b : _GEN_21541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21543 = 10'h1c5 == r_count_28_io_out ? io_r_453_b : _GEN_21542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21544 = 10'h1c6 == r_count_28_io_out ? io_r_454_b : _GEN_21543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21545 = 10'h1c7 == r_count_28_io_out ? io_r_455_b : _GEN_21544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21546 = 10'h1c8 == r_count_28_io_out ? io_r_456_b : _GEN_21545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21547 = 10'h1c9 == r_count_28_io_out ? io_r_457_b : _GEN_21546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21548 = 10'h1ca == r_count_28_io_out ? io_r_458_b : _GEN_21547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21549 = 10'h1cb == r_count_28_io_out ? io_r_459_b : _GEN_21548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21550 = 10'h1cc == r_count_28_io_out ? io_r_460_b : _GEN_21549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21551 = 10'h1cd == r_count_28_io_out ? io_r_461_b : _GEN_21550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21552 = 10'h1ce == r_count_28_io_out ? io_r_462_b : _GEN_21551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21553 = 10'h1cf == r_count_28_io_out ? io_r_463_b : _GEN_21552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21554 = 10'h1d0 == r_count_28_io_out ? io_r_464_b : _GEN_21553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21555 = 10'h1d1 == r_count_28_io_out ? io_r_465_b : _GEN_21554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21556 = 10'h1d2 == r_count_28_io_out ? io_r_466_b : _GEN_21555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21557 = 10'h1d3 == r_count_28_io_out ? io_r_467_b : _GEN_21556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21558 = 10'h1d4 == r_count_28_io_out ? io_r_468_b : _GEN_21557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21559 = 10'h1d5 == r_count_28_io_out ? io_r_469_b : _GEN_21558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21560 = 10'h1d6 == r_count_28_io_out ? io_r_470_b : _GEN_21559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21561 = 10'h1d7 == r_count_28_io_out ? io_r_471_b : _GEN_21560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21562 = 10'h1d8 == r_count_28_io_out ? io_r_472_b : _GEN_21561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21563 = 10'h1d9 == r_count_28_io_out ? io_r_473_b : _GEN_21562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21564 = 10'h1da == r_count_28_io_out ? io_r_474_b : _GEN_21563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21565 = 10'h1db == r_count_28_io_out ? io_r_475_b : _GEN_21564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21566 = 10'h1dc == r_count_28_io_out ? io_r_476_b : _GEN_21565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21567 = 10'h1dd == r_count_28_io_out ? io_r_477_b : _GEN_21566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21568 = 10'h1de == r_count_28_io_out ? io_r_478_b : _GEN_21567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21569 = 10'h1df == r_count_28_io_out ? io_r_479_b : _GEN_21568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21570 = 10'h1e0 == r_count_28_io_out ? io_r_480_b : _GEN_21569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21571 = 10'h1e1 == r_count_28_io_out ? io_r_481_b : _GEN_21570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21572 = 10'h1e2 == r_count_28_io_out ? io_r_482_b : _GEN_21571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21573 = 10'h1e3 == r_count_28_io_out ? io_r_483_b : _GEN_21572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21574 = 10'h1e4 == r_count_28_io_out ? io_r_484_b : _GEN_21573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21575 = 10'h1e5 == r_count_28_io_out ? io_r_485_b : _GEN_21574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21576 = 10'h1e6 == r_count_28_io_out ? io_r_486_b : _GEN_21575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21577 = 10'h1e7 == r_count_28_io_out ? io_r_487_b : _GEN_21576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21578 = 10'h1e8 == r_count_28_io_out ? io_r_488_b : _GEN_21577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21579 = 10'h1e9 == r_count_28_io_out ? io_r_489_b : _GEN_21578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21580 = 10'h1ea == r_count_28_io_out ? io_r_490_b : _GEN_21579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21581 = 10'h1eb == r_count_28_io_out ? io_r_491_b : _GEN_21580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21582 = 10'h1ec == r_count_28_io_out ? io_r_492_b : _GEN_21581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21583 = 10'h1ed == r_count_28_io_out ? io_r_493_b : _GEN_21582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21584 = 10'h1ee == r_count_28_io_out ? io_r_494_b : _GEN_21583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21585 = 10'h1ef == r_count_28_io_out ? io_r_495_b : _GEN_21584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21586 = 10'h1f0 == r_count_28_io_out ? io_r_496_b : _GEN_21585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21587 = 10'h1f1 == r_count_28_io_out ? io_r_497_b : _GEN_21586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21588 = 10'h1f2 == r_count_28_io_out ? io_r_498_b : _GEN_21587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21589 = 10'h1f3 == r_count_28_io_out ? io_r_499_b : _GEN_21588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21590 = 10'h1f4 == r_count_28_io_out ? io_r_500_b : _GEN_21589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21591 = 10'h1f5 == r_count_28_io_out ? io_r_501_b : _GEN_21590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21592 = 10'h1f6 == r_count_28_io_out ? io_r_502_b : _GEN_21591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21593 = 10'h1f7 == r_count_28_io_out ? io_r_503_b : _GEN_21592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21594 = 10'h1f8 == r_count_28_io_out ? io_r_504_b : _GEN_21593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21595 = 10'h1f9 == r_count_28_io_out ? io_r_505_b : _GEN_21594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21596 = 10'h1fa == r_count_28_io_out ? io_r_506_b : _GEN_21595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21597 = 10'h1fb == r_count_28_io_out ? io_r_507_b : _GEN_21596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21598 = 10'h1fc == r_count_28_io_out ? io_r_508_b : _GEN_21597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21599 = 10'h1fd == r_count_28_io_out ? io_r_509_b : _GEN_21598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21600 = 10'h1fe == r_count_28_io_out ? io_r_510_b : _GEN_21599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21601 = 10'h1ff == r_count_28_io_out ? io_r_511_b : _GEN_21600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21602 = 10'h200 == r_count_28_io_out ? io_r_512_b : _GEN_21601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21603 = 10'h201 == r_count_28_io_out ? io_r_513_b : _GEN_21602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21604 = 10'h202 == r_count_28_io_out ? io_r_514_b : _GEN_21603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21605 = 10'h203 == r_count_28_io_out ? io_r_515_b : _GEN_21604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21606 = 10'h204 == r_count_28_io_out ? io_r_516_b : _GEN_21605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21607 = 10'h205 == r_count_28_io_out ? io_r_517_b : _GEN_21606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21608 = 10'h206 == r_count_28_io_out ? io_r_518_b : _GEN_21607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21609 = 10'h207 == r_count_28_io_out ? io_r_519_b : _GEN_21608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21610 = 10'h208 == r_count_28_io_out ? io_r_520_b : _GEN_21609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21611 = 10'h209 == r_count_28_io_out ? io_r_521_b : _GEN_21610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21612 = 10'h20a == r_count_28_io_out ? io_r_522_b : _GEN_21611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21613 = 10'h20b == r_count_28_io_out ? io_r_523_b : _GEN_21612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21614 = 10'h20c == r_count_28_io_out ? io_r_524_b : _GEN_21613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21615 = 10'h20d == r_count_28_io_out ? io_r_525_b : _GEN_21614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21616 = 10'h20e == r_count_28_io_out ? io_r_526_b : _GEN_21615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21617 = 10'h20f == r_count_28_io_out ? io_r_527_b : _GEN_21616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21618 = 10'h210 == r_count_28_io_out ? io_r_528_b : _GEN_21617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21619 = 10'h211 == r_count_28_io_out ? io_r_529_b : _GEN_21618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21620 = 10'h212 == r_count_28_io_out ? io_r_530_b : _GEN_21619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21621 = 10'h213 == r_count_28_io_out ? io_r_531_b : _GEN_21620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21622 = 10'h214 == r_count_28_io_out ? io_r_532_b : _GEN_21621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21623 = 10'h215 == r_count_28_io_out ? io_r_533_b : _GEN_21622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21624 = 10'h216 == r_count_28_io_out ? io_r_534_b : _GEN_21623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21625 = 10'h217 == r_count_28_io_out ? io_r_535_b : _GEN_21624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21626 = 10'h218 == r_count_28_io_out ? io_r_536_b : _GEN_21625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21627 = 10'h219 == r_count_28_io_out ? io_r_537_b : _GEN_21626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21628 = 10'h21a == r_count_28_io_out ? io_r_538_b : _GEN_21627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21629 = 10'h21b == r_count_28_io_out ? io_r_539_b : _GEN_21628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21630 = 10'h21c == r_count_28_io_out ? io_r_540_b : _GEN_21629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21631 = 10'h21d == r_count_28_io_out ? io_r_541_b : _GEN_21630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21632 = 10'h21e == r_count_28_io_out ? io_r_542_b : _GEN_21631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21633 = 10'h21f == r_count_28_io_out ? io_r_543_b : _GEN_21632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21634 = 10'h220 == r_count_28_io_out ? io_r_544_b : _GEN_21633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21635 = 10'h221 == r_count_28_io_out ? io_r_545_b : _GEN_21634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21636 = 10'h222 == r_count_28_io_out ? io_r_546_b : _GEN_21635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21637 = 10'h223 == r_count_28_io_out ? io_r_547_b : _GEN_21636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21638 = 10'h224 == r_count_28_io_out ? io_r_548_b : _GEN_21637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21639 = 10'h225 == r_count_28_io_out ? io_r_549_b : _GEN_21638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21640 = 10'h226 == r_count_28_io_out ? io_r_550_b : _GEN_21639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21641 = 10'h227 == r_count_28_io_out ? io_r_551_b : _GEN_21640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21642 = 10'h228 == r_count_28_io_out ? io_r_552_b : _GEN_21641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21643 = 10'h229 == r_count_28_io_out ? io_r_553_b : _GEN_21642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21644 = 10'h22a == r_count_28_io_out ? io_r_554_b : _GEN_21643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21645 = 10'h22b == r_count_28_io_out ? io_r_555_b : _GEN_21644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21646 = 10'h22c == r_count_28_io_out ? io_r_556_b : _GEN_21645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21647 = 10'h22d == r_count_28_io_out ? io_r_557_b : _GEN_21646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21648 = 10'h22e == r_count_28_io_out ? io_r_558_b : _GEN_21647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21649 = 10'h22f == r_count_28_io_out ? io_r_559_b : _GEN_21648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21650 = 10'h230 == r_count_28_io_out ? io_r_560_b : _GEN_21649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21651 = 10'h231 == r_count_28_io_out ? io_r_561_b : _GEN_21650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21652 = 10'h232 == r_count_28_io_out ? io_r_562_b : _GEN_21651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21653 = 10'h233 == r_count_28_io_out ? io_r_563_b : _GEN_21652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21654 = 10'h234 == r_count_28_io_out ? io_r_564_b : _GEN_21653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21655 = 10'h235 == r_count_28_io_out ? io_r_565_b : _GEN_21654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21656 = 10'h236 == r_count_28_io_out ? io_r_566_b : _GEN_21655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21657 = 10'h237 == r_count_28_io_out ? io_r_567_b : _GEN_21656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21658 = 10'h238 == r_count_28_io_out ? io_r_568_b : _GEN_21657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21659 = 10'h239 == r_count_28_io_out ? io_r_569_b : _GEN_21658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21660 = 10'h23a == r_count_28_io_out ? io_r_570_b : _GEN_21659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21661 = 10'h23b == r_count_28_io_out ? io_r_571_b : _GEN_21660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21662 = 10'h23c == r_count_28_io_out ? io_r_572_b : _GEN_21661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21663 = 10'h23d == r_count_28_io_out ? io_r_573_b : _GEN_21662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21664 = 10'h23e == r_count_28_io_out ? io_r_574_b : _GEN_21663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21665 = 10'h23f == r_count_28_io_out ? io_r_575_b : _GEN_21664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21666 = 10'h240 == r_count_28_io_out ? io_r_576_b : _GEN_21665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21667 = 10'h241 == r_count_28_io_out ? io_r_577_b : _GEN_21666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21668 = 10'h242 == r_count_28_io_out ? io_r_578_b : _GEN_21667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21669 = 10'h243 == r_count_28_io_out ? io_r_579_b : _GEN_21668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21670 = 10'h244 == r_count_28_io_out ? io_r_580_b : _GEN_21669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21671 = 10'h245 == r_count_28_io_out ? io_r_581_b : _GEN_21670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21672 = 10'h246 == r_count_28_io_out ? io_r_582_b : _GEN_21671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21673 = 10'h247 == r_count_28_io_out ? io_r_583_b : _GEN_21672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21674 = 10'h248 == r_count_28_io_out ? io_r_584_b : _GEN_21673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21675 = 10'h249 == r_count_28_io_out ? io_r_585_b : _GEN_21674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21676 = 10'h24a == r_count_28_io_out ? io_r_586_b : _GEN_21675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21677 = 10'h24b == r_count_28_io_out ? io_r_587_b : _GEN_21676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21678 = 10'h24c == r_count_28_io_out ? io_r_588_b : _GEN_21677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21679 = 10'h24d == r_count_28_io_out ? io_r_589_b : _GEN_21678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21680 = 10'h24e == r_count_28_io_out ? io_r_590_b : _GEN_21679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21681 = 10'h24f == r_count_28_io_out ? io_r_591_b : _GEN_21680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21682 = 10'h250 == r_count_28_io_out ? io_r_592_b : _GEN_21681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21683 = 10'h251 == r_count_28_io_out ? io_r_593_b : _GEN_21682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21684 = 10'h252 == r_count_28_io_out ? io_r_594_b : _GEN_21683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21685 = 10'h253 == r_count_28_io_out ? io_r_595_b : _GEN_21684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21686 = 10'h254 == r_count_28_io_out ? io_r_596_b : _GEN_21685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21687 = 10'h255 == r_count_28_io_out ? io_r_597_b : _GEN_21686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21688 = 10'h256 == r_count_28_io_out ? io_r_598_b : _GEN_21687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21689 = 10'h257 == r_count_28_io_out ? io_r_599_b : _GEN_21688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21690 = 10'h258 == r_count_28_io_out ? io_r_600_b : _GEN_21689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21691 = 10'h259 == r_count_28_io_out ? io_r_601_b : _GEN_21690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21692 = 10'h25a == r_count_28_io_out ? io_r_602_b : _GEN_21691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21693 = 10'h25b == r_count_28_io_out ? io_r_603_b : _GEN_21692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21694 = 10'h25c == r_count_28_io_out ? io_r_604_b : _GEN_21693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21695 = 10'h25d == r_count_28_io_out ? io_r_605_b : _GEN_21694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21696 = 10'h25e == r_count_28_io_out ? io_r_606_b : _GEN_21695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21697 = 10'h25f == r_count_28_io_out ? io_r_607_b : _GEN_21696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21698 = 10'h260 == r_count_28_io_out ? io_r_608_b : _GEN_21697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21699 = 10'h261 == r_count_28_io_out ? io_r_609_b : _GEN_21698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21700 = 10'h262 == r_count_28_io_out ? io_r_610_b : _GEN_21699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21701 = 10'h263 == r_count_28_io_out ? io_r_611_b : _GEN_21700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21702 = 10'h264 == r_count_28_io_out ? io_r_612_b : _GEN_21701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21703 = 10'h265 == r_count_28_io_out ? io_r_613_b : _GEN_21702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21704 = 10'h266 == r_count_28_io_out ? io_r_614_b : _GEN_21703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21705 = 10'h267 == r_count_28_io_out ? io_r_615_b : _GEN_21704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21706 = 10'h268 == r_count_28_io_out ? io_r_616_b : _GEN_21705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21707 = 10'h269 == r_count_28_io_out ? io_r_617_b : _GEN_21706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21708 = 10'h26a == r_count_28_io_out ? io_r_618_b : _GEN_21707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21709 = 10'h26b == r_count_28_io_out ? io_r_619_b : _GEN_21708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21710 = 10'h26c == r_count_28_io_out ? io_r_620_b : _GEN_21709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21711 = 10'h26d == r_count_28_io_out ? io_r_621_b : _GEN_21710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21712 = 10'h26e == r_count_28_io_out ? io_r_622_b : _GEN_21711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21713 = 10'h26f == r_count_28_io_out ? io_r_623_b : _GEN_21712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21714 = 10'h270 == r_count_28_io_out ? io_r_624_b : _GEN_21713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21715 = 10'h271 == r_count_28_io_out ? io_r_625_b : _GEN_21714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21716 = 10'h272 == r_count_28_io_out ? io_r_626_b : _GEN_21715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21717 = 10'h273 == r_count_28_io_out ? io_r_627_b : _GEN_21716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21718 = 10'h274 == r_count_28_io_out ? io_r_628_b : _GEN_21717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21719 = 10'h275 == r_count_28_io_out ? io_r_629_b : _GEN_21718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21720 = 10'h276 == r_count_28_io_out ? io_r_630_b : _GEN_21719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21721 = 10'h277 == r_count_28_io_out ? io_r_631_b : _GEN_21720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21722 = 10'h278 == r_count_28_io_out ? io_r_632_b : _GEN_21721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21723 = 10'h279 == r_count_28_io_out ? io_r_633_b : _GEN_21722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21724 = 10'h27a == r_count_28_io_out ? io_r_634_b : _GEN_21723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21725 = 10'h27b == r_count_28_io_out ? io_r_635_b : _GEN_21724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21726 = 10'h27c == r_count_28_io_out ? io_r_636_b : _GEN_21725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21727 = 10'h27d == r_count_28_io_out ? io_r_637_b : _GEN_21726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21728 = 10'h27e == r_count_28_io_out ? io_r_638_b : _GEN_21727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21729 = 10'h27f == r_count_28_io_out ? io_r_639_b : _GEN_21728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21730 = 10'h280 == r_count_28_io_out ? io_r_640_b : _GEN_21729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21731 = 10'h281 == r_count_28_io_out ? io_r_641_b : _GEN_21730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21732 = 10'h282 == r_count_28_io_out ? io_r_642_b : _GEN_21731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21733 = 10'h283 == r_count_28_io_out ? io_r_643_b : _GEN_21732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21734 = 10'h284 == r_count_28_io_out ? io_r_644_b : _GEN_21733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21735 = 10'h285 == r_count_28_io_out ? io_r_645_b : _GEN_21734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21736 = 10'h286 == r_count_28_io_out ? io_r_646_b : _GEN_21735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21737 = 10'h287 == r_count_28_io_out ? io_r_647_b : _GEN_21736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21738 = 10'h288 == r_count_28_io_out ? io_r_648_b : _GEN_21737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21739 = 10'h289 == r_count_28_io_out ? io_r_649_b : _GEN_21738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21740 = 10'h28a == r_count_28_io_out ? io_r_650_b : _GEN_21739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21741 = 10'h28b == r_count_28_io_out ? io_r_651_b : _GEN_21740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21742 = 10'h28c == r_count_28_io_out ? io_r_652_b : _GEN_21741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21743 = 10'h28d == r_count_28_io_out ? io_r_653_b : _GEN_21742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21744 = 10'h28e == r_count_28_io_out ? io_r_654_b : _GEN_21743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21745 = 10'h28f == r_count_28_io_out ? io_r_655_b : _GEN_21744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21746 = 10'h290 == r_count_28_io_out ? io_r_656_b : _GEN_21745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21747 = 10'h291 == r_count_28_io_out ? io_r_657_b : _GEN_21746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21748 = 10'h292 == r_count_28_io_out ? io_r_658_b : _GEN_21747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21749 = 10'h293 == r_count_28_io_out ? io_r_659_b : _GEN_21748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21750 = 10'h294 == r_count_28_io_out ? io_r_660_b : _GEN_21749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21751 = 10'h295 == r_count_28_io_out ? io_r_661_b : _GEN_21750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21752 = 10'h296 == r_count_28_io_out ? io_r_662_b : _GEN_21751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21753 = 10'h297 == r_count_28_io_out ? io_r_663_b : _GEN_21752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21754 = 10'h298 == r_count_28_io_out ? io_r_664_b : _GEN_21753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21755 = 10'h299 == r_count_28_io_out ? io_r_665_b : _GEN_21754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21756 = 10'h29a == r_count_28_io_out ? io_r_666_b : _GEN_21755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21757 = 10'h29b == r_count_28_io_out ? io_r_667_b : _GEN_21756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21758 = 10'h29c == r_count_28_io_out ? io_r_668_b : _GEN_21757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21759 = 10'h29d == r_count_28_io_out ? io_r_669_b : _GEN_21758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21760 = 10'h29e == r_count_28_io_out ? io_r_670_b : _GEN_21759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21761 = 10'h29f == r_count_28_io_out ? io_r_671_b : _GEN_21760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21762 = 10'h2a0 == r_count_28_io_out ? io_r_672_b : _GEN_21761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21763 = 10'h2a1 == r_count_28_io_out ? io_r_673_b : _GEN_21762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21764 = 10'h2a2 == r_count_28_io_out ? io_r_674_b : _GEN_21763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21765 = 10'h2a3 == r_count_28_io_out ? io_r_675_b : _GEN_21764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21766 = 10'h2a4 == r_count_28_io_out ? io_r_676_b : _GEN_21765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21767 = 10'h2a5 == r_count_28_io_out ? io_r_677_b : _GEN_21766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21768 = 10'h2a6 == r_count_28_io_out ? io_r_678_b : _GEN_21767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21769 = 10'h2a7 == r_count_28_io_out ? io_r_679_b : _GEN_21768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21770 = 10'h2a8 == r_count_28_io_out ? io_r_680_b : _GEN_21769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21771 = 10'h2a9 == r_count_28_io_out ? io_r_681_b : _GEN_21770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21772 = 10'h2aa == r_count_28_io_out ? io_r_682_b : _GEN_21771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21773 = 10'h2ab == r_count_28_io_out ? io_r_683_b : _GEN_21772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21774 = 10'h2ac == r_count_28_io_out ? io_r_684_b : _GEN_21773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21775 = 10'h2ad == r_count_28_io_out ? io_r_685_b : _GEN_21774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21776 = 10'h2ae == r_count_28_io_out ? io_r_686_b : _GEN_21775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21777 = 10'h2af == r_count_28_io_out ? io_r_687_b : _GEN_21776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21778 = 10'h2b0 == r_count_28_io_out ? io_r_688_b : _GEN_21777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21779 = 10'h2b1 == r_count_28_io_out ? io_r_689_b : _GEN_21778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21780 = 10'h2b2 == r_count_28_io_out ? io_r_690_b : _GEN_21779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21781 = 10'h2b3 == r_count_28_io_out ? io_r_691_b : _GEN_21780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21782 = 10'h2b4 == r_count_28_io_out ? io_r_692_b : _GEN_21781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21783 = 10'h2b5 == r_count_28_io_out ? io_r_693_b : _GEN_21782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21784 = 10'h2b6 == r_count_28_io_out ? io_r_694_b : _GEN_21783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21785 = 10'h2b7 == r_count_28_io_out ? io_r_695_b : _GEN_21784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21786 = 10'h2b8 == r_count_28_io_out ? io_r_696_b : _GEN_21785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21787 = 10'h2b9 == r_count_28_io_out ? io_r_697_b : _GEN_21786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21788 = 10'h2ba == r_count_28_io_out ? io_r_698_b : _GEN_21787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21789 = 10'h2bb == r_count_28_io_out ? io_r_699_b : _GEN_21788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21790 = 10'h2bc == r_count_28_io_out ? io_r_700_b : _GEN_21789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21791 = 10'h2bd == r_count_28_io_out ? io_r_701_b : _GEN_21790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21792 = 10'h2be == r_count_28_io_out ? io_r_702_b : _GEN_21791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21793 = 10'h2bf == r_count_28_io_out ? io_r_703_b : _GEN_21792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21794 = 10'h2c0 == r_count_28_io_out ? io_r_704_b : _GEN_21793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21795 = 10'h2c1 == r_count_28_io_out ? io_r_705_b : _GEN_21794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21796 = 10'h2c2 == r_count_28_io_out ? io_r_706_b : _GEN_21795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21797 = 10'h2c3 == r_count_28_io_out ? io_r_707_b : _GEN_21796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21798 = 10'h2c4 == r_count_28_io_out ? io_r_708_b : _GEN_21797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21799 = 10'h2c5 == r_count_28_io_out ? io_r_709_b : _GEN_21798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21800 = 10'h2c6 == r_count_28_io_out ? io_r_710_b : _GEN_21799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21801 = 10'h2c7 == r_count_28_io_out ? io_r_711_b : _GEN_21800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21802 = 10'h2c8 == r_count_28_io_out ? io_r_712_b : _GEN_21801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21803 = 10'h2c9 == r_count_28_io_out ? io_r_713_b : _GEN_21802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21804 = 10'h2ca == r_count_28_io_out ? io_r_714_b : _GEN_21803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21805 = 10'h2cb == r_count_28_io_out ? io_r_715_b : _GEN_21804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21806 = 10'h2cc == r_count_28_io_out ? io_r_716_b : _GEN_21805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21807 = 10'h2cd == r_count_28_io_out ? io_r_717_b : _GEN_21806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21808 = 10'h2ce == r_count_28_io_out ? io_r_718_b : _GEN_21807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21809 = 10'h2cf == r_count_28_io_out ? io_r_719_b : _GEN_21808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21810 = 10'h2d0 == r_count_28_io_out ? io_r_720_b : _GEN_21809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21811 = 10'h2d1 == r_count_28_io_out ? io_r_721_b : _GEN_21810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21812 = 10'h2d2 == r_count_28_io_out ? io_r_722_b : _GEN_21811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21813 = 10'h2d3 == r_count_28_io_out ? io_r_723_b : _GEN_21812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21814 = 10'h2d4 == r_count_28_io_out ? io_r_724_b : _GEN_21813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21815 = 10'h2d5 == r_count_28_io_out ? io_r_725_b : _GEN_21814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21816 = 10'h2d6 == r_count_28_io_out ? io_r_726_b : _GEN_21815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21817 = 10'h2d7 == r_count_28_io_out ? io_r_727_b : _GEN_21816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21818 = 10'h2d8 == r_count_28_io_out ? io_r_728_b : _GEN_21817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21819 = 10'h2d9 == r_count_28_io_out ? io_r_729_b : _GEN_21818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21820 = 10'h2da == r_count_28_io_out ? io_r_730_b : _GEN_21819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21821 = 10'h2db == r_count_28_io_out ? io_r_731_b : _GEN_21820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21822 = 10'h2dc == r_count_28_io_out ? io_r_732_b : _GEN_21821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21823 = 10'h2dd == r_count_28_io_out ? io_r_733_b : _GEN_21822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21824 = 10'h2de == r_count_28_io_out ? io_r_734_b : _GEN_21823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21825 = 10'h2df == r_count_28_io_out ? io_r_735_b : _GEN_21824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21826 = 10'h2e0 == r_count_28_io_out ? io_r_736_b : _GEN_21825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21827 = 10'h2e1 == r_count_28_io_out ? io_r_737_b : _GEN_21826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21828 = 10'h2e2 == r_count_28_io_out ? io_r_738_b : _GEN_21827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21829 = 10'h2e3 == r_count_28_io_out ? io_r_739_b : _GEN_21828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21830 = 10'h2e4 == r_count_28_io_out ? io_r_740_b : _GEN_21829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21831 = 10'h2e5 == r_count_28_io_out ? io_r_741_b : _GEN_21830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21832 = 10'h2e6 == r_count_28_io_out ? io_r_742_b : _GEN_21831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21833 = 10'h2e7 == r_count_28_io_out ? io_r_743_b : _GEN_21832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21834 = 10'h2e8 == r_count_28_io_out ? io_r_744_b : _GEN_21833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21835 = 10'h2e9 == r_count_28_io_out ? io_r_745_b : _GEN_21834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21836 = 10'h2ea == r_count_28_io_out ? io_r_746_b : _GEN_21835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21837 = 10'h2eb == r_count_28_io_out ? io_r_747_b : _GEN_21836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21838 = 10'h2ec == r_count_28_io_out ? io_r_748_b : _GEN_21837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21841 = 10'h1 == r_count_29_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21842 = 10'h2 == r_count_29_io_out ? io_r_2_b : _GEN_21841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21843 = 10'h3 == r_count_29_io_out ? io_r_3_b : _GEN_21842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21844 = 10'h4 == r_count_29_io_out ? io_r_4_b : _GEN_21843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21845 = 10'h5 == r_count_29_io_out ? io_r_5_b : _GEN_21844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21846 = 10'h6 == r_count_29_io_out ? io_r_6_b : _GEN_21845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21847 = 10'h7 == r_count_29_io_out ? io_r_7_b : _GEN_21846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21848 = 10'h8 == r_count_29_io_out ? io_r_8_b : _GEN_21847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21849 = 10'h9 == r_count_29_io_out ? io_r_9_b : _GEN_21848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21850 = 10'ha == r_count_29_io_out ? io_r_10_b : _GEN_21849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21851 = 10'hb == r_count_29_io_out ? io_r_11_b : _GEN_21850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21852 = 10'hc == r_count_29_io_out ? io_r_12_b : _GEN_21851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21853 = 10'hd == r_count_29_io_out ? io_r_13_b : _GEN_21852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21854 = 10'he == r_count_29_io_out ? io_r_14_b : _GEN_21853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21855 = 10'hf == r_count_29_io_out ? io_r_15_b : _GEN_21854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21856 = 10'h10 == r_count_29_io_out ? io_r_16_b : _GEN_21855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21857 = 10'h11 == r_count_29_io_out ? io_r_17_b : _GEN_21856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21858 = 10'h12 == r_count_29_io_out ? io_r_18_b : _GEN_21857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21859 = 10'h13 == r_count_29_io_out ? io_r_19_b : _GEN_21858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21860 = 10'h14 == r_count_29_io_out ? io_r_20_b : _GEN_21859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21861 = 10'h15 == r_count_29_io_out ? io_r_21_b : _GEN_21860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21862 = 10'h16 == r_count_29_io_out ? io_r_22_b : _GEN_21861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21863 = 10'h17 == r_count_29_io_out ? io_r_23_b : _GEN_21862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21864 = 10'h18 == r_count_29_io_out ? io_r_24_b : _GEN_21863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21865 = 10'h19 == r_count_29_io_out ? io_r_25_b : _GEN_21864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21866 = 10'h1a == r_count_29_io_out ? io_r_26_b : _GEN_21865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21867 = 10'h1b == r_count_29_io_out ? io_r_27_b : _GEN_21866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21868 = 10'h1c == r_count_29_io_out ? io_r_28_b : _GEN_21867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21869 = 10'h1d == r_count_29_io_out ? io_r_29_b : _GEN_21868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21870 = 10'h1e == r_count_29_io_out ? io_r_30_b : _GEN_21869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21871 = 10'h1f == r_count_29_io_out ? io_r_31_b : _GEN_21870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21872 = 10'h20 == r_count_29_io_out ? io_r_32_b : _GEN_21871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21873 = 10'h21 == r_count_29_io_out ? io_r_33_b : _GEN_21872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21874 = 10'h22 == r_count_29_io_out ? io_r_34_b : _GEN_21873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21875 = 10'h23 == r_count_29_io_out ? io_r_35_b : _GEN_21874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21876 = 10'h24 == r_count_29_io_out ? io_r_36_b : _GEN_21875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21877 = 10'h25 == r_count_29_io_out ? io_r_37_b : _GEN_21876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21878 = 10'h26 == r_count_29_io_out ? io_r_38_b : _GEN_21877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21879 = 10'h27 == r_count_29_io_out ? io_r_39_b : _GEN_21878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21880 = 10'h28 == r_count_29_io_out ? io_r_40_b : _GEN_21879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21881 = 10'h29 == r_count_29_io_out ? io_r_41_b : _GEN_21880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21882 = 10'h2a == r_count_29_io_out ? io_r_42_b : _GEN_21881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21883 = 10'h2b == r_count_29_io_out ? io_r_43_b : _GEN_21882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21884 = 10'h2c == r_count_29_io_out ? io_r_44_b : _GEN_21883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21885 = 10'h2d == r_count_29_io_out ? io_r_45_b : _GEN_21884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21886 = 10'h2e == r_count_29_io_out ? io_r_46_b : _GEN_21885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21887 = 10'h2f == r_count_29_io_out ? io_r_47_b : _GEN_21886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21888 = 10'h30 == r_count_29_io_out ? io_r_48_b : _GEN_21887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21889 = 10'h31 == r_count_29_io_out ? io_r_49_b : _GEN_21888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21890 = 10'h32 == r_count_29_io_out ? io_r_50_b : _GEN_21889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21891 = 10'h33 == r_count_29_io_out ? io_r_51_b : _GEN_21890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21892 = 10'h34 == r_count_29_io_out ? io_r_52_b : _GEN_21891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21893 = 10'h35 == r_count_29_io_out ? io_r_53_b : _GEN_21892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21894 = 10'h36 == r_count_29_io_out ? io_r_54_b : _GEN_21893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21895 = 10'h37 == r_count_29_io_out ? io_r_55_b : _GEN_21894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21896 = 10'h38 == r_count_29_io_out ? io_r_56_b : _GEN_21895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21897 = 10'h39 == r_count_29_io_out ? io_r_57_b : _GEN_21896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21898 = 10'h3a == r_count_29_io_out ? io_r_58_b : _GEN_21897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21899 = 10'h3b == r_count_29_io_out ? io_r_59_b : _GEN_21898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21900 = 10'h3c == r_count_29_io_out ? io_r_60_b : _GEN_21899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21901 = 10'h3d == r_count_29_io_out ? io_r_61_b : _GEN_21900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21902 = 10'h3e == r_count_29_io_out ? io_r_62_b : _GEN_21901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21903 = 10'h3f == r_count_29_io_out ? io_r_63_b : _GEN_21902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21904 = 10'h40 == r_count_29_io_out ? io_r_64_b : _GEN_21903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21905 = 10'h41 == r_count_29_io_out ? io_r_65_b : _GEN_21904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21906 = 10'h42 == r_count_29_io_out ? io_r_66_b : _GEN_21905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21907 = 10'h43 == r_count_29_io_out ? io_r_67_b : _GEN_21906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21908 = 10'h44 == r_count_29_io_out ? io_r_68_b : _GEN_21907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21909 = 10'h45 == r_count_29_io_out ? io_r_69_b : _GEN_21908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21910 = 10'h46 == r_count_29_io_out ? io_r_70_b : _GEN_21909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21911 = 10'h47 == r_count_29_io_out ? io_r_71_b : _GEN_21910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21912 = 10'h48 == r_count_29_io_out ? io_r_72_b : _GEN_21911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21913 = 10'h49 == r_count_29_io_out ? io_r_73_b : _GEN_21912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21914 = 10'h4a == r_count_29_io_out ? io_r_74_b : _GEN_21913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21915 = 10'h4b == r_count_29_io_out ? io_r_75_b : _GEN_21914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21916 = 10'h4c == r_count_29_io_out ? io_r_76_b : _GEN_21915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21917 = 10'h4d == r_count_29_io_out ? io_r_77_b : _GEN_21916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21918 = 10'h4e == r_count_29_io_out ? io_r_78_b : _GEN_21917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21919 = 10'h4f == r_count_29_io_out ? io_r_79_b : _GEN_21918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21920 = 10'h50 == r_count_29_io_out ? io_r_80_b : _GEN_21919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21921 = 10'h51 == r_count_29_io_out ? io_r_81_b : _GEN_21920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21922 = 10'h52 == r_count_29_io_out ? io_r_82_b : _GEN_21921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21923 = 10'h53 == r_count_29_io_out ? io_r_83_b : _GEN_21922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21924 = 10'h54 == r_count_29_io_out ? io_r_84_b : _GEN_21923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21925 = 10'h55 == r_count_29_io_out ? io_r_85_b : _GEN_21924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21926 = 10'h56 == r_count_29_io_out ? io_r_86_b : _GEN_21925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21927 = 10'h57 == r_count_29_io_out ? io_r_87_b : _GEN_21926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21928 = 10'h58 == r_count_29_io_out ? io_r_88_b : _GEN_21927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21929 = 10'h59 == r_count_29_io_out ? io_r_89_b : _GEN_21928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21930 = 10'h5a == r_count_29_io_out ? io_r_90_b : _GEN_21929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21931 = 10'h5b == r_count_29_io_out ? io_r_91_b : _GEN_21930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21932 = 10'h5c == r_count_29_io_out ? io_r_92_b : _GEN_21931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21933 = 10'h5d == r_count_29_io_out ? io_r_93_b : _GEN_21932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21934 = 10'h5e == r_count_29_io_out ? io_r_94_b : _GEN_21933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21935 = 10'h5f == r_count_29_io_out ? io_r_95_b : _GEN_21934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21936 = 10'h60 == r_count_29_io_out ? io_r_96_b : _GEN_21935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21937 = 10'h61 == r_count_29_io_out ? io_r_97_b : _GEN_21936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21938 = 10'h62 == r_count_29_io_out ? io_r_98_b : _GEN_21937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21939 = 10'h63 == r_count_29_io_out ? io_r_99_b : _GEN_21938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21940 = 10'h64 == r_count_29_io_out ? io_r_100_b : _GEN_21939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21941 = 10'h65 == r_count_29_io_out ? io_r_101_b : _GEN_21940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21942 = 10'h66 == r_count_29_io_out ? io_r_102_b : _GEN_21941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21943 = 10'h67 == r_count_29_io_out ? io_r_103_b : _GEN_21942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21944 = 10'h68 == r_count_29_io_out ? io_r_104_b : _GEN_21943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21945 = 10'h69 == r_count_29_io_out ? io_r_105_b : _GEN_21944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21946 = 10'h6a == r_count_29_io_out ? io_r_106_b : _GEN_21945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21947 = 10'h6b == r_count_29_io_out ? io_r_107_b : _GEN_21946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21948 = 10'h6c == r_count_29_io_out ? io_r_108_b : _GEN_21947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21949 = 10'h6d == r_count_29_io_out ? io_r_109_b : _GEN_21948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21950 = 10'h6e == r_count_29_io_out ? io_r_110_b : _GEN_21949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21951 = 10'h6f == r_count_29_io_out ? io_r_111_b : _GEN_21950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21952 = 10'h70 == r_count_29_io_out ? io_r_112_b : _GEN_21951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21953 = 10'h71 == r_count_29_io_out ? io_r_113_b : _GEN_21952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21954 = 10'h72 == r_count_29_io_out ? io_r_114_b : _GEN_21953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21955 = 10'h73 == r_count_29_io_out ? io_r_115_b : _GEN_21954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21956 = 10'h74 == r_count_29_io_out ? io_r_116_b : _GEN_21955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21957 = 10'h75 == r_count_29_io_out ? io_r_117_b : _GEN_21956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21958 = 10'h76 == r_count_29_io_out ? io_r_118_b : _GEN_21957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21959 = 10'h77 == r_count_29_io_out ? io_r_119_b : _GEN_21958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21960 = 10'h78 == r_count_29_io_out ? io_r_120_b : _GEN_21959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21961 = 10'h79 == r_count_29_io_out ? io_r_121_b : _GEN_21960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21962 = 10'h7a == r_count_29_io_out ? io_r_122_b : _GEN_21961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21963 = 10'h7b == r_count_29_io_out ? io_r_123_b : _GEN_21962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21964 = 10'h7c == r_count_29_io_out ? io_r_124_b : _GEN_21963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21965 = 10'h7d == r_count_29_io_out ? io_r_125_b : _GEN_21964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21966 = 10'h7e == r_count_29_io_out ? io_r_126_b : _GEN_21965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21967 = 10'h7f == r_count_29_io_out ? io_r_127_b : _GEN_21966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21968 = 10'h80 == r_count_29_io_out ? io_r_128_b : _GEN_21967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21969 = 10'h81 == r_count_29_io_out ? io_r_129_b : _GEN_21968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21970 = 10'h82 == r_count_29_io_out ? io_r_130_b : _GEN_21969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21971 = 10'h83 == r_count_29_io_out ? io_r_131_b : _GEN_21970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21972 = 10'h84 == r_count_29_io_out ? io_r_132_b : _GEN_21971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21973 = 10'h85 == r_count_29_io_out ? io_r_133_b : _GEN_21972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21974 = 10'h86 == r_count_29_io_out ? io_r_134_b : _GEN_21973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21975 = 10'h87 == r_count_29_io_out ? io_r_135_b : _GEN_21974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21976 = 10'h88 == r_count_29_io_out ? io_r_136_b : _GEN_21975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21977 = 10'h89 == r_count_29_io_out ? io_r_137_b : _GEN_21976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21978 = 10'h8a == r_count_29_io_out ? io_r_138_b : _GEN_21977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21979 = 10'h8b == r_count_29_io_out ? io_r_139_b : _GEN_21978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21980 = 10'h8c == r_count_29_io_out ? io_r_140_b : _GEN_21979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21981 = 10'h8d == r_count_29_io_out ? io_r_141_b : _GEN_21980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21982 = 10'h8e == r_count_29_io_out ? io_r_142_b : _GEN_21981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21983 = 10'h8f == r_count_29_io_out ? io_r_143_b : _GEN_21982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21984 = 10'h90 == r_count_29_io_out ? io_r_144_b : _GEN_21983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21985 = 10'h91 == r_count_29_io_out ? io_r_145_b : _GEN_21984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21986 = 10'h92 == r_count_29_io_out ? io_r_146_b : _GEN_21985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21987 = 10'h93 == r_count_29_io_out ? io_r_147_b : _GEN_21986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21988 = 10'h94 == r_count_29_io_out ? io_r_148_b : _GEN_21987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21989 = 10'h95 == r_count_29_io_out ? io_r_149_b : _GEN_21988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21990 = 10'h96 == r_count_29_io_out ? io_r_150_b : _GEN_21989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21991 = 10'h97 == r_count_29_io_out ? io_r_151_b : _GEN_21990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21992 = 10'h98 == r_count_29_io_out ? io_r_152_b : _GEN_21991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21993 = 10'h99 == r_count_29_io_out ? io_r_153_b : _GEN_21992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21994 = 10'h9a == r_count_29_io_out ? io_r_154_b : _GEN_21993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21995 = 10'h9b == r_count_29_io_out ? io_r_155_b : _GEN_21994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21996 = 10'h9c == r_count_29_io_out ? io_r_156_b : _GEN_21995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21997 = 10'h9d == r_count_29_io_out ? io_r_157_b : _GEN_21996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21998 = 10'h9e == r_count_29_io_out ? io_r_158_b : _GEN_21997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_21999 = 10'h9f == r_count_29_io_out ? io_r_159_b : _GEN_21998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22000 = 10'ha0 == r_count_29_io_out ? io_r_160_b : _GEN_21999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22001 = 10'ha1 == r_count_29_io_out ? io_r_161_b : _GEN_22000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22002 = 10'ha2 == r_count_29_io_out ? io_r_162_b : _GEN_22001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22003 = 10'ha3 == r_count_29_io_out ? io_r_163_b : _GEN_22002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22004 = 10'ha4 == r_count_29_io_out ? io_r_164_b : _GEN_22003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22005 = 10'ha5 == r_count_29_io_out ? io_r_165_b : _GEN_22004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22006 = 10'ha6 == r_count_29_io_out ? io_r_166_b : _GEN_22005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22007 = 10'ha7 == r_count_29_io_out ? io_r_167_b : _GEN_22006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22008 = 10'ha8 == r_count_29_io_out ? io_r_168_b : _GEN_22007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22009 = 10'ha9 == r_count_29_io_out ? io_r_169_b : _GEN_22008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22010 = 10'haa == r_count_29_io_out ? io_r_170_b : _GEN_22009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22011 = 10'hab == r_count_29_io_out ? io_r_171_b : _GEN_22010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22012 = 10'hac == r_count_29_io_out ? io_r_172_b : _GEN_22011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22013 = 10'had == r_count_29_io_out ? io_r_173_b : _GEN_22012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22014 = 10'hae == r_count_29_io_out ? io_r_174_b : _GEN_22013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22015 = 10'haf == r_count_29_io_out ? io_r_175_b : _GEN_22014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22016 = 10'hb0 == r_count_29_io_out ? io_r_176_b : _GEN_22015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22017 = 10'hb1 == r_count_29_io_out ? io_r_177_b : _GEN_22016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22018 = 10'hb2 == r_count_29_io_out ? io_r_178_b : _GEN_22017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22019 = 10'hb3 == r_count_29_io_out ? io_r_179_b : _GEN_22018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22020 = 10'hb4 == r_count_29_io_out ? io_r_180_b : _GEN_22019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22021 = 10'hb5 == r_count_29_io_out ? io_r_181_b : _GEN_22020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22022 = 10'hb6 == r_count_29_io_out ? io_r_182_b : _GEN_22021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22023 = 10'hb7 == r_count_29_io_out ? io_r_183_b : _GEN_22022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22024 = 10'hb8 == r_count_29_io_out ? io_r_184_b : _GEN_22023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22025 = 10'hb9 == r_count_29_io_out ? io_r_185_b : _GEN_22024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22026 = 10'hba == r_count_29_io_out ? io_r_186_b : _GEN_22025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22027 = 10'hbb == r_count_29_io_out ? io_r_187_b : _GEN_22026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22028 = 10'hbc == r_count_29_io_out ? io_r_188_b : _GEN_22027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22029 = 10'hbd == r_count_29_io_out ? io_r_189_b : _GEN_22028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22030 = 10'hbe == r_count_29_io_out ? io_r_190_b : _GEN_22029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22031 = 10'hbf == r_count_29_io_out ? io_r_191_b : _GEN_22030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22032 = 10'hc0 == r_count_29_io_out ? io_r_192_b : _GEN_22031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22033 = 10'hc1 == r_count_29_io_out ? io_r_193_b : _GEN_22032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22034 = 10'hc2 == r_count_29_io_out ? io_r_194_b : _GEN_22033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22035 = 10'hc3 == r_count_29_io_out ? io_r_195_b : _GEN_22034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22036 = 10'hc4 == r_count_29_io_out ? io_r_196_b : _GEN_22035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22037 = 10'hc5 == r_count_29_io_out ? io_r_197_b : _GEN_22036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22038 = 10'hc6 == r_count_29_io_out ? io_r_198_b : _GEN_22037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22039 = 10'hc7 == r_count_29_io_out ? io_r_199_b : _GEN_22038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22040 = 10'hc8 == r_count_29_io_out ? io_r_200_b : _GEN_22039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22041 = 10'hc9 == r_count_29_io_out ? io_r_201_b : _GEN_22040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22042 = 10'hca == r_count_29_io_out ? io_r_202_b : _GEN_22041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22043 = 10'hcb == r_count_29_io_out ? io_r_203_b : _GEN_22042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22044 = 10'hcc == r_count_29_io_out ? io_r_204_b : _GEN_22043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22045 = 10'hcd == r_count_29_io_out ? io_r_205_b : _GEN_22044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22046 = 10'hce == r_count_29_io_out ? io_r_206_b : _GEN_22045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22047 = 10'hcf == r_count_29_io_out ? io_r_207_b : _GEN_22046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22048 = 10'hd0 == r_count_29_io_out ? io_r_208_b : _GEN_22047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22049 = 10'hd1 == r_count_29_io_out ? io_r_209_b : _GEN_22048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22050 = 10'hd2 == r_count_29_io_out ? io_r_210_b : _GEN_22049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22051 = 10'hd3 == r_count_29_io_out ? io_r_211_b : _GEN_22050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22052 = 10'hd4 == r_count_29_io_out ? io_r_212_b : _GEN_22051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22053 = 10'hd5 == r_count_29_io_out ? io_r_213_b : _GEN_22052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22054 = 10'hd6 == r_count_29_io_out ? io_r_214_b : _GEN_22053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22055 = 10'hd7 == r_count_29_io_out ? io_r_215_b : _GEN_22054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22056 = 10'hd8 == r_count_29_io_out ? io_r_216_b : _GEN_22055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22057 = 10'hd9 == r_count_29_io_out ? io_r_217_b : _GEN_22056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22058 = 10'hda == r_count_29_io_out ? io_r_218_b : _GEN_22057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22059 = 10'hdb == r_count_29_io_out ? io_r_219_b : _GEN_22058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22060 = 10'hdc == r_count_29_io_out ? io_r_220_b : _GEN_22059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22061 = 10'hdd == r_count_29_io_out ? io_r_221_b : _GEN_22060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22062 = 10'hde == r_count_29_io_out ? io_r_222_b : _GEN_22061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22063 = 10'hdf == r_count_29_io_out ? io_r_223_b : _GEN_22062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22064 = 10'he0 == r_count_29_io_out ? io_r_224_b : _GEN_22063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22065 = 10'he1 == r_count_29_io_out ? io_r_225_b : _GEN_22064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22066 = 10'he2 == r_count_29_io_out ? io_r_226_b : _GEN_22065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22067 = 10'he3 == r_count_29_io_out ? io_r_227_b : _GEN_22066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22068 = 10'he4 == r_count_29_io_out ? io_r_228_b : _GEN_22067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22069 = 10'he5 == r_count_29_io_out ? io_r_229_b : _GEN_22068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22070 = 10'he6 == r_count_29_io_out ? io_r_230_b : _GEN_22069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22071 = 10'he7 == r_count_29_io_out ? io_r_231_b : _GEN_22070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22072 = 10'he8 == r_count_29_io_out ? io_r_232_b : _GEN_22071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22073 = 10'he9 == r_count_29_io_out ? io_r_233_b : _GEN_22072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22074 = 10'hea == r_count_29_io_out ? io_r_234_b : _GEN_22073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22075 = 10'heb == r_count_29_io_out ? io_r_235_b : _GEN_22074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22076 = 10'hec == r_count_29_io_out ? io_r_236_b : _GEN_22075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22077 = 10'hed == r_count_29_io_out ? io_r_237_b : _GEN_22076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22078 = 10'hee == r_count_29_io_out ? io_r_238_b : _GEN_22077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22079 = 10'hef == r_count_29_io_out ? io_r_239_b : _GEN_22078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22080 = 10'hf0 == r_count_29_io_out ? io_r_240_b : _GEN_22079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22081 = 10'hf1 == r_count_29_io_out ? io_r_241_b : _GEN_22080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22082 = 10'hf2 == r_count_29_io_out ? io_r_242_b : _GEN_22081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22083 = 10'hf3 == r_count_29_io_out ? io_r_243_b : _GEN_22082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22084 = 10'hf4 == r_count_29_io_out ? io_r_244_b : _GEN_22083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22085 = 10'hf5 == r_count_29_io_out ? io_r_245_b : _GEN_22084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22086 = 10'hf6 == r_count_29_io_out ? io_r_246_b : _GEN_22085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22087 = 10'hf7 == r_count_29_io_out ? io_r_247_b : _GEN_22086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22088 = 10'hf8 == r_count_29_io_out ? io_r_248_b : _GEN_22087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22089 = 10'hf9 == r_count_29_io_out ? io_r_249_b : _GEN_22088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22090 = 10'hfa == r_count_29_io_out ? io_r_250_b : _GEN_22089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22091 = 10'hfb == r_count_29_io_out ? io_r_251_b : _GEN_22090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22092 = 10'hfc == r_count_29_io_out ? io_r_252_b : _GEN_22091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22093 = 10'hfd == r_count_29_io_out ? io_r_253_b : _GEN_22092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22094 = 10'hfe == r_count_29_io_out ? io_r_254_b : _GEN_22093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22095 = 10'hff == r_count_29_io_out ? io_r_255_b : _GEN_22094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22096 = 10'h100 == r_count_29_io_out ? io_r_256_b : _GEN_22095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22097 = 10'h101 == r_count_29_io_out ? io_r_257_b : _GEN_22096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22098 = 10'h102 == r_count_29_io_out ? io_r_258_b : _GEN_22097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22099 = 10'h103 == r_count_29_io_out ? io_r_259_b : _GEN_22098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22100 = 10'h104 == r_count_29_io_out ? io_r_260_b : _GEN_22099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22101 = 10'h105 == r_count_29_io_out ? io_r_261_b : _GEN_22100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22102 = 10'h106 == r_count_29_io_out ? io_r_262_b : _GEN_22101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22103 = 10'h107 == r_count_29_io_out ? io_r_263_b : _GEN_22102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22104 = 10'h108 == r_count_29_io_out ? io_r_264_b : _GEN_22103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22105 = 10'h109 == r_count_29_io_out ? io_r_265_b : _GEN_22104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22106 = 10'h10a == r_count_29_io_out ? io_r_266_b : _GEN_22105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22107 = 10'h10b == r_count_29_io_out ? io_r_267_b : _GEN_22106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22108 = 10'h10c == r_count_29_io_out ? io_r_268_b : _GEN_22107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22109 = 10'h10d == r_count_29_io_out ? io_r_269_b : _GEN_22108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22110 = 10'h10e == r_count_29_io_out ? io_r_270_b : _GEN_22109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22111 = 10'h10f == r_count_29_io_out ? io_r_271_b : _GEN_22110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22112 = 10'h110 == r_count_29_io_out ? io_r_272_b : _GEN_22111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22113 = 10'h111 == r_count_29_io_out ? io_r_273_b : _GEN_22112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22114 = 10'h112 == r_count_29_io_out ? io_r_274_b : _GEN_22113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22115 = 10'h113 == r_count_29_io_out ? io_r_275_b : _GEN_22114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22116 = 10'h114 == r_count_29_io_out ? io_r_276_b : _GEN_22115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22117 = 10'h115 == r_count_29_io_out ? io_r_277_b : _GEN_22116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22118 = 10'h116 == r_count_29_io_out ? io_r_278_b : _GEN_22117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22119 = 10'h117 == r_count_29_io_out ? io_r_279_b : _GEN_22118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22120 = 10'h118 == r_count_29_io_out ? io_r_280_b : _GEN_22119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22121 = 10'h119 == r_count_29_io_out ? io_r_281_b : _GEN_22120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22122 = 10'h11a == r_count_29_io_out ? io_r_282_b : _GEN_22121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22123 = 10'h11b == r_count_29_io_out ? io_r_283_b : _GEN_22122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22124 = 10'h11c == r_count_29_io_out ? io_r_284_b : _GEN_22123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22125 = 10'h11d == r_count_29_io_out ? io_r_285_b : _GEN_22124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22126 = 10'h11e == r_count_29_io_out ? io_r_286_b : _GEN_22125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22127 = 10'h11f == r_count_29_io_out ? io_r_287_b : _GEN_22126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22128 = 10'h120 == r_count_29_io_out ? io_r_288_b : _GEN_22127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22129 = 10'h121 == r_count_29_io_out ? io_r_289_b : _GEN_22128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22130 = 10'h122 == r_count_29_io_out ? io_r_290_b : _GEN_22129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22131 = 10'h123 == r_count_29_io_out ? io_r_291_b : _GEN_22130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22132 = 10'h124 == r_count_29_io_out ? io_r_292_b : _GEN_22131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22133 = 10'h125 == r_count_29_io_out ? io_r_293_b : _GEN_22132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22134 = 10'h126 == r_count_29_io_out ? io_r_294_b : _GEN_22133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22135 = 10'h127 == r_count_29_io_out ? io_r_295_b : _GEN_22134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22136 = 10'h128 == r_count_29_io_out ? io_r_296_b : _GEN_22135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22137 = 10'h129 == r_count_29_io_out ? io_r_297_b : _GEN_22136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22138 = 10'h12a == r_count_29_io_out ? io_r_298_b : _GEN_22137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22139 = 10'h12b == r_count_29_io_out ? io_r_299_b : _GEN_22138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22140 = 10'h12c == r_count_29_io_out ? io_r_300_b : _GEN_22139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22141 = 10'h12d == r_count_29_io_out ? io_r_301_b : _GEN_22140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22142 = 10'h12e == r_count_29_io_out ? io_r_302_b : _GEN_22141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22143 = 10'h12f == r_count_29_io_out ? io_r_303_b : _GEN_22142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22144 = 10'h130 == r_count_29_io_out ? io_r_304_b : _GEN_22143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22145 = 10'h131 == r_count_29_io_out ? io_r_305_b : _GEN_22144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22146 = 10'h132 == r_count_29_io_out ? io_r_306_b : _GEN_22145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22147 = 10'h133 == r_count_29_io_out ? io_r_307_b : _GEN_22146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22148 = 10'h134 == r_count_29_io_out ? io_r_308_b : _GEN_22147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22149 = 10'h135 == r_count_29_io_out ? io_r_309_b : _GEN_22148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22150 = 10'h136 == r_count_29_io_out ? io_r_310_b : _GEN_22149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22151 = 10'h137 == r_count_29_io_out ? io_r_311_b : _GEN_22150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22152 = 10'h138 == r_count_29_io_out ? io_r_312_b : _GEN_22151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22153 = 10'h139 == r_count_29_io_out ? io_r_313_b : _GEN_22152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22154 = 10'h13a == r_count_29_io_out ? io_r_314_b : _GEN_22153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22155 = 10'h13b == r_count_29_io_out ? io_r_315_b : _GEN_22154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22156 = 10'h13c == r_count_29_io_out ? io_r_316_b : _GEN_22155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22157 = 10'h13d == r_count_29_io_out ? io_r_317_b : _GEN_22156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22158 = 10'h13e == r_count_29_io_out ? io_r_318_b : _GEN_22157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22159 = 10'h13f == r_count_29_io_out ? io_r_319_b : _GEN_22158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22160 = 10'h140 == r_count_29_io_out ? io_r_320_b : _GEN_22159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22161 = 10'h141 == r_count_29_io_out ? io_r_321_b : _GEN_22160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22162 = 10'h142 == r_count_29_io_out ? io_r_322_b : _GEN_22161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22163 = 10'h143 == r_count_29_io_out ? io_r_323_b : _GEN_22162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22164 = 10'h144 == r_count_29_io_out ? io_r_324_b : _GEN_22163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22165 = 10'h145 == r_count_29_io_out ? io_r_325_b : _GEN_22164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22166 = 10'h146 == r_count_29_io_out ? io_r_326_b : _GEN_22165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22167 = 10'h147 == r_count_29_io_out ? io_r_327_b : _GEN_22166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22168 = 10'h148 == r_count_29_io_out ? io_r_328_b : _GEN_22167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22169 = 10'h149 == r_count_29_io_out ? io_r_329_b : _GEN_22168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22170 = 10'h14a == r_count_29_io_out ? io_r_330_b : _GEN_22169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22171 = 10'h14b == r_count_29_io_out ? io_r_331_b : _GEN_22170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22172 = 10'h14c == r_count_29_io_out ? io_r_332_b : _GEN_22171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22173 = 10'h14d == r_count_29_io_out ? io_r_333_b : _GEN_22172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22174 = 10'h14e == r_count_29_io_out ? io_r_334_b : _GEN_22173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22175 = 10'h14f == r_count_29_io_out ? io_r_335_b : _GEN_22174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22176 = 10'h150 == r_count_29_io_out ? io_r_336_b : _GEN_22175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22177 = 10'h151 == r_count_29_io_out ? io_r_337_b : _GEN_22176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22178 = 10'h152 == r_count_29_io_out ? io_r_338_b : _GEN_22177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22179 = 10'h153 == r_count_29_io_out ? io_r_339_b : _GEN_22178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22180 = 10'h154 == r_count_29_io_out ? io_r_340_b : _GEN_22179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22181 = 10'h155 == r_count_29_io_out ? io_r_341_b : _GEN_22180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22182 = 10'h156 == r_count_29_io_out ? io_r_342_b : _GEN_22181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22183 = 10'h157 == r_count_29_io_out ? io_r_343_b : _GEN_22182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22184 = 10'h158 == r_count_29_io_out ? io_r_344_b : _GEN_22183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22185 = 10'h159 == r_count_29_io_out ? io_r_345_b : _GEN_22184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22186 = 10'h15a == r_count_29_io_out ? io_r_346_b : _GEN_22185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22187 = 10'h15b == r_count_29_io_out ? io_r_347_b : _GEN_22186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22188 = 10'h15c == r_count_29_io_out ? io_r_348_b : _GEN_22187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22189 = 10'h15d == r_count_29_io_out ? io_r_349_b : _GEN_22188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22190 = 10'h15e == r_count_29_io_out ? io_r_350_b : _GEN_22189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22191 = 10'h15f == r_count_29_io_out ? io_r_351_b : _GEN_22190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22192 = 10'h160 == r_count_29_io_out ? io_r_352_b : _GEN_22191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22193 = 10'h161 == r_count_29_io_out ? io_r_353_b : _GEN_22192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22194 = 10'h162 == r_count_29_io_out ? io_r_354_b : _GEN_22193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22195 = 10'h163 == r_count_29_io_out ? io_r_355_b : _GEN_22194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22196 = 10'h164 == r_count_29_io_out ? io_r_356_b : _GEN_22195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22197 = 10'h165 == r_count_29_io_out ? io_r_357_b : _GEN_22196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22198 = 10'h166 == r_count_29_io_out ? io_r_358_b : _GEN_22197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22199 = 10'h167 == r_count_29_io_out ? io_r_359_b : _GEN_22198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22200 = 10'h168 == r_count_29_io_out ? io_r_360_b : _GEN_22199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22201 = 10'h169 == r_count_29_io_out ? io_r_361_b : _GEN_22200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22202 = 10'h16a == r_count_29_io_out ? io_r_362_b : _GEN_22201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22203 = 10'h16b == r_count_29_io_out ? io_r_363_b : _GEN_22202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22204 = 10'h16c == r_count_29_io_out ? io_r_364_b : _GEN_22203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22205 = 10'h16d == r_count_29_io_out ? io_r_365_b : _GEN_22204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22206 = 10'h16e == r_count_29_io_out ? io_r_366_b : _GEN_22205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22207 = 10'h16f == r_count_29_io_out ? io_r_367_b : _GEN_22206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22208 = 10'h170 == r_count_29_io_out ? io_r_368_b : _GEN_22207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22209 = 10'h171 == r_count_29_io_out ? io_r_369_b : _GEN_22208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22210 = 10'h172 == r_count_29_io_out ? io_r_370_b : _GEN_22209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22211 = 10'h173 == r_count_29_io_out ? io_r_371_b : _GEN_22210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22212 = 10'h174 == r_count_29_io_out ? io_r_372_b : _GEN_22211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22213 = 10'h175 == r_count_29_io_out ? io_r_373_b : _GEN_22212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22214 = 10'h176 == r_count_29_io_out ? io_r_374_b : _GEN_22213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22215 = 10'h177 == r_count_29_io_out ? io_r_375_b : _GEN_22214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22216 = 10'h178 == r_count_29_io_out ? io_r_376_b : _GEN_22215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22217 = 10'h179 == r_count_29_io_out ? io_r_377_b : _GEN_22216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22218 = 10'h17a == r_count_29_io_out ? io_r_378_b : _GEN_22217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22219 = 10'h17b == r_count_29_io_out ? io_r_379_b : _GEN_22218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22220 = 10'h17c == r_count_29_io_out ? io_r_380_b : _GEN_22219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22221 = 10'h17d == r_count_29_io_out ? io_r_381_b : _GEN_22220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22222 = 10'h17e == r_count_29_io_out ? io_r_382_b : _GEN_22221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22223 = 10'h17f == r_count_29_io_out ? io_r_383_b : _GEN_22222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22224 = 10'h180 == r_count_29_io_out ? io_r_384_b : _GEN_22223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22225 = 10'h181 == r_count_29_io_out ? io_r_385_b : _GEN_22224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22226 = 10'h182 == r_count_29_io_out ? io_r_386_b : _GEN_22225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22227 = 10'h183 == r_count_29_io_out ? io_r_387_b : _GEN_22226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22228 = 10'h184 == r_count_29_io_out ? io_r_388_b : _GEN_22227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22229 = 10'h185 == r_count_29_io_out ? io_r_389_b : _GEN_22228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22230 = 10'h186 == r_count_29_io_out ? io_r_390_b : _GEN_22229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22231 = 10'h187 == r_count_29_io_out ? io_r_391_b : _GEN_22230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22232 = 10'h188 == r_count_29_io_out ? io_r_392_b : _GEN_22231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22233 = 10'h189 == r_count_29_io_out ? io_r_393_b : _GEN_22232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22234 = 10'h18a == r_count_29_io_out ? io_r_394_b : _GEN_22233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22235 = 10'h18b == r_count_29_io_out ? io_r_395_b : _GEN_22234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22236 = 10'h18c == r_count_29_io_out ? io_r_396_b : _GEN_22235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22237 = 10'h18d == r_count_29_io_out ? io_r_397_b : _GEN_22236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22238 = 10'h18e == r_count_29_io_out ? io_r_398_b : _GEN_22237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22239 = 10'h18f == r_count_29_io_out ? io_r_399_b : _GEN_22238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22240 = 10'h190 == r_count_29_io_out ? io_r_400_b : _GEN_22239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22241 = 10'h191 == r_count_29_io_out ? io_r_401_b : _GEN_22240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22242 = 10'h192 == r_count_29_io_out ? io_r_402_b : _GEN_22241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22243 = 10'h193 == r_count_29_io_out ? io_r_403_b : _GEN_22242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22244 = 10'h194 == r_count_29_io_out ? io_r_404_b : _GEN_22243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22245 = 10'h195 == r_count_29_io_out ? io_r_405_b : _GEN_22244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22246 = 10'h196 == r_count_29_io_out ? io_r_406_b : _GEN_22245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22247 = 10'h197 == r_count_29_io_out ? io_r_407_b : _GEN_22246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22248 = 10'h198 == r_count_29_io_out ? io_r_408_b : _GEN_22247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22249 = 10'h199 == r_count_29_io_out ? io_r_409_b : _GEN_22248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22250 = 10'h19a == r_count_29_io_out ? io_r_410_b : _GEN_22249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22251 = 10'h19b == r_count_29_io_out ? io_r_411_b : _GEN_22250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22252 = 10'h19c == r_count_29_io_out ? io_r_412_b : _GEN_22251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22253 = 10'h19d == r_count_29_io_out ? io_r_413_b : _GEN_22252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22254 = 10'h19e == r_count_29_io_out ? io_r_414_b : _GEN_22253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22255 = 10'h19f == r_count_29_io_out ? io_r_415_b : _GEN_22254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22256 = 10'h1a0 == r_count_29_io_out ? io_r_416_b : _GEN_22255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22257 = 10'h1a1 == r_count_29_io_out ? io_r_417_b : _GEN_22256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22258 = 10'h1a2 == r_count_29_io_out ? io_r_418_b : _GEN_22257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22259 = 10'h1a3 == r_count_29_io_out ? io_r_419_b : _GEN_22258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22260 = 10'h1a4 == r_count_29_io_out ? io_r_420_b : _GEN_22259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22261 = 10'h1a5 == r_count_29_io_out ? io_r_421_b : _GEN_22260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22262 = 10'h1a6 == r_count_29_io_out ? io_r_422_b : _GEN_22261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22263 = 10'h1a7 == r_count_29_io_out ? io_r_423_b : _GEN_22262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22264 = 10'h1a8 == r_count_29_io_out ? io_r_424_b : _GEN_22263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22265 = 10'h1a9 == r_count_29_io_out ? io_r_425_b : _GEN_22264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22266 = 10'h1aa == r_count_29_io_out ? io_r_426_b : _GEN_22265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22267 = 10'h1ab == r_count_29_io_out ? io_r_427_b : _GEN_22266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22268 = 10'h1ac == r_count_29_io_out ? io_r_428_b : _GEN_22267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22269 = 10'h1ad == r_count_29_io_out ? io_r_429_b : _GEN_22268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22270 = 10'h1ae == r_count_29_io_out ? io_r_430_b : _GEN_22269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22271 = 10'h1af == r_count_29_io_out ? io_r_431_b : _GEN_22270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22272 = 10'h1b0 == r_count_29_io_out ? io_r_432_b : _GEN_22271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22273 = 10'h1b1 == r_count_29_io_out ? io_r_433_b : _GEN_22272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22274 = 10'h1b2 == r_count_29_io_out ? io_r_434_b : _GEN_22273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22275 = 10'h1b3 == r_count_29_io_out ? io_r_435_b : _GEN_22274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22276 = 10'h1b4 == r_count_29_io_out ? io_r_436_b : _GEN_22275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22277 = 10'h1b5 == r_count_29_io_out ? io_r_437_b : _GEN_22276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22278 = 10'h1b6 == r_count_29_io_out ? io_r_438_b : _GEN_22277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22279 = 10'h1b7 == r_count_29_io_out ? io_r_439_b : _GEN_22278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22280 = 10'h1b8 == r_count_29_io_out ? io_r_440_b : _GEN_22279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22281 = 10'h1b9 == r_count_29_io_out ? io_r_441_b : _GEN_22280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22282 = 10'h1ba == r_count_29_io_out ? io_r_442_b : _GEN_22281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22283 = 10'h1bb == r_count_29_io_out ? io_r_443_b : _GEN_22282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22284 = 10'h1bc == r_count_29_io_out ? io_r_444_b : _GEN_22283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22285 = 10'h1bd == r_count_29_io_out ? io_r_445_b : _GEN_22284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22286 = 10'h1be == r_count_29_io_out ? io_r_446_b : _GEN_22285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22287 = 10'h1bf == r_count_29_io_out ? io_r_447_b : _GEN_22286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22288 = 10'h1c0 == r_count_29_io_out ? io_r_448_b : _GEN_22287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22289 = 10'h1c1 == r_count_29_io_out ? io_r_449_b : _GEN_22288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22290 = 10'h1c2 == r_count_29_io_out ? io_r_450_b : _GEN_22289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22291 = 10'h1c3 == r_count_29_io_out ? io_r_451_b : _GEN_22290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22292 = 10'h1c4 == r_count_29_io_out ? io_r_452_b : _GEN_22291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22293 = 10'h1c5 == r_count_29_io_out ? io_r_453_b : _GEN_22292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22294 = 10'h1c6 == r_count_29_io_out ? io_r_454_b : _GEN_22293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22295 = 10'h1c7 == r_count_29_io_out ? io_r_455_b : _GEN_22294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22296 = 10'h1c8 == r_count_29_io_out ? io_r_456_b : _GEN_22295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22297 = 10'h1c9 == r_count_29_io_out ? io_r_457_b : _GEN_22296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22298 = 10'h1ca == r_count_29_io_out ? io_r_458_b : _GEN_22297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22299 = 10'h1cb == r_count_29_io_out ? io_r_459_b : _GEN_22298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22300 = 10'h1cc == r_count_29_io_out ? io_r_460_b : _GEN_22299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22301 = 10'h1cd == r_count_29_io_out ? io_r_461_b : _GEN_22300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22302 = 10'h1ce == r_count_29_io_out ? io_r_462_b : _GEN_22301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22303 = 10'h1cf == r_count_29_io_out ? io_r_463_b : _GEN_22302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22304 = 10'h1d0 == r_count_29_io_out ? io_r_464_b : _GEN_22303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22305 = 10'h1d1 == r_count_29_io_out ? io_r_465_b : _GEN_22304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22306 = 10'h1d2 == r_count_29_io_out ? io_r_466_b : _GEN_22305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22307 = 10'h1d3 == r_count_29_io_out ? io_r_467_b : _GEN_22306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22308 = 10'h1d4 == r_count_29_io_out ? io_r_468_b : _GEN_22307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22309 = 10'h1d5 == r_count_29_io_out ? io_r_469_b : _GEN_22308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22310 = 10'h1d6 == r_count_29_io_out ? io_r_470_b : _GEN_22309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22311 = 10'h1d7 == r_count_29_io_out ? io_r_471_b : _GEN_22310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22312 = 10'h1d8 == r_count_29_io_out ? io_r_472_b : _GEN_22311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22313 = 10'h1d9 == r_count_29_io_out ? io_r_473_b : _GEN_22312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22314 = 10'h1da == r_count_29_io_out ? io_r_474_b : _GEN_22313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22315 = 10'h1db == r_count_29_io_out ? io_r_475_b : _GEN_22314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22316 = 10'h1dc == r_count_29_io_out ? io_r_476_b : _GEN_22315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22317 = 10'h1dd == r_count_29_io_out ? io_r_477_b : _GEN_22316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22318 = 10'h1de == r_count_29_io_out ? io_r_478_b : _GEN_22317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22319 = 10'h1df == r_count_29_io_out ? io_r_479_b : _GEN_22318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22320 = 10'h1e0 == r_count_29_io_out ? io_r_480_b : _GEN_22319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22321 = 10'h1e1 == r_count_29_io_out ? io_r_481_b : _GEN_22320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22322 = 10'h1e2 == r_count_29_io_out ? io_r_482_b : _GEN_22321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22323 = 10'h1e3 == r_count_29_io_out ? io_r_483_b : _GEN_22322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22324 = 10'h1e4 == r_count_29_io_out ? io_r_484_b : _GEN_22323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22325 = 10'h1e5 == r_count_29_io_out ? io_r_485_b : _GEN_22324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22326 = 10'h1e6 == r_count_29_io_out ? io_r_486_b : _GEN_22325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22327 = 10'h1e7 == r_count_29_io_out ? io_r_487_b : _GEN_22326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22328 = 10'h1e8 == r_count_29_io_out ? io_r_488_b : _GEN_22327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22329 = 10'h1e9 == r_count_29_io_out ? io_r_489_b : _GEN_22328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22330 = 10'h1ea == r_count_29_io_out ? io_r_490_b : _GEN_22329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22331 = 10'h1eb == r_count_29_io_out ? io_r_491_b : _GEN_22330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22332 = 10'h1ec == r_count_29_io_out ? io_r_492_b : _GEN_22331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22333 = 10'h1ed == r_count_29_io_out ? io_r_493_b : _GEN_22332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22334 = 10'h1ee == r_count_29_io_out ? io_r_494_b : _GEN_22333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22335 = 10'h1ef == r_count_29_io_out ? io_r_495_b : _GEN_22334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22336 = 10'h1f0 == r_count_29_io_out ? io_r_496_b : _GEN_22335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22337 = 10'h1f1 == r_count_29_io_out ? io_r_497_b : _GEN_22336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22338 = 10'h1f2 == r_count_29_io_out ? io_r_498_b : _GEN_22337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22339 = 10'h1f3 == r_count_29_io_out ? io_r_499_b : _GEN_22338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22340 = 10'h1f4 == r_count_29_io_out ? io_r_500_b : _GEN_22339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22341 = 10'h1f5 == r_count_29_io_out ? io_r_501_b : _GEN_22340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22342 = 10'h1f6 == r_count_29_io_out ? io_r_502_b : _GEN_22341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22343 = 10'h1f7 == r_count_29_io_out ? io_r_503_b : _GEN_22342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22344 = 10'h1f8 == r_count_29_io_out ? io_r_504_b : _GEN_22343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22345 = 10'h1f9 == r_count_29_io_out ? io_r_505_b : _GEN_22344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22346 = 10'h1fa == r_count_29_io_out ? io_r_506_b : _GEN_22345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22347 = 10'h1fb == r_count_29_io_out ? io_r_507_b : _GEN_22346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22348 = 10'h1fc == r_count_29_io_out ? io_r_508_b : _GEN_22347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22349 = 10'h1fd == r_count_29_io_out ? io_r_509_b : _GEN_22348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22350 = 10'h1fe == r_count_29_io_out ? io_r_510_b : _GEN_22349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22351 = 10'h1ff == r_count_29_io_out ? io_r_511_b : _GEN_22350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22352 = 10'h200 == r_count_29_io_out ? io_r_512_b : _GEN_22351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22353 = 10'h201 == r_count_29_io_out ? io_r_513_b : _GEN_22352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22354 = 10'h202 == r_count_29_io_out ? io_r_514_b : _GEN_22353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22355 = 10'h203 == r_count_29_io_out ? io_r_515_b : _GEN_22354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22356 = 10'h204 == r_count_29_io_out ? io_r_516_b : _GEN_22355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22357 = 10'h205 == r_count_29_io_out ? io_r_517_b : _GEN_22356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22358 = 10'h206 == r_count_29_io_out ? io_r_518_b : _GEN_22357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22359 = 10'h207 == r_count_29_io_out ? io_r_519_b : _GEN_22358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22360 = 10'h208 == r_count_29_io_out ? io_r_520_b : _GEN_22359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22361 = 10'h209 == r_count_29_io_out ? io_r_521_b : _GEN_22360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22362 = 10'h20a == r_count_29_io_out ? io_r_522_b : _GEN_22361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22363 = 10'h20b == r_count_29_io_out ? io_r_523_b : _GEN_22362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22364 = 10'h20c == r_count_29_io_out ? io_r_524_b : _GEN_22363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22365 = 10'h20d == r_count_29_io_out ? io_r_525_b : _GEN_22364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22366 = 10'h20e == r_count_29_io_out ? io_r_526_b : _GEN_22365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22367 = 10'h20f == r_count_29_io_out ? io_r_527_b : _GEN_22366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22368 = 10'h210 == r_count_29_io_out ? io_r_528_b : _GEN_22367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22369 = 10'h211 == r_count_29_io_out ? io_r_529_b : _GEN_22368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22370 = 10'h212 == r_count_29_io_out ? io_r_530_b : _GEN_22369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22371 = 10'h213 == r_count_29_io_out ? io_r_531_b : _GEN_22370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22372 = 10'h214 == r_count_29_io_out ? io_r_532_b : _GEN_22371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22373 = 10'h215 == r_count_29_io_out ? io_r_533_b : _GEN_22372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22374 = 10'h216 == r_count_29_io_out ? io_r_534_b : _GEN_22373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22375 = 10'h217 == r_count_29_io_out ? io_r_535_b : _GEN_22374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22376 = 10'h218 == r_count_29_io_out ? io_r_536_b : _GEN_22375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22377 = 10'h219 == r_count_29_io_out ? io_r_537_b : _GEN_22376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22378 = 10'h21a == r_count_29_io_out ? io_r_538_b : _GEN_22377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22379 = 10'h21b == r_count_29_io_out ? io_r_539_b : _GEN_22378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22380 = 10'h21c == r_count_29_io_out ? io_r_540_b : _GEN_22379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22381 = 10'h21d == r_count_29_io_out ? io_r_541_b : _GEN_22380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22382 = 10'h21e == r_count_29_io_out ? io_r_542_b : _GEN_22381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22383 = 10'h21f == r_count_29_io_out ? io_r_543_b : _GEN_22382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22384 = 10'h220 == r_count_29_io_out ? io_r_544_b : _GEN_22383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22385 = 10'h221 == r_count_29_io_out ? io_r_545_b : _GEN_22384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22386 = 10'h222 == r_count_29_io_out ? io_r_546_b : _GEN_22385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22387 = 10'h223 == r_count_29_io_out ? io_r_547_b : _GEN_22386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22388 = 10'h224 == r_count_29_io_out ? io_r_548_b : _GEN_22387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22389 = 10'h225 == r_count_29_io_out ? io_r_549_b : _GEN_22388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22390 = 10'h226 == r_count_29_io_out ? io_r_550_b : _GEN_22389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22391 = 10'h227 == r_count_29_io_out ? io_r_551_b : _GEN_22390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22392 = 10'h228 == r_count_29_io_out ? io_r_552_b : _GEN_22391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22393 = 10'h229 == r_count_29_io_out ? io_r_553_b : _GEN_22392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22394 = 10'h22a == r_count_29_io_out ? io_r_554_b : _GEN_22393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22395 = 10'h22b == r_count_29_io_out ? io_r_555_b : _GEN_22394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22396 = 10'h22c == r_count_29_io_out ? io_r_556_b : _GEN_22395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22397 = 10'h22d == r_count_29_io_out ? io_r_557_b : _GEN_22396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22398 = 10'h22e == r_count_29_io_out ? io_r_558_b : _GEN_22397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22399 = 10'h22f == r_count_29_io_out ? io_r_559_b : _GEN_22398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22400 = 10'h230 == r_count_29_io_out ? io_r_560_b : _GEN_22399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22401 = 10'h231 == r_count_29_io_out ? io_r_561_b : _GEN_22400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22402 = 10'h232 == r_count_29_io_out ? io_r_562_b : _GEN_22401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22403 = 10'h233 == r_count_29_io_out ? io_r_563_b : _GEN_22402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22404 = 10'h234 == r_count_29_io_out ? io_r_564_b : _GEN_22403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22405 = 10'h235 == r_count_29_io_out ? io_r_565_b : _GEN_22404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22406 = 10'h236 == r_count_29_io_out ? io_r_566_b : _GEN_22405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22407 = 10'h237 == r_count_29_io_out ? io_r_567_b : _GEN_22406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22408 = 10'h238 == r_count_29_io_out ? io_r_568_b : _GEN_22407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22409 = 10'h239 == r_count_29_io_out ? io_r_569_b : _GEN_22408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22410 = 10'h23a == r_count_29_io_out ? io_r_570_b : _GEN_22409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22411 = 10'h23b == r_count_29_io_out ? io_r_571_b : _GEN_22410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22412 = 10'h23c == r_count_29_io_out ? io_r_572_b : _GEN_22411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22413 = 10'h23d == r_count_29_io_out ? io_r_573_b : _GEN_22412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22414 = 10'h23e == r_count_29_io_out ? io_r_574_b : _GEN_22413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22415 = 10'h23f == r_count_29_io_out ? io_r_575_b : _GEN_22414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22416 = 10'h240 == r_count_29_io_out ? io_r_576_b : _GEN_22415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22417 = 10'h241 == r_count_29_io_out ? io_r_577_b : _GEN_22416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22418 = 10'h242 == r_count_29_io_out ? io_r_578_b : _GEN_22417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22419 = 10'h243 == r_count_29_io_out ? io_r_579_b : _GEN_22418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22420 = 10'h244 == r_count_29_io_out ? io_r_580_b : _GEN_22419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22421 = 10'h245 == r_count_29_io_out ? io_r_581_b : _GEN_22420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22422 = 10'h246 == r_count_29_io_out ? io_r_582_b : _GEN_22421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22423 = 10'h247 == r_count_29_io_out ? io_r_583_b : _GEN_22422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22424 = 10'h248 == r_count_29_io_out ? io_r_584_b : _GEN_22423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22425 = 10'h249 == r_count_29_io_out ? io_r_585_b : _GEN_22424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22426 = 10'h24a == r_count_29_io_out ? io_r_586_b : _GEN_22425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22427 = 10'h24b == r_count_29_io_out ? io_r_587_b : _GEN_22426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22428 = 10'h24c == r_count_29_io_out ? io_r_588_b : _GEN_22427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22429 = 10'h24d == r_count_29_io_out ? io_r_589_b : _GEN_22428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22430 = 10'h24e == r_count_29_io_out ? io_r_590_b : _GEN_22429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22431 = 10'h24f == r_count_29_io_out ? io_r_591_b : _GEN_22430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22432 = 10'h250 == r_count_29_io_out ? io_r_592_b : _GEN_22431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22433 = 10'h251 == r_count_29_io_out ? io_r_593_b : _GEN_22432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22434 = 10'h252 == r_count_29_io_out ? io_r_594_b : _GEN_22433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22435 = 10'h253 == r_count_29_io_out ? io_r_595_b : _GEN_22434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22436 = 10'h254 == r_count_29_io_out ? io_r_596_b : _GEN_22435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22437 = 10'h255 == r_count_29_io_out ? io_r_597_b : _GEN_22436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22438 = 10'h256 == r_count_29_io_out ? io_r_598_b : _GEN_22437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22439 = 10'h257 == r_count_29_io_out ? io_r_599_b : _GEN_22438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22440 = 10'h258 == r_count_29_io_out ? io_r_600_b : _GEN_22439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22441 = 10'h259 == r_count_29_io_out ? io_r_601_b : _GEN_22440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22442 = 10'h25a == r_count_29_io_out ? io_r_602_b : _GEN_22441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22443 = 10'h25b == r_count_29_io_out ? io_r_603_b : _GEN_22442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22444 = 10'h25c == r_count_29_io_out ? io_r_604_b : _GEN_22443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22445 = 10'h25d == r_count_29_io_out ? io_r_605_b : _GEN_22444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22446 = 10'h25e == r_count_29_io_out ? io_r_606_b : _GEN_22445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22447 = 10'h25f == r_count_29_io_out ? io_r_607_b : _GEN_22446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22448 = 10'h260 == r_count_29_io_out ? io_r_608_b : _GEN_22447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22449 = 10'h261 == r_count_29_io_out ? io_r_609_b : _GEN_22448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22450 = 10'h262 == r_count_29_io_out ? io_r_610_b : _GEN_22449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22451 = 10'h263 == r_count_29_io_out ? io_r_611_b : _GEN_22450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22452 = 10'h264 == r_count_29_io_out ? io_r_612_b : _GEN_22451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22453 = 10'h265 == r_count_29_io_out ? io_r_613_b : _GEN_22452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22454 = 10'h266 == r_count_29_io_out ? io_r_614_b : _GEN_22453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22455 = 10'h267 == r_count_29_io_out ? io_r_615_b : _GEN_22454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22456 = 10'h268 == r_count_29_io_out ? io_r_616_b : _GEN_22455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22457 = 10'h269 == r_count_29_io_out ? io_r_617_b : _GEN_22456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22458 = 10'h26a == r_count_29_io_out ? io_r_618_b : _GEN_22457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22459 = 10'h26b == r_count_29_io_out ? io_r_619_b : _GEN_22458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22460 = 10'h26c == r_count_29_io_out ? io_r_620_b : _GEN_22459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22461 = 10'h26d == r_count_29_io_out ? io_r_621_b : _GEN_22460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22462 = 10'h26e == r_count_29_io_out ? io_r_622_b : _GEN_22461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22463 = 10'h26f == r_count_29_io_out ? io_r_623_b : _GEN_22462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22464 = 10'h270 == r_count_29_io_out ? io_r_624_b : _GEN_22463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22465 = 10'h271 == r_count_29_io_out ? io_r_625_b : _GEN_22464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22466 = 10'h272 == r_count_29_io_out ? io_r_626_b : _GEN_22465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22467 = 10'h273 == r_count_29_io_out ? io_r_627_b : _GEN_22466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22468 = 10'h274 == r_count_29_io_out ? io_r_628_b : _GEN_22467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22469 = 10'h275 == r_count_29_io_out ? io_r_629_b : _GEN_22468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22470 = 10'h276 == r_count_29_io_out ? io_r_630_b : _GEN_22469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22471 = 10'h277 == r_count_29_io_out ? io_r_631_b : _GEN_22470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22472 = 10'h278 == r_count_29_io_out ? io_r_632_b : _GEN_22471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22473 = 10'h279 == r_count_29_io_out ? io_r_633_b : _GEN_22472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22474 = 10'h27a == r_count_29_io_out ? io_r_634_b : _GEN_22473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22475 = 10'h27b == r_count_29_io_out ? io_r_635_b : _GEN_22474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22476 = 10'h27c == r_count_29_io_out ? io_r_636_b : _GEN_22475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22477 = 10'h27d == r_count_29_io_out ? io_r_637_b : _GEN_22476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22478 = 10'h27e == r_count_29_io_out ? io_r_638_b : _GEN_22477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22479 = 10'h27f == r_count_29_io_out ? io_r_639_b : _GEN_22478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22480 = 10'h280 == r_count_29_io_out ? io_r_640_b : _GEN_22479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22481 = 10'h281 == r_count_29_io_out ? io_r_641_b : _GEN_22480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22482 = 10'h282 == r_count_29_io_out ? io_r_642_b : _GEN_22481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22483 = 10'h283 == r_count_29_io_out ? io_r_643_b : _GEN_22482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22484 = 10'h284 == r_count_29_io_out ? io_r_644_b : _GEN_22483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22485 = 10'h285 == r_count_29_io_out ? io_r_645_b : _GEN_22484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22486 = 10'h286 == r_count_29_io_out ? io_r_646_b : _GEN_22485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22487 = 10'h287 == r_count_29_io_out ? io_r_647_b : _GEN_22486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22488 = 10'h288 == r_count_29_io_out ? io_r_648_b : _GEN_22487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22489 = 10'h289 == r_count_29_io_out ? io_r_649_b : _GEN_22488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22490 = 10'h28a == r_count_29_io_out ? io_r_650_b : _GEN_22489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22491 = 10'h28b == r_count_29_io_out ? io_r_651_b : _GEN_22490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22492 = 10'h28c == r_count_29_io_out ? io_r_652_b : _GEN_22491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22493 = 10'h28d == r_count_29_io_out ? io_r_653_b : _GEN_22492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22494 = 10'h28e == r_count_29_io_out ? io_r_654_b : _GEN_22493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22495 = 10'h28f == r_count_29_io_out ? io_r_655_b : _GEN_22494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22496 = 10'h290 == r_count_29_io_out ? io_r_656_b : _GEN_22495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22497 = 10'h291 == r_count_29_io_out ? io_r_657_b : _GEN_22496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22498 = 10'h292 == r_count_29_io_out ? io_r_658_b : _GEN_22497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22499 = 10'h293 == r_count_29_io_out ? io_r_659_b : _GEN_22498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22500 = 10'h294 == r_count_29_io_out ? io_r_660_b : _GEN_22499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22501 = 10'h295 == r_count_29_io_out ? io_r_661_b : _GEN_22500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22502 = 10'h296 == r_count_29_io_out ? io_r_662_b : _GEN_22501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22503 = 10'h297 == r_count_29_io_out ? io_r_663_b : _GEN_22502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22504 = 10'h298 == r_count_29_io_out ? io_r_664_b : _GEN_22503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22505 = 10'h299 == r_count_29_io_out ? io_r_665_b : _GEN_22504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22506 = 10'h29a == r_count_29_io_out ? io_r_666_b : _GEN_22505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22507 = 10'h29b == r_count_29_io_out ? io_r_667_b : _GEN_22506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22508 = 10'h29c == r_count_29_io_out ? io_r_668_b : _GEN_22507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22509 = 10'h29d == r_count_29_io_out ? io_r_669_b : _GEN_22508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22510 = 10'h29e == r_count_29_io_out ? io_r_670_b : _GEN_22509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22511 = 10'h29f == r_count_29_io_out ? io_r_671_b : _GEN_22510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22512 = 10'h2a0 == r_count_29_io_out ? io_r_672_b : _GEN_22511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22513 = 10'h2a1 == r_count_29_io_out ? io_r_673_b : _GEN_22512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22514 = 10'h2a2 == r_count_29_io_out ? io_r_674_b : _GEN_22513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22515 = 10'h2a3 == r_count_29_io_out ? io_r_675_b : _GEN_22514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22516 = 10'h2a4 == r_count_29_io_out ? io_r_676_b : _GEN_22515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22517 = 10'h2a5 == r_count_29_io_out ? io_r_677_b : _GEN_22516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22518 = 10'h2a6 == r_count_29_io_out ? io_r_678_b : _GEN_22517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22519 = 10'h2a7 == r_count_29_io_out ? io_r_679_b : _GEN_22518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22520 = 10'h2a8 == r_count_29_io_out ? io_r_680_b : _GEN_22519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22521 = 10'h2a9 == r_count_29_io_out ? io_r_681_b : _GEN_22520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22522 = 10'h2aa == r_count_29_io_out ? io_r_682_b : _GEN_22521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22523 = 10'h2ab == r_count_29_io_out ? io_r_683_b : _GEN_22522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22524 = 10'h2ac == r_count_29_io_out ? io_r_684_b : _GEN_22523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22525 = 10'h2ad == r_count_29_io_out ? io_r_685_b : _GEN_22524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22526 = 10'h2ae == r_count_29_io_out ? io_r_686_b : _GEN_22525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22527 = 10'h2af == r_count_29_io_out ? io_r_687_b : _GEN_22526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22528 = 10'h2b0 == r_count_29_io_out ? io_r_688_b : _GEN_22527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22529 = 10'h2b1 == r_count_29_io_out ? io_r_689_b : _GEN_22528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22530 = 10'h2b2 == r_count_29_io_out ? io_r_690_b : _GEN_22529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22531 = 10'h2b3 == r_count_29_io_out ? io_r_691_b : _GEN_22530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22532 = 10'h2b4 == r_count_29_io_out ? io_r_692_b : _GEN_22531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22533 = 10'h2b5 == r_count_29_io_out ? io_r_693_b : _GEN_22532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22534 = 10'h2b6 == r_count_29_io_out ? io_r_694_b : _GEN_22533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22535 = 10'h2b7 == r_count_29_io_out ? io_r_695_b : _GEN_22534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22536 = 10'h2b8 == r_count_29_io_out ? io_r_696_b : _GEN_22535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22537 = 10'h2b9 == r_count_29_io_out ? io_r_697_b : _GEN_22536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22538 = 10'h2ba == r_count_29_io_out ? io_r_698_b : _GEN_22537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22539 = 10'h2bb == r_count_29_io_out ? io_r_699_b : _GEN_22538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22540 = 10'h2bc == r_count_29_io_out ? io_r_700_b : _GEN_22539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22541 = 10'h2bd == r_count_29_io_out ? io_r_701_b : _GEN_22540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22542 = 10'h2be == r_count_29_io_out ? io_r_702_b : _GEN_22541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22543 = 10'h2bf == r_count_29_io_out ? io_r_703_b : _GEN_22542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22544 = 10'h2c0 == r_count_29_io_out ? io_r_704_b : _GEN_22543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22545 = 10'h2c1 == r_count_29_io_out ? io_r_705_b : _GEN_22544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22546 = 10'h2c2 == r_count_29_io_out ? io_r_706_b : _GEN_22545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22547 = 10'h2c3 == r_count_29_io_out ? io_r_707_b : _GEN_22546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22548 = 10'h2c4 == r_count_29_io_out ? io_r_708_b : _GEN_22547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22549 = 10'h2c5 == r_count_29_io_out ? io_r_709_b : _GEN_22548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22550 = 10'h2c6 == r_count_29_io_out ? io_r_710_b : _GEN_22549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22551 = 10'h2c7 == r_count_29_io_out ? io_r_711_b : _GEN_22550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22552 = 10'h2c8 == r_count_29_io_out ? io_r_712_b : _GEN_22551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22553 = 10'h2c9 == r_count_29_io_out ? io_r_713_b : _GEN_22552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22554 = 10'h2ca == r_count_29_io_out ? io_r_714_b : _GEN_22553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22555 = 10'h2cb == r_count_29_io_out ? io_r_715_b : _GEN_22554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22556 = 10'h2cc == r_count_29_io_out ? io_r_716_b : _GEN_22555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22557 = 10'h2cd == r_count_29_io_out ? io_r_717_b : _GEN_22556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22558 = 10'h2ce == r_count_29_io_out ? io_r_718_b : _GEN_22557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22559 = 10'h2cf == r_count_29_io_out ? io_r_719_b : _GEN_22558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22560 = 10'h2d0 == r_count_29_io_out ? io_r_720_b : _GEN_22559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22561 = 10'h2d1 == r_count_29_io_out ? io_r_721_b : _GEN_22560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22562 = 10'h2d2 == r_count_29_io_out ? io_r_722_b : _GEN_22561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22563 = 10'h2d3 == r_count_29_io_out ? io_r_723_b : _GEN_22562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22564 = 10'h2d4 == r_count_29_io_out ? io_r_724_b : _GEN_22563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22565 = 10'h2d5 == r_count_29_io_out ? io_r_725_b : _GEN_22564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22566 = 10'h2d6 == r_count_29_io_out ? io_r_726_b : _GEN_22565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22567 = 10'h2d7 == r_count_29_io_out ? io_r_727_b : _GEN_22566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22568 = 10'h2d8 == r_count_29_io_out ? io_r_728_b : _GEN_22567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22569 = 10'h2d9 == r_count_29_io_out ? io_r_729_b : _GEN_22568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22570 = 10'h2da == r_count_29_io_out ? io_r_730_b : _GEN_22569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22571 = 10'h2db == r_count_29_io_out ? io_r_731_b : _GEN_22570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22572 = 10'h2dc == r_count_29_io_out ? io_r_732_b : _GEN_22571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22573 = 10'h2dd == r_count_29_io_out ? io_r_733_b : _GEN_22572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22574 = 10'h2de == r_count_29_io_out ? io_r_734_b : _GEN_22573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22575 = 10'h2df == r_count_29_io_out ? io_r_735_b : _GEN_22574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22576 = 10'h2e0 == r_count_29_io_out ? io_r_736_b : _GEN_22575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22577 = 10'h2e1 == r_count_29_io_out ? io_r_737_b : _GEN_22576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22578 = 10'h2e2 == r_count_29_io_out ? io_r_738_b : _GEN_22577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22579 = 10'h2e3 == r_count_29_io_out ? io_r_739_b : _GEN_22578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22580 = 10'h2e4 == r_count_29_io_out ? io_r_740_b : _GEN_22579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22581 = 10'h2e5 == r_count_29_io_out ? io_r_741_b : _GEN_22580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22582 = 10'h2e6 == r_count_29_io_out ? io_r_742_b : _GEN_22581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22583 = 10'h2e7 == r_count_29_io_out ? io_r_743_b : _GEN_22582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22584 = 10'h2e8 == r_count_29_io_out ? io_r_744_b : _GEN_22583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22585 = 10'h2e9 == r_count_29_io_out ? io_r_745_b : _GEN_22584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22586 = 10'h2ea == r_count_29_io_out ? io_r_746_b : _GEN_22585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22587 = 10'h2eb == r_count_29_io_out ? io_r_747_b : _GEN_22586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_22588 = 10'h2ec == r_count_29_io_out ? io_r_748_b : _GEN_22587; // @[SWChisel.scala 221:{19,19}]
  SWCell array_0 ( // @[SWChisel.scala 170:39]
    .io_q(array_0_io_q),
    .io_r(array_0_io_r),
    .io_e_i(array_0_io_e_i),
    .io_f_i(array_0_io_f_i),
    .io_ve_i(array_0_io_ve_i),
    .io_vf_i(array_0_io_vf_i),
    .io_vv_i(array_0_io_vv_i),
    .io_e_o(array_0_io_e_o),
    .io_f_o(array_0_io_f_o),
    .io_v_o(array_0_io_v_o)
  );
  SWCell array_1 ( // @[SWChisel.scala 170:39]
    .io_q(array_1_io_q),
    .io_r(array_1_io_r),
    .io_e_i(array_1_io_e_i),
    .io_f_i(array_1_io_f_i),
    .io_ve_i(array_1_io_ve_i),
    .io_vf_i(array_1_io_vf_i),
    .io_vv_i(array_1_io_vv_i),
    .io_e_o(array_1_io_e_o),
    .io_f_o(array_1_io_f_o),
    .io_v_o(array_1_io_v_o)
  );
  SWCell array_2 ( // @[SWChisel.scala 170:39]
    .io_q(array_2_io_q),
    .io_r(array_2_io_r),
    .io_e_i(array_2_io_e_i),
    .io_f_i(array_2_io_f_i),
    .io_ve_i(array_2_io_ve_i),
    .io_vf_i(array_2_io_vf_i),
    .io_vv_i(array_2_io_vv_i),
    .io_e_o(array_2_io_e_o),
    .io_f_o(array_2_io_f_o),
    .io_v_o(array_2_io_v_o)
  );
  SWCell array_3 ( // @[SWChisel.scala 170:39]
    .io_q(array_3_io_q),
    .io_r(array_3_io_r),
    .io_e_i(array_3_io_e_i),
    .io_f_i(array_3_io_f_i),
    .io_ve_i(array_3_io_ve_i),
    .io_vf_i(array_3_io_vf_i),
    .io_vv_i(array_3_io_vv_i),
    .io_e_o(array_3_io_e_o),
    .io_f_o(array_3_io_f_o),
    .io_v_o(array_3_io_v_o)
  );
  SWCell array_4 ( // @[SWChisel.scala 170:39]
    .io_q(array_4_io_q),
    .io_r(array_4_io_r),
    .io_e_i(array_4_io_e_i),
    .io_f_i(array_4_io_f_i),
    .io_ve_i(array_4_io_ve_i),
    .io_vf_i(array_4_io_vf_i),
    .io_vv_i(array_4_io_vv_i),
    .io_e_o(array_4_io_e_o),
    .io_f_o(array_4_io_f_o),
    .io_v_o(array_4_io_v_o)
  );
  SWCell array_5 ( // @[SWChisel.scala 170:39]
    .io_q(array_5_io_q),
    .io_r(array_5_io_r),
    .io_e_i(array_5_io_e_i),
    .io_f_i(array_5_io_f_i),
    .io_ve_i(array_5_io_ve_i),
    .io_vf_i(array_5_io_vf_i),
    .io_vv_i(array_5_io_vv_i),
    .io_e_o(array_5_io_e_o),
    .io_f_o(array_5_io_f_o),
    .io_v_o(array_5_io_v_o)
  );
  SWCell array_6 ( // @[SWChisel.scala 170:39]
    .io_q(array_6_io_q),
    .io_r(array_6_io_r),
    .io_e_i(array_6_io_e_i),
    .io_f_i(array_6_io_f_i),
    .io_ve_i(array_6_io_ve_i),
    .io_vf_i(array_6_io_vf_i),
    .io_vv_i(array_6_io_vv_i),
    .io_e_o(array_6_io_e_o),
    .io_f_o(array_6_io_f_o),
    .io_v_o(array_6_io_v_o)
  );
  SWCell array_7 ( // @[SWChisel.scala 170:39]
    .io_q(array_7_io_q),
    .io_r(array_7_io_r),
    .io_e_i(array_7_io_e_i),
    .io_f_i(array_7_io_f_i),
    .io_ve_i(array_7_io_ve_i),
    .io_vf_i(array_7_io_vf_i),
    .io_vv_i(array_7_io_vv_i),
    .io_e_o(array_7_io_e_o),
    .io_f_o(array_7_io_f_o),
    .io_v_o(array_7_io_v_o)
  );
  SWCell array_8 ( // @[SWChisel.scala 170:39]
    .io_q(array_8_io_q),
    .io_r(array_8_io_r),
    .io_e_i(array_8_io_e_i),
    .io_f_i(array_8_io_f_i),
    .io_ve_i(array_8_io_ve_i),
    .io_vf_i(array_8_io_vf_i),
    .io_vv_i(array_8_io_vv_i),
    .io_e_o(array_8_io_e_o),
    .io_f_o(array_8_io_f_o),
    .io_v_o(array_8_io_v_o)
  );
  SWCell array_9 ( // @[SWChisel.scala 170:39]
    .io_q(array_9_io_q),
    .io_r(array_9_io_r),
    .io_e_i(array_9_io_e_i),
    .io_f_i(array_9_io_f_i),
    .io_ve_i(array_9_io_ve_i),
    .io_vf_i(array_9_io_vf_i),
    .io_vv_i(array_9_io_vv_i),
    .io_e_o(array_9_io_e_o),
    .io_f_o(array_9_io_f_o),
    .io_v_o(array_9_io_v_o)
  );
  SWCell array_10 ( // @[SWChisel.scala 170:39]
    .io_q(array_10_io_q),
    .io_r(array_10_io_r),
    .io_e_i(array_10_io_e_i),
    .io_f_i(array_10_io_f_i),
    .io_ve_i(array_10_io_ve_i),
    .io_vf_i(array_10_io_vf_i),
    .io_vv_i(array_10_io_vv_i),
    .io_e_o(array_10_io_e_o),
    .io_f_o(array_10_io_f_o),
    .io_v_o(array_10_io_v_o)
  );
  SWCell array_11 ( // @[SWChisel.scala 170:39]
    .io_q(array_11_io_q),
    .io_r(array_11_io_r),
    .io_e_i(array_11_io_e_i),
    .io_f_i(array_11_io_f_i),
    .io_ve_i(array_11_io_ve_i),
    .io_vf_i(array_11_io_vf_i),
    .io_vv_i(array_11_io_vv_i),
    .io_e_o(array_11_io_e_o),
    .io_f_o(array_11_io_f_o),
    .io_v_o(array_11_io_v_o)
  );
  SWCell array_12 ( // @[SWChisel.scala 170:39]
    .io_q(array_12_io_q),
    .io_r(array_12_io_r),
    .io_e_i(array_12_io_e_i),
    .io_f_i(array_12_io_f_i),
    .io_ve_i(array_12_io_ve_i),
    .io_vf_i(array_12_io_vf_i),
    .io_vv_i(array_12_io_vv_i),
    .io_e_o(array_12_io_e_o),
    .io_f_o(array_12_io_f_o),
    .io_v_o(array_12_io_v_o)
  );
  SWCell array_13 ( // @[SWChisel.scala 170:39]
    .io_q(array_13_io_q),
    .io_r(array_13_io_r),
    .io_e_i(array_13_io_e_i),
    .io_f_i(array_13_io_f_i),
    .io_ve_i(array_13_io_ve_i),
    .io_vf_i(array_13_io_vf_i),
    .io_vv_i(array_13_io_vv_i),
    .io_e_o(array_13_io_e_o),
    .io_f_o(array_13_io_f_o),
    .io_v_o(array_13_io_v_o)
  );
  SWCell array_14 ( // @[SWChisel.scala 170:39]
    .io_q(array_14_io_q),
    .io_r(array_14_io_r),
    .io_e_i(array_14_io_e_i),
    .io_f_i(array_14_io_f_i),
    .io_ve_i(array_14_io_ve_i),
    .io_vf_i(array_14_io_vf_i),
    .io_vv_i(array_14_io_vv_i),
    .io_e_o(array_14_io_e_o),
    .io_f_o(array_14_io_f_o),
    .io_v_o(array_14_io_v_o)
  );
  SWCell array_15 ( // @[SWChisel.scala 170:39]
    .io_q(array_15_io_q),
    .io_r(array_15_io_r),
    .io_e_i(array_15_io_e_i),
    .io_f_i(array_15_io_f_i),
    .io_ve_i(array_15_io_ve_i),
    .io_vf_i(array_15_io_vf_i),
    .io_vv_i(array_15_io_vv_i),
    .io_e_o(array_15_io_e_o),
    .io_f_o(array_15_io_f_o),
    .io_v_o(array_15_io_v_o)
  );
  SWCell array_16 ( // @[SWChisel.scala 170:39]
    .io_q(array_16_io_q),
    .io_r(array_16_io_r),
    .io_e_i(array_16_io_e_i),
    .io_f_i(array_16_io_f_i),
    .io_ve_i(array_16_io_ve_i),
    .io_vf_i(array_16_io_vf_i),
    .io_vv_i(array_16_io_vv_i),
    .io_e_o(array_16_io_e_o),
    .io_f_o(array_16_io_f_o),
    .io_v_o(array_16_io_v_o)
  );
  SWCell array_17 ( // @[SWChisel.scala 170:39]
    .io_q(array_17_io_q),
    .io_r(array_17_io_r),
    .io_e_i(array_17_io_e_i),
    .io_f_i(array_17_io_f_i),
    .io_ve_i(array_17_io_ve_i),
    .io_vf_i(array_17_io_vf_i),
    .io_vv_i(array_17_io_vv_i),
    .io_e_o(array_17_io_e_o),
    .io_f_o(array_17_io_f_o),
    .io_v_o(array_17_io_v_o)
  );
  SWCell array_18 ( // @[SWChisel.scala 170:39]
    .io_q(array_18_io_q),
    .io_r(array_18_io_r),
    .io_e_i(array_18_io_e_i),
    .io_f_i(array_18_io_f_i),
    .io_ve_i(array_18_io_ve_i),
    .io_vf_i(array_18_io_vf_i),
    .io_vv_i(array_18_io_vv_i),
    .io_e_o(array_18_io_e_o),
    .io_f_o(array_18_io_f_o),
    .io_v_o(array_18_io_v_o)
  );
  SWCell array_19 ( // @[SWChisel.scala 170:39]
    .io_q(array_19_io_q),
    .io_r(array_19_io_r),
    .io_e_i(array_19_io_e_i),
    .io_f_i(array_19_io_f_i),
    .io_ve_i(array_19_io_ve_i),
    .io_vf_i(array_19_io_vf_i),
    .io_vv_i(array_19_io_vv_i),
    .io_e_o(array_19_io_e_o),
    .io_f_o(array_19_io_f_o),
    .io_v_o(array_19_io_v_o)
  );
  SWCell array_20 ( // @[SWChisel.scala 170:39]
    .io_q(array_20_io_q),
    .io_r(array_20_io_r),
    .io_e_i(array_20_io_e_i),
    .io_f_i(array_20_io_f_i),
    .io_ve_i(array_20_io_ve_i),
    .io_vf_i(array_20_io_vf_i),
    .io_vv_i(array_20_io_vv_i),
    .io_e_o(array_20_io_e_o),
    .io_f_o(array_20_io_f_o),
    .io_v_o(array_20_io_v_o)
  );
  SWCell array_21 ( // @[SWChisel.scala 170:39]
    .io_q(array_21_io_q),
    .io_r(array_21_io_r),
    .io_e_i(array_21_io_e_i),
    .io_f_i(array_21_io_f_i),
    .io_ve_i(array_21_io_ve_i),
    .io_vf_i(array_21_io_vf_i),
    .io_vv_i(array_21_io_vv_i),
    .io_e_o(array_21_io_e_o),
    .io_f_o(array_21_io_f_o),
    .io_v_o(array_21_io_v_o)
  );
  SWCell array_22 ( // @[SWChisel.scala 170:39]
    .io_q(array_22_io_q),
    .io_r(array_22_io_r),
    .io_e_i(array_22_io_e_i),
    .io_f_i(array_22_io_f_i),
    .io_ve_i(array_22_io_ve_i),
    .io_vf_i(array_22_io_vf_i),
    .io_vv_i(array_22_io_vv_i),
    .io_e_o(array_22_io_e_o),
    .io_f_o(array_22_io_f_o),
    .io_v_o(array_22_io_v_o)
  );
  SWCell array_23 ( // @[SWChisel.scala 170:39]
    .io_q(array_23_io_q),
    .io_r(array_23_io_r),
    .io_e_i(array_23_io_e_i),
    .io_f_i(array_23_io_f_i),
    .io_ve_i(array_23_io_ve_i),
    .io_vf_i(array_23_io_vf_i),
    .io_vv_i(array_23_io_vv_i),
    .io_e_o(array_23_io_e_o),
    .io_f_o(array_23_io_f_o),
    .io_v_o(array_23_io_v_o)
  );
  SWCell array_24 ( // @[SWChisel.scala 170:39]
    .io_q(array_24_io_q),
    .io_r(array_24_io_r),
    .io_e_i(array_24_io_e_i),
    .io_f_i(array_24_io_f_i),
    .io_ve_i(array_24_io_ve_i),
    .io_vf_i(array_24_io_vf_i),
    .io_vv_i(array_24_io_vv_i),
    .io_e_o(array_24_io_e_o),
    .io_f_o(array_24_io_f_o),
    .io_v_o(array_24_io_v_o)
  );
  SWCell array_25 ( // @[SWChisel.scala 170:39]
    .io_q(array_25_io_q),
    .io_r(array_25_io_r),
    .io_e_i(array_25_io_e_i),
    .io_f_i(array_25_io_f_i),
    .io_ve_i(array_25_io_ve_i),
    .io_vf_i(array_25_io_vf_i),
    .io_vv_i(array_25_io_vv_i),
    .io_e_o(array_25_io_e_o),
    .io_f_o(array_25_io_f_o),
    .io_v_o(array_25_io_v_o)
  );
  SWCell array_26 ( // @[SWChisel.scala 170:39]
    .io_q(array_26_io_q),
    .io_r(array_26_io_r),
    .io_e_i(array_26_io_e_i),
    .io_f_i(array_26_io_f_i),
    .io_ve_i(array_26_io_ve_i),
    .io_vf_i(array_26_io_vf_i),
    .io_vv_i(array_26_io_vv_i),
    .io_e_o(array_26_io_e_o),
    .io_f_o(array_26_io_f_o),
    .io_v_o(array_26_io_v_o)
  );
  SWCell array_27 ( // @[SWChisel.scala 170:39]
    .io_q(array_27_io_q),
    .io_r(array_27_io_r),
    .io_e_i(array_27_io_e_i),
    .io_f_i(array_27_io_f_i),
    .io_ve_i(array_27_io_ve_i),
    .io_vf_i(array_27_io_vf_i),
    .io_vv_i(array_27_io_vv_i),
    .io_e_o(array_27_io_e_o),
    .io_f_o(array_27_io_f_o),
    .io_v_o(array_27_io_v_o)
  );
  SWCell array_28 ( // @[SWChisel.scala 170:39]
    .io_q(array_28_io_q),
    .io_r(array_28_io_r),
    .io_e_i(array_28_io_e_i),
    .io_f_i(array_28_io_f_i),
    .io_ve_i(array_28_io_ve_i),
    .io_vf_i(array_28_io_vf_i),
    .io_vv_i(array_28_io_vv_i),
    .io_e_o(array_28_io_e_o),
    .io_f_o(array_28_io_f_o),
    .io_v_o(array_28_io_v_o)
  );
  SWCell array_29 ( // @[SWChisel.scala 170:39]
    .io_q(array_29_io_q),
    .io_r(array_29_io_r),
    .io_e_i(array_29_io_e_i),
    .io_f_i(array_29_io_f_i),
    .io_ve_i(array_29_io_ve_i),
    .io_vf_i(array_29_io_vf_i),
    .io_vv_i(array_29_io_vv_i),
    .io_e_o(array_29_io_e_o),
    .io_f_o(array_29_io_f_o),
    .io_v_o(array_29_io_v_o)
  );
  MyCounter r_count_0 ( // @[SWChisel.scala 171:41]
    .clock(r_count_0_clock),
    .reset(r_count_0_reset),
    .io_en(r_count_0_io_en),
    .io_out(r_count_0_io_out)
  );
  MyCounter r_count_1 ( // @[SWChisel.scala 171:41]
    .clock(r_count_1_clock),
    .reset(r_count_1_reset),
    .io_en(r_count_1_io_en),
    .io_out(r_count_1_io_out)
  );
  MyCounter r_count_2 ( // @[SWChisel.scala 171:41]
    .clock(r_count_2_clock),
    .reset(r_count_2_reset),
    .io_en(r_count_2_io_en),
    .io_out(r_count_2_io_out)
  );
  MyCounter r_count_3 ( // @[SWChisel.scala 171:41]
    .clock(r_count_3_clock),
    .reset(r_count_3_reset),
    .io_en(r_count_3_io_en),
    .io_out(r_count_3_io_out)
  );
  MyCounter r_count_4 ( // @[SWChisel.scala 171:41]
    .clock(r_count_4_clock),
    .reset(r_count_4_reset),
    .io_en(r_count_4_io_en),
    .io_out(r_count_4_io_out)
  );
  MyCounter r_count_5 ( // @[SWChisel.scala 171:41]
    .clock(r_count_5_clock),
    .reset(r_count_5_reset),
    .io_en(r_count_5_io_en),
    .io_out(r_count_5_io_out)
  );
  MyCounter r_count_6 ( // @[SWChisel.scala 171:41]
    .clock(r_count_6_clock),
    .reset(r_count_6_reset),
    .io_en(r_count_6_io_en),
    .io_out(r_count_6_io_out)
  );
  MyCounter r_count_7 ( // @[SWChisel.scala 171:41]
    .clock(r_count_7_clock),
    .reset(r_count_7_reset),
    .io_en(r_count_7_io_en),
    .io_out(r_count_7_io_out)
  );
  MyCounter r_count_8 ( // @[SWChisel.scala 171:41]
    .clock(r_count_8_clock),
    .reset(r_count_8_reset),
    .io_en(r_count_8_io_en),
    .io_out(r_count_8_io_out)
  );
  MyCounter r_count_9 ( // @[SWChisel.scala 171:41]
    .clock(r_count_9_clock),
    .reset(r_count_9_reset),
    .io_en(r_count_9_io_en),
    .io_out(r_count_9_io_out)
  );
  MyCounter r_count_10 ( // @[SWChisel.scala 171:41]
    .clock(r_count_10_clock),
    .reset(r_count_10_reset),
    .io_en(r_count_10_io_en),
    .io_out(r_count_10_io_out)
  );
  MyCounter r_count_11 ( // @[SWChisel.scala 171:41]
    .clock(r_count_11_clock),
    .reset(r_count_11_reset),
    .io_en(r_count_11_io_en),
    .io_out(r_count_11_io_out)
  );
  MyCounter r_count_12 ( // @[SWChisel.scala 171:41]
    .clock(r_count_12_clock),
    .reset(r_count_12_reset),
    .io_en(r_count_12_io_en),
    .io_out(r_count_12_io_out)
  );
  MyCounter r_count_13 ( // @[SWChisel.scala 171:41]
    .clock(r_count_13_clock),
    .reset(r_count_13_reset),
    .io_en(r_count_13_io_en),
    .io_out(r_count_13_io_out)
  );
  MyCounter r_count_14 ( // @[SWChisel.scala 171:41]
    .clock(r_count_14_clock),
    .reset(r_count_14_reset),
    .io_en(r_count_14_io_en),
    .io_out(r_count_14_io_out)
  );
  MyCounter r_count_15 ( // @[SWChisel.scala 171:41]
    .clock(r_count_15_clock),
    .reset(r_count_15_reset),
    .io_en(r_count_15_io_en),
    .io_out(r_count_15_io_out)
  );
  MyCounter r_count_16 ( // @[SWChisel.scala 171:41]
    .clock(r_count_16_clock),
    .reset(r_count_16_reset),
    .io_en(r_count_16_io_en),
    .io_out(r_count_16_io_out)
  );
  MyCounter r_count_17 ( // @[SWChisel.scala 171:41]
    .clock(r_count_17_clock),
    .reset(r_count_17_reset),
    .io_en(r_count_17_io_en),
    .io_out(r_count_17_io_out)
  );
  MyCounter r_count_18 ( // @[SWChisel.scala 171:41]
    .clock(r_count_18_clock),
    .reset(r_count_18_reset),
    .io_en(r_count_18_io_en),
    .io_out(r_count_18_io_out)
  );
  MyCounter r_count_19 ( // @[SWChisel.scala 171:41]
    .clock(r_count_19_clock),
    .reset(r_count_19_reset),
    .io_en(r_count_19_io_en),
    .io_out(r_count_19_io_out)
  );
  MyCounter r_count_20 ( // @[SWChisel.scala 171:41]
    .clock(r_count_20_clock),
    .reset(r_count_20_reset),
    .io_en(r_count_20_io_en),
    .io_out(r_count_20_io_out)
  );
  MyCounter r_count_21 ( // @[SWChisel.scala 171:41]
    .clock(r_count_21_clock),
    .reset(r_count_21_reset),
    .io_en(r_count_21_io_en),
    .io_out(r_count_21_io_out)
  );
  MyCounter r_count_22 ( // @[SWChisel.scala 171:41]
    .clock(r_count_22_clock),
    .reset(r_count_22_reset),
    .io_en(r_count_22_io_en),
    .io_out(r_count_22_io_out)
  );
  MyCounter r_count_23 ( // @[SWChisel.scala 171:41]
    .clock(r_count_23_clock),
    .reset(r_count_23_reset),
    .io_en(r_count_23_io_en),
    .io_out(r_count_23_io_out)
  );
  MyCounter r_count_24 ( // @[SWChisel.scala 171:41]
    .clock(r_count_24_clock),
    .reset(r_count_24_reset),
    .io_en(r_count_24_io_en),
    .io_out(r_count_24_io_out)
  );
  MyCounter r_count_25 ( // @[SWChisel.scala 171:41]
    .clock(r_count_25_clock),
    .reset(r_count_25_reset),
    .io_en(r_count_25_io_en),
    .io_out(r_count_25_io_out)
  );
  MyCounter r_count_26 ( // @[SWChisel.scala 171:41]
    .clock(r_count_26_clock),
    .reset(r_count_26_reset),
    .io_en(r_count_26_io_en),
    .io_out(r_count_26_io_out)
  );
  MyCounter r_count_27 ( // @[SWChisel.scala 171:41]
    .clock(r_count_27_clock),
    .reset(r_count_27_reset),
    .io_en(r_count_27_io_en),
    .io_out(r_count_27_io_out)
  );
  MyCounter r_count_28 ( // @[SWChisel.scala 171:41]
    .clock(r_count_28_clock),
    .reset(r_count_28_reset),
    .io_en(r_count_28_io_en),
    .io_out(r_count_28_io_out)
  );
  MyCounter r_count_29 ( // @[SWChisel.scala 171:41]
    .clock(r_count_29_clock),
    .reset(r_count_29_reset),
    .io_en(r_count_29_io_en),
    .io_out(r_count_29_io_out)
  );
  MAX max ( // @[SWChisel.scala 174:19]
    .clock(max_clock),
    .reset(max_reset),
    .io_start(max_io_start),
    .io_in(max_io_in),
    .io_done(max_io_done),
    .io_out(max_io_out)
  );
  assign io_result = max_io_out; // @[SWChisel.scala 181:13]
  assign io_done = max_io_done; // @[SWChisel.scala 182:11]
  assign array_0_io_q = io_q_0_b; // @[SWChisel.scala 220:19]
  assign array_0_io_r = 10'h2ed == r_count_0_io_out ? io_r_749_b : _GEN_838; // @[SWChisel.scala 221:{19,19}]
  assign array_0_io_e_i = E_0; // @[SWChisel.scala 196:21]
  assign array_0_io_f_i = 16'sh0; // @[SWChisel.scala 198:21]
  assign array_0_io_ve_i = V1_1; // @[SWChisel.scala 197:22]
  assign array_0_io_vf_i = V1_0; // @[SWChisel.scala 199:22]
  assign array_0_io_vv_i = V2_0; // @[SWChisel.scala 200:22]
  assign array_1_io_q = io_q_1_b; // @[SWChisel.scala 220:19]
  assign array_1_io_r = 10'h2ed == r_count_1_io_out ? io_r_749_b : _GEN_1588; // @[SWChisel.scala 221:{19,19}]
  assign array_1_io_e_i = E_1; // @[SWChisel.scala 196:21]
  assign array_1_io_f_i = F_1; // @[SWChisel.scala 198:21]
  assign array_1_io_ve_i = V1_2; // @[SWChisel.scala 197:22]
  assign array_1_io_vf_i = V1_1; // @[SWChisel.scala 199:22]
  assign array_1_io_vv_i = V2_1; // @[SWChisel.scala 200:22]
  assign array_2_io_q = io_q_2_b; // @[SWChisel.scala 220:19]
  assign array_2_io_r = 10'h2ed == r_count_2_io_out ? io_r_749_b : _GEN_2338; // @[SWChisel.scala 221:{19,19}]
  assign array_2_io_e_i = E_2; // @[SWChisel.scala 196:21]
  assign array_2_io_f_i = F_2; // @[SWChisel.scala 198:21]
  assign array_2_io_ve_i = V1_3; // @[SWChisel.scala 197:22]
  assign array_2_io_vf_i = V1_2; // @[SWChisel.scala 199:22]
  assign array_2_io_vv_i = V2_2; // @[SWChisel.scala 200:22]
  assign array_3_io_q = io_q_3_b; // @[SWChisel.scala 220:19]
  assign array_3_io_r = 10'h2ed == r_count_3_io_out ? io_r_749_b : _GEN_3088; // @[SWChisel.scala 221:{19,19}]
  assign array_3_io_e_i = E_3; // @[SWChisel.scala 196:21]
  assign array_3_io_f_i = F_3; // @[SWChisel.scala 198:21]
  assign array_3_io_ve_i = V1_4; // @[SWChisel.scala 197:22]
  assign array_3_io_vf_i = V1_3; // @[SWChisel.scala 199:22]
  assign array_3_io_vv_i = V2_3; // @[SWChisel.scala 200:22]
  assign array_4_io_q = io_q_4_b; // @[SWChisel.scala 220:19]
  assign array_4_io_r = 10'h2ed == r_count_4_io_out ? io_r_749_b : _GEN_3838; // @[SWChisel.scala 221:{19,19}]
  assign array_4_io_e_i = E_4; // @[SWChisel.scala 196:21]
  assign array_4_io_f_i = F_4; // @[SWChisel.scala 198:21]
  assign array_4_io_ve_i = V1_5; // @[SWChisel.scala 197:22]
  assign array_4_io_vf_i = V1_4; // @[SWChisel.scala 199:22]
  assign array_4_io_vv_i = V2_4; // @[SWChisel.scala 200:22]
  assign array_5_io_q = io_q_5_b; // @[SWChisel.scala 220:19]
  assign array_5_io_r = 10'h2ed == r_count_5_io_out ? io_r_749_b : _GEN_4588; // @[SWChisel.scala 221:{19,19}]
  assign array_5_io_e_i = E_5; // @[SWChisel.scala 196:21]
  assign array_5_io_f_i = F_5; // @[SWChisel.scala 198:21]
  assign array_5_io_ve_i = V1_6; // @[SWChisel.scala 197:22]
  assign array_5_io_vf_i = V1_5; // @[SWChisel.scala 199:22]
  assign array_5_io_vv_i = V2_5; // @[SWChisel.scala 200:22]
  assign array_6_io_q = io_q_6_b; // @[SWChisel.scala 220:19]
  assign array_6_io_r = 10'h2ed == r_count_6_io_out ? io_r_749_b : _GEN_5338; // @[SWChisel.scala 221:{19,19}]
  assign array_6_io_e_i = E_6; // @[SWChisel.scala 196:21]
  assign array_6_io_f_i = F_6; // @[SWChisel.scala 198:21]
  assign array_6_io_ve_i = V1_7; // @[SWChisel.scala 197:22]
  assign array_6_io_vf_i = V1_6; // @[SWChisel.scala 199:22]
  assign array_6_io_vv_i = V2_6; // @[SWChisel.scala 200:22]
  assign array_7_io_q = io_q_7_b; // @[SWChisel.scala 220:19]
  assign array_7_io_r = 10'h2ed == r_count_7_io_out ? io_r_749_b : _GEN_6088; // @[SWChisel.scala 221:{19,19}]
  assign array_7_io_e_i = E_7; // @[SWChisel.scala 196:21]
  assign array_7_io_f_i = F_7; // @[SWChisel.scala 198:21]
  assign array_7_io_ve_i = V1_8; // @[SWChisel.scala 197:22]
  assign array_7_io_vf_i = V1_7; // @[SWChisel.scala 199:22]
  assign array_7_io_vv_i = V2_7; // @[SWChisel.scala 200:22]
  assign array_8_io_q = io_q_8_b; // @[SWChisel.scala 220:19]
  assign array_8_io_r = 10'h2ed == r_count_8_io_out ? io_r_749_b : _GEN_6838; // @[SWChisel.scala 221:{19,19}]
  assign array_8_io_e_i = E_8; // @[SWChisel.scala 196:21]
  assign array_8_io_f_i = F_8; // @[SWChisel.scala 198:21]
  assign array_8_io_ve_i = V1_9; // @[SWChisel.scala 197:22]
  assign array_8_io_vf_i = V1_8; // @[SWChisel.scala 199:22]
  assign array_8_io_vv_i = V2_8; // @[SWChisel.scala 200:22]
  assign array_9_io_q = io_q_9_b; // @[SWChisel.scala 220:19]
  assign array_9_io_r = 10'h2ed == r_count_9_io_out ? io_r_749_b : _GEN_7588; // @[SWChisel.scala 221:{19,19}]
  assign array_9_io_e_i = E_9; // @[SWChisel.scala 196:21]
  assign array_9_io_f_i = F_9; // @[SWChisel.scala 198:21]
  assign array_9_io_ve_i = V1_10; // @[SWChisel.scala 197:22]
  assign array_9_io_vf_i = V1_9; // @[SWChisel.scala 199:22]
  assign array_9_io_vv_i = V2_9; // @[SWChisel.scala 200:22]
  assign array_10_io_q = io_q_10_b; // @[SWChisel.scala 220:19]
  assign array_10_io_r = 10'h2ed == r_count_10_io_out ? io_r_749_b : _GEN_8338; // @[SWChisel.scala 221:{19,19}]
  assign array_10_io_e_i = E_10; // @[SWChisel.scala 196:21]
  assign array_10_io_f_i = F_10; // @[SWChisel.scala 198:21]
  assign array_10_io_ve_i = V1_11; // @[SWChisel.scala 197:22]
  assign array_10_io_vf_i = V1_10; // @[SWChisel.scala 199:22]
  assign array_10_io_vv_i = V2_10; // @[SWChisel.scala 200:22]
  assign array_11_io_q = io_q_11_b; // @[SWChisel.scala 220:19]
  assign array_11_io_r = 10'h2ed == r_count_11_io_out ? io_r_749_b : _GEN_9088; // @[SWChisel.scala 221:{19,19}]
  assign array_11_io_e_i = E_11; // @[SWChisel.scala 196:21]
  assign array_11_io_f_i = F_11; // @[SWChisel.scala 198:21]
  assign array_11_io_ve_i = V1_12; // @[SWChisel.scala 197:22]
  assign array_11_io_vf_i = V1_11; // @[SWChisel.scala 199:22]
  assign array_11_io_vv_i = V2_11; // @[SWChisel.scala 200:22]
  assign array_12_io_q = io_q_12_b; // @[SWChisel.scala 220:19]
  assign array_12_io_r = 10'h2ed == r_count_12_io_out ? io_r_749_b : _GEN_9838; // @[SWChisel.scala 221:{19,19}]
  assign array_12_io_e_i = E_12; // @[SWChisel.scala 196:21]
  assign array_12_io_f_i = F_12; // @[SWChisel.scala 198:21]
  assign array_12_io_ve_i = V1_13; // @[SWChisel.scala 197:22]
  assign array_12_io_vf_i = V1_12; // @[SWChisel.scala 199:22]
  assign array_12_io_vv_i = V2_12; // @[SWChisel.scala 200:22]
  assign array_13_io_q = io_q_13_b; // @[SWChisel.scala 220:19]
  assign array_13_io_r = 10'h2ed == r_count_13_io_out ? io_r_749_b : _GEN_10588; // @[SWChisel.scala 221:{19,19}]
  assign array_13_io_e_i = E_13; // @[SWChisel.scala 196:21]
  assign array_13_io_f_i = F_13; // @[SWChisel.scala 198:21]
  assign array_13_io_ve_i = V1_14; // @[SWChisel.scala 197:22]
  assign array_13_io_vf_i = V1_13; // @[SWChisel.scala 199:22]
  assign array_13_io_vv_i = V2_13; // @[SWChisel.scala 200:22]
  assign array_14_io_q = io_q_14_b; // @[SWChisel.scala 220:19]
  assign array_14_io_r = 10'h2ed == r_count_14_io_out ? io_r_749_b : _GEN_11338; // @[SWChisel.scala 221:{19,19}]
  assign array_14_io_e_i = E_14; // @[SWChisel.scala 196:21]
  assign array_14_io_f_i = F_14; // @[SWChisel.scala 198:21]
  assign array_14_io_ve_i = V1_15; // @[SWChisel.scala 197:22]
  assign array_14_io_vf_i = V1_14; // @[SWChisel.scala 199:22]
  assign array_14_io_vv_i = V2_14; // @[SWChisel.scala 200:22]
  assign array_15_io_q = io_q_15_b; // @[SWChisel.scala 220:19]
  assign array_15_io_r = 10'h2ed == r_count_15_io_out ? io_r_749_b : _GEN_12088; // @[SWChisel.scala 221:{19,19}]
  assign array_15_io_e_i = E_15; // @[SWChisel.scala 196:21]
  assign array_15_io_f_i = F_15; // @[SWChisel.scala 198:21]
  assign array_15_io_ve_i = V1_16; // @[SWChisel.scala 197:22]
  assign array_15_io_vf_i = V1_15; // @[SWChisel.scala 199:22]
  assign array_15_io_vv_i = V2_15; // @[SWChisel.scala 200:22]
  assign array_16_io_q = io_q_16_b; // @[SWChisel.scala 220:19]
  assign array_16_io_r = 10'h2ed == r_count_16_io_out ? io_r_749_b : _GEN_12838; // @[SWChisel.scala 221:{19,19}]
  assign array_16_io_e_i = E_16; // @[SWChisel.scala 196:21]
  assign array_16_io_f_i = F_16; // @[SWChisel.scala 198:21]
  assign array_16_io_ve_i = V1_17; // @[SWChisel.scala 197:22]
  assign array_16_io_vf_i = V1_16; // @[SWChisel.scala 199:22]
  assign array_16_io_vv_i = V2_16; // @[SWChisel.scala 200:22]
  assign array_17_io_q = io_q_17_b; // @[SWChisel.scala 220:19]
  assign array_17_io_r = 10'h2ed == r_count_17_io_out ? io_r_749_b : _GEN_13588; // @[SWChisel.scala 221:{19,19}]
  assign array_17_io_e_i = E_17; // @[SWChisel.scala 196:21]
  assign array_17_io_f_i = F_17; // @[SWChisel.scala 198:21]
  assign array_17_io_ve_i = V1_18; // @[SWChisel.scala 197:22]
  assign array_17_io_vf_i = V1_17; // @[SWChisel.scala 199:22]
  assign array_17_io_vv_i = V2_17; // @[SWChisel.scala 200:22]
  assign array_18_io_q = io_q_18_b; // @[SWChisel.scala 220:19]
  assign array_18_io_r = 10'h2ed == r_count_18_io_out ? io_r_749_b : _GEN_14338; // @[SWChisel.scala 221:{19,19}]
  assign array_18_io_e_i = E_18; // @[SWChisel.scala 196:21]
  assign array_18_io_f_i = F_18; // @[SWChisel.scala 198:21]
  assign array_18_io_ve_i = V1_19; // @[SWChisel.scala 197:22]
  assign array_18_io_vf_i = V1_18; // @[SWChisel.scala 199:22]
  assign array_18_io_vv_i = V2_18; // @[SWChisel.scala 200:22]
  assign array_19_io_q = io_q_19_b; // @[SWChisel.scala 220:19]
  assign array_19_io_r = 10'h2ed == r_count_19_io_out ? io_r_749_b : _GEN_15088; // @[SWChisel.scala 221:{19,19}]
  assign array_19_io_e_i = E_19; // @[SWChisel.scala 196:21]
  assign array_19_io_f_i = F_19; // @[SWChisel.scala 198:21]
  assign array_19_io_ve_i = V1_20; // @[SWChisel.scala 197:22]
  assign array_19_io_vf_i = V1_19; // @[SWChisel.scala 199:22]
  assign array_19_io_vv_i = V2_19; // @[SWChisel.scala 200:22]
  assign array_20_io_q = io_q_20_b; // @[SWChisel.scala 220:19]
  assign array_20_io_r = 10'h2ed == r_count_20_io_out ? io_r_749_b : _GEN_15838; // @[SWChisel.scala 221:{19,19}]
  assign array_20_io_e_i = E_20; // @[SWChisel.scala 196:21]
  assign array_20_io_f_i = F_20; // @[SWChisel.scala 198:21]
  assign array_20_io_ve_i = V1_21; // @[SWChisel.scala 197:22]
  assign array_20_io_vf_i = V1_20; // @[SWChisel.scala 199:22]
  assign array_20_io_vv_i = V2_20; // @[SWChisel.scala 200:22]
  assign array_21_io_q = io_q_21_b; // @[SWChisel.scala 220:19]
  assign array_21_io_r = 10'h2ed == r_count_21_io_out ? io_r_749_b : _GEN_16588; // @[SWChisel.scala 221:{19,19}]
  assign array_21_io_e_i = E_21; // @[SWChisel.scala 196:21]
  assign array_21_io_f_i = F_21; // @[SWChisel.scala 198:21]
  assign array_21_io_ve_i = V1_22; // @[SWChisel.scala 197:22]
  assign array_21_io_vf_i = V1_21; // @[SWChisel.scala 199:22]
  assign array_21_io_vv_i = V2_21; // @[SWChisel.scala 200:22]
  assign array_22_io_q = io_q_22_b; // @[SWChisel.scala 220:19]
  assign array_22_io_r = 10'h2ed == r_count_22_io_out ? io_r_749_b : _GEN_17338; // @[SWChisel.scala 221:{19,19}]
  assign array_22_io_e_i = E_22; // @[SWChisel.scala 196:21]
  assign array_22_io_f_i = F_22; // @[SWChisel.scala 198:21]
  assign array_22_io_ve_i = V1_23; // @[SWChisel.scala 197:22]
  assign array_22_io_vf_i = V1_22; // @[SWChisel.scala 199:22]
  assign array_22_io_vv_i = V2_22; // @[SWChisel.scala 200:22]
  assign array_23_io_q = io_q_23_b; // @[SWChisel.scala 220:19]
  assign array_23_io_r = 10'h2ed == r_count_23_io_out ? io_r_749_b : _GEN_18088; // @[SWChisel.scala 221:{19,19}]
  assign array_23_io_e_i = E_23; // @[SWChisel.scala 196:21]
  assign array_23_io_f_i = F_23; // @[SWChisel.scala 198:21]
  assign array_23_io_ve_i = V1_24; // @[SWChisel.scala 197:22]
  assign array_23_io_vf_i = V1_23; // @[SWChisel.scala 199:22]
  assign array_23_io_vv_i = V2_23; // @[SWChisel.scala 200:22]
  assign array_24_io_q = io_q_24_b; // @[SWChisel.scala 220:19]
  assign array_24_io_r = 10'h2ed == r_count_24_io_out ? io_r_749_b : _GEN_18838; // @[SWChisel.scala 221:{19,19}]
  assign array_24_io_e_i = E_24; // @[SWChisel.scala 196:21]
  assign array_24_io_f_i = F_24; // @[SWChisel.scala 198:21]
  assign array_24_io_ve_i = V1_25; // @[SWChisel.scala 197:22]
  assign array_24_io_vf_i = V1_24; // @[SWChisel.scala 199:22]
  assign array_24_io_vv_i = V2_24; // @[SWChisel.scala 200:22]
  assign array_25_io_q = io_q_25_b; // @[SWChisel.scala 220:19]
  assign array_25_io_r = 10'h2ed == r_count_25_io_out ? io_r_749_b : _GEN_19588; // @[SWChisel.scala 221:{19,19}]
  assign array_25_io_e_i = E_25; // @[SWChisel.scala 196:21]
  assign array_25_io_f_i = F_25; // @[SWChisel.scala 198:21]
  assign array_25_io_ve_i = V1_26; // @[SWChisel.scala 197:22]
  assign array_25_io_vf_i = V1_25; // @[SWChisel.scala 199:22]
  assign array_25_io_vv_i = V2_25; // @[SWChisel.scala 200:22]
  assign array_26_io_q = io_q_26_b; // @[SWChisel.scala 220:19]
  assign array_26_io_r = 10'h2ed == r_count_26_io_out ? io_r_749_b : _GEN_20338; // @[SWChisel.scala 221:{19,19}]
  assign array_26_io_e_i = E_26; // @[SWChisel.scala 196:21]
  assign array_26_io_f_i = F_26; // @[SWChisel.scala 198:21]
  assign array_26_io_ve_i = V1_27; // @[SWChisel.scala 197:22]
  assign array_26_io_vf_i = V1_26; // @[SWChisel.scala 199:22]
  assign array_26_io_vv_i = V2_26; // @[SWChisel.scala 200:22]
  assign array_27_io_q = io_q_27_b; // @[SWChisel.scala 220:19]
  assign array_27_io_r = 10'h2ed == r_count_27_io_out ? io_r_749_b : _GEN_21088; // @[SWChisel.scala 221:{19,19}]
  assign array_27_io_e_i = E_27; // @[SWChisel.scala 196:21]
  assign array_27_io_f_i = F_27; // @[SWChisel.scala 198:21]
  assign array_27_io_ve_i = V1_28; // @[SWChisel.scala 197:22]
  assign array_27_io_vf_i = V1_27; // @[SWChisel.scala 199:22]
  assign array_27_io_vv_i = V2_27; // @[SWChisel.scala 200:22]
  assign array_28_io_q = io_q_28_b; // @[SWChisel.scala 220:19]
  assign array_28_io_r = 10'h2ed == r_count_28_io_out ? io_r_749_b : _GEN_21838; // @[SWChisel.scala 221:{19,19}]
  assign array_28_io_e_i = E_28; // @[SWChisel.scala 196:21]
  assign array_28_io_f_i = F_28; // @[SWChisel.scala 198:21]
  assign array_28_io_ve_i = V1_29; // @[SWChisel.scala 197:22]
  assign array_28_io_vf_i = V1_28; // @[SWChisel.scala 199:22]
  assign array_28_io_vv_i = V2_28; // @[SWChisel.scala 200:22]
  assign array_29_io_q = io_q_29_b; // @[SWChisel.scala 220:19]
  assign array_29_io_r = 10'h2ed == r_count_29_io_out ? io_r_749_b : _GEN_22588; // @[SWChisel.scala 221:{19,19}]
  assign array_29_io_e_i = E_29; // @[SWChisel.scala 196:21]
  assign array_29_io_f_i = F_29; // @[SWChisel.scala 198:21]
  assign array_29_io_ve_i = V1_30; // @[SWChisel.scala 197:22]
  assign array_29_io_vf_i = V1_29; // @[SWChisel.scala 199:22]
  assign array_29_io_vv_i = V2_29; // @[SWChisel.scala 200:22]
  assign r_count_0_clock = clock;
  assign r_count_0_reset = reset;
  assign r_count_0_io_en = start_reg_0; // @[SWChisel.scala 192:22]
  assign r_count_1_clock = clock;
  assign r_count_1_reset = reset;
  assign r_count_1_io_en = start_reg_1; // @[SWChisel.scala 192:22]
  assign r_count_2_clock = clock;
  assign r_count_2_reset = reset;
  assign r_count_2_io_en = start_reg_2; // @[SWChisel.scala 192:22]
  assign r_count_3_clock = clock;
  assign r_count_3_reset = reset;
  assign r_count_3_io_en = start_reg_3; // @[SWChisel.scala 192:22]
  assign r_count_4_clock = clock;
  assign r_count_4_reset = reset;
  assign r_count_4_io_en = start_reg_4; // @[SWChisel.scala 192:22]
  assign r_count_5_clock = clock;
  assign r_count_5_reset = reset;
  assign r_count_5_io_en = start_reg_5; // @[SWChisel.scala 192:22]
  assign r_count_6_clock = clock;
  assign r_count_6_reset = reset;
  assign r_count_6_io_en = start_reg_6; // @[SWChisel.scala 192:22]
  assign r_count_7_clock = clock;
  assign r_count_7_reset = reset;
  assign r_count_7_io_en = start_reg_7; // @[SWChisel.scala 192:22]
  assign r_count_8_clock = clock;
  assign r_count_8_reset = reset;
  assign r_count_8_io_en = start_reg_8; // @[SWChisel.scala 192:22]
  assign r_count_9_clock = clock;
  assign r_count_9_reset = reset;
  assign r_count_9_io_en = start_reg_9; // @[SWChisel.scala 192:22]
  assign r_count_10_clock = clock;
  assign r_count_10_reset = reset;
  assign r_count_10_io_en = start_reg_10; // @[SWChisel.scala 192:22]
  assign r_count_11_clock = clock;
  assign r_count_11_reset = reset;
  assign r_count_11_io_en = start_reg_11; // @[SWChisel.scala 192:22]
  assign r_count_12_clock = clock;
  assign r_count_12_reset = reset;
  assign r_count_12_io_en = start_reg_12; // @[SWChisel.scala 192:22]
  assign r_count_13_clock = clock;
  assign r_count_13_reset = reset;
  assign r_count_13_io_en = start_reg_13; // @[SWChisel.scala 192:22]
  assign r_count_14_clock = clock;
  assign r_count_14_reset = reset;
  assign r_count_14_io_en = start_reg_14; // @[SWChisel.scala 192:22]
  assign r_count_15_clock = clock;
  assign r_count_15_reset = reset;
  assign r_count_15_io_en = start_reg_15; // @[SWChisel.scala 192:22]
  assign r_count_16_clock = clock;
  assign r_count_16_reset = reset;
  assign r_count_16_io_en = start_reg_16; // @[SWChisel.scala 192:22]
  assign r_count_17_clock = clock;
  assign r_count_17_reset = reset;
  assign r_count_17_io_en = start_reg_17; // @[SWChisel.scala 192:22]
  assign r_count_18_clock = clock;
  assign r_count_18_reset = reset;
  assign r_count_18_io_en = start_reg_18; // @[SWChisel.scala 192:22]
  assign r_count_19_clock = clock;
  assign r_count_19_reset = reset;
  assign r_count_19_io_en = start_reg_19; // @[SWChisel.scala 192:22]
  assign r_count_20_clock = clock;
  assign r_count_20_reset = reset;
  assign r_count_20_io_en = start_reg_20; // @[SWChisel.scala 192:22]
  assign r_count_21_clock = clock;
  assign r_count_21_reset = reset;
  assign r_count_21_io_en = start_reg_21; // @[SWChisel.scala 192:22]
  assign r_count_22_clock = clock;
  assign r_count_22_reset = reset;
  assign r_count_22_io_en = start_reg_22; // @[SWChisel.scala 192:22]
  assign r_count_23_clock = clock;
  assign r_count_23_reset = reset;
  assign r_count_23_io_en = start_reg_23; // @[SWChisel.scala 192:22]
  assign r_count_24_clock = clock;
  assign r_count_24_reset = reset;
  assign r_count_24_io_en = start_reg_24; // @[SWChisel.scala 192:22]
  assign r_count_25_clock = clock;
  assign r_count_25_reset = reset;
  assign r_count_25_io_en = start_reg_25; // @[SWChisel.scala 192:22]
  assign r_count_26_clock = clock;
  assign r_count_26_reset = reset;
  assign r_count_26_io_en = start_reg_26; // @[SWChisel.scala 192:22]
  assign r_count_27_clock = clock;
  assign r_count_27_reset = reset;
  assign r_count_27_io_en = start_reg_27; // @[SWChisel.scala 192:22]
  assign r_count_28_clock = clock;
  assign r_count_28_reset = reset;
  assign r_count_28_io_en = start_reg_28; // @[SWChisel.scala 192:22]
  assign r_count_29_clock = clock;
  assign r_count_29_reset = reset;
  assign r_count_29_io_en = start_reg_29; // @[SWChisel.scala 192:22]
  assign max_clock = clock;
  assign max_reset = reset;
  assign max_io_start = start_reg_29; // @[SWChisel.scala 178:16]
  assign max_io_in = V1_30; // @[SWChisel.scala 177:13]
  always @(posedge clock) begin
    if (reset) begin // @[SWChisel.scala 162:18]
      E_0 <= -16'sh2; // @[SWChisel.scala 162:18]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      E_0 <= array_0_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_1 <= -16'sh3; // @[SWChisel.scala 162:18]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      E_1 <= array_1_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_2 <= -16'sh4; // @[SWChisel.scala 162:18]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      E_2 <= array_2_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_3 <= -16'sh5; // @[SWChisel.scala 162:18]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      E_3 <= array_3_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_4 <= -16'sh6; // @[SWChisel.scala 162:18]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      E_4 <= array_4_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_5 <= -16'sh7; // @[SWChisel.scala 162:18]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      E_5 <= array_5_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_6 <= -16'sh8; // @[SWChisel.scala 162:18]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      E_6 <= array_6_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_7 <= -16'sh9; // @[SWChisel.scala 162:18]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      E_7 <= array_7_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_8 <= -16'sha; // @[SWChisel.scala 162:18]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      E_8 <= array_8_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_9 <= -16'shb; // @[SWChisel.scala 162:18]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      E_9 <= array_9_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_10 <= -16'shc; // @[SWChisel.scala 162:18]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      E_10 <= array_10_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_11 <= -16'shd; // @[SWChisel.scala 162:18]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      E_11 <= array_11_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_12 <= -16'she; // @[SWChisel.scala 162:18]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      E_12 <= array_12_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_13 <= -16'shf; // @[SWChisel.scala 162:18]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      E_13 <= array_13_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_14 <= -16'sh10; // @[SWChisel.scala 162:18]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      E_14 <= array_14_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_15 <= -16'sh11; // @[SWChisel.scala 162:18]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      E_15 <= array_15_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_16 <= -16'sh12; // @[SWChisel.scala 162:18]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      E_16 <= array_16_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_17 <= -16'sh13; // @[SWChisel.scala 162:18]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      E_17 <= array_17_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_18 <= -16'sh14; // @[SWChisel.scala 162:18]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      E_18 <= array_18_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_19 <= -16'sh15; // @[SWChisel.scala 162:18]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      E_19 <= array_19_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_20 <= -16'sh16; // @[SWChisel.scala 162:18]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      E_20 <= array_20_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_21 <= -16'sh17; // @[SWChisel.scala 162:18]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      E_21 <= array_21_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_22 <= -16'sh18; // @[SWChisel.scala 162:18]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      E_22 <= array_22_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_23 <= -16'sh19; // @[SWChisel.scala 162:18]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      E_23 <= array_23_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_24 <= -16'sh1a; // @[SWChisel.scala 162:18]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      E_24 <= array_24_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_25 <= -16'sh1b; // @[SWChisel.scala 162:18]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      E_25 <= array_25_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_26 <= -16'sh1c; // @[SWChisel.scala 162:18]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      E_26 <= array_26_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_27 <= -16'sh1d; // @[SWChisel.scala 162:18]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      E_27 <= array_27_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_28 <= -16'sh1e; // @[SWChisel.scala 162:18]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      E_28 <= array_28_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_29 <= -16'sh1f; // @[SWChisel.scala 162:18]
    end else if (start_reg_29) begin // @[SWChisel.scala 207:25]
      E_29 <= array_29_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_1 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      F_1 <= array_0_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_2 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      F_2 <= array_1_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_3 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      F_3 <= array_2_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_4 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      F_4 <= array_3_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_5 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      F_5 <= array_4_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_6 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      F_6 <= array_5_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_7 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      F_7 <= array_6_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_8 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      F_8 <= array_7_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_9 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      F_9 <= array_8_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_10 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      F_10 <= array_9_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_11 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      F_11 <= array_10_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_12 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      F_12 <= array_11_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_13 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      F_13 <= array_12_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_14 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      F_14 <= array_13_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_15 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      F_15 <= array_14_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_16 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      F_16 <= array_15_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_17 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      F_17 <= array_16_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_18 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      F_18 <= array_17_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_19 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      F_19 <= array_18_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_20 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      F_20 <= array_19_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_21 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      F_21 <= array_20_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_22 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      F_22 <= array_21_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_23 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      F_23 <= array_22_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_24 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      F_24 <= array_23_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_25 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      F_25 <= array_24_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_26 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      F_26 <= array_25_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_27 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      F_27 <= array_26_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_28 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      F_28 <= array_27_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_29 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      F_29 <= array_28_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_0 <= -16'sh1; // @[SWChisel.scala 164:19]
    end else begin
      V1_0 <= 16'sh0; // @[SWChisel.scala 165:9]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_1 <= -16'sh2; // @[SWChisel.scala 164:19]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      V1_1 <= array_0_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_2 <= -16'sh3; // @[SWChisel.scala 164:19]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      V1_2 <= array_1_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_3 <= -16'sh4; // @[SWChisel.scala 164:19]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      V1_3 <= array_2_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_4 <= -16'sh5; // @[SWChisel.scala 164:19]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      V1_4 <= array_3_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_5 <= -16'sh6; // @[SWChisel.scala 164:19]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      V1_5 <= array_4_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_6 <= -16'sh7; // @[SWChisel.scala 164:19]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      V1_6 <= array_5_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_7 <= -16'sh8; // @[SWChisel.scala 164:19]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      V1_7 <= array_6_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_8 <= -16'sh9; // @[SWChisel.scala 164:19]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      V1_8 <= array_7_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_9 <= -16'sha; // @[SWChisel.scala 164:19]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      V1_9 <= array_8_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_10 <= -16'shb; // @[SWChisel.scala 164:19]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      V1_10 <= array_9_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_11 <= -16'shc; // @[SWChisel.scala 164:19]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      V1_11 <= array_10_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_12 <= -16'shd; // @[SWChisel.scala 164:19]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      V1_12 <= array_11_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_13 <= -16'she; // @[SWChisel.scala 164:19]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      V1_13 <= array_12_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_14 <= -16'shf; // @[SWChisel.scala 164:19]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      V1_14 <= array_13_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_15 <= -16'sh10; // @[SWChisel.scala 164:19]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      V1_15 <= array_14_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_16 <= -16'sh11; // @[SWChisel.scala 164:19]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      V1_16 <= array_15_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_17 <= -16'sh12; // @[SWChisel.scala 164:19]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      V1_17 <= array_16_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_18 <= -16'sh13; // @[SWChisel.scala 164:19]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      V1_18 <= array_17_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_19 <= -16'sh14; // @[SWChisel.scala 164:19]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      V1_19 <= array_18_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_20 <= -16'sh15; // @[SWChisel.scala 164:19]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      V1_20 <= array_19_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_21 <= -16'sh16; // @[SWChisel.scala 164:19]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      V1_21 <= array_20_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_22 <= -16'sh17; // @[SWChisel.scala 164:19]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      V1_22 <= array_21_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_23 <= -16'sh18; // @[SWChisel.scala 164:19]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      V1_23 <= array_22_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_24 <= -16'sh19; // @[SWChisel.scala 164:19]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      V1_24 <= array_23_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_25 <= -16'sh1a; // @[SWChisel.scala 164:19]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      V1_25 <= array_24_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_26 <= -16'sh1b; // @[SWChisel.scala 164:19]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      V1_26 <= array_25_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_27 <= -16'sh1c; // @[SWChisel.scala 164:19]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      V1_27 <= array_26_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_28 <= -16'sh1d; // @[SWChisel.scala 164:19]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      V1_28 <= array_27_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_29 <= -16'sh1e; // @[SWChisel.scala 164:19]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      V1_29 <= array_28_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_30 <= -16'sh1f; // @[SWChisel.scala 164:19]
    end else if (start_reg_29) begin // @[SWChisel.scala 207:25]
      V1_30 <= array_29_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_0 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_0 <= V1_0; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_1 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_1 <= V1_1; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_2 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_2 <= V1_2; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_3 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_3 <= V1_3; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_4 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_4 <= V1_4; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_5 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_5 <= V1_5; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_6 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_6 <= V1_6; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_7 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_7 <= V1_7; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_8 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_8 <= V1_8; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_9 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_9 <= V1_9; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_10 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_10 <= V1_10; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_11 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_11 <= V1_11; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_12 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_12 <= V1_12; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_13 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_13 <= V1_13; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_14 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_14 <= V1_14; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_15 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_15 <= V1_15; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_16 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_16 <= V1_16; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_17 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_17 <= V1_17; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_18 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_18 <= V1_18; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_19 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_19 <= V1_19; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_20 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_20 <= V1_20; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_21 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_21 <= V1_21; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_22 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_22 <= V1_22; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_23 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_23 <= V1_23; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_24 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_24 <= V1_24; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_25 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_25 <= V1_25; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_26 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_26 <= V1_26; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_27 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_27 <= V1_27; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_28 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_28 <= V1_28; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_29 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_29 <= V1_29; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_0 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_0 <= io_start; // @[SWChisel.scala 185:16]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_1 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_1 <= start_reg_0; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_2 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_2 <= start_reg_1; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_3 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_3 <= start_reg_2; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_4 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_4 <= start_reg_3; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_5 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_5 <= start_reg_4; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_6 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_6 <= start_reg_5; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_7 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_7 <= start_reg_6; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_8 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_8 <= start_reg_7; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_9 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_9 <= start_reg_8; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_10 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_10 <= start_reg_9; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_11 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_11 <= start_reg_10; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_12 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_12 <= start_reg_11; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_13 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_13 <= start_reg_12; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_14 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_14 <= start_reg_13; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_15 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_15 <= start_reg_14; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_16 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_16 <= start_reg_15; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_17 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_17 <= start_reg_16; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_18 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_18 <= start_reg_17; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_19 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_19 <= start_reg_18; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_20 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_20 <= start_reg_19; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_21 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_21 <= start_reg_20; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_22 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_22 <= start_reg_21; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_23 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_23 <= start_reg_22; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_24 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_24 <= start_reg_23; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_25 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_25 <= start_reg_24; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_26 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_26 <= start_reg_25; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_27 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_27 <= start_reg_26; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_28 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_28 <= start_reg_27; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_29 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_29 <= start_reg_28; // @[SWChisel.scala 187:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  E_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  E_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  E_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  E_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  E_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  E_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  E_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  E_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  E_8 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  E_9 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  E_10 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  E_11 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  E_12 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  E_13 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  E_14 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  E_15 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  E_16 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  E_17 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  E_18 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  E_19 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  E_20 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  E_21 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  E_22 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  E_23 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  E_24 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  E_25 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  E_26 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  E_27 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  E_28 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  E_29 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  F_1 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  F_2 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  F_3 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  F_4 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  F_5 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  F_6 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  F_7 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  F_8 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  F_9 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  F_10 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  F_11 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  F_12 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  F_13 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  F_14 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  F_15 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  F_16 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  F_17 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  F_18 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  F_19 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  F_20 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  F_21 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  F_22 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  F_23 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  F_24 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  F_25 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  F_26 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  F_27 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  F_28 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  F_29 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  V1_0 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  V1_1 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  V1_2 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  V1_3 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  V1_4 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  V1_5 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  V1_6 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  V1_7 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  V1_8 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  V1_9 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  V1_10 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  V1_11 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  V1_12 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  V1_13 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  V1_14 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  V1_15 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  V1_16 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  V1_17 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  V1_18 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  V1_19 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  V1_20 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  V1_21 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  V1_22 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  V1_23 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  V1_24 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  V1_25 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  V1_26 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  V1_27 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  V1_28 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  V1_29 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  V1_30 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  V2_0 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  V2_1 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  V2_2 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  V2_3 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  V2_4 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  V2_5 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  V2_6 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  V2_7 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  V2_8 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  V2_9 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  V2_10 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  V2_11 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  V2_12 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  V2_13 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  V2_14 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  V2_15 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  V2_16 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  V2_17 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  V2_18 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  V2_19 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  V2_20 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  V2_21 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  V2_22 = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  V2_23 = _RAND_113[15:0];
  _RAND_114 = {1{`RANDOM}};
  V2_24 = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  V2_25 = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  V2_26 = _RAND_116[15:0];
  _RAND_117 = {1{`RANDOM}};
  V2_27 = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  V2_28 = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  V2_29 = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  start_reg_0 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  start_reg_1 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  start_reg_2 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  start_reg_3 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  start_reg_4 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  start_reg_5 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  start_reg_6 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  start_reg_7 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  start_reg_8 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  start_reg_9 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  start_reg_10 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  start_reg_11 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  start_reg_12 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  start_reg_13 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  start_reg_14 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  start_reg_15 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  start_reg_16 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  start_reg_17 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  start_reg_18 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  start_reg_19 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  start_reg_20 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  start_reg_21 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  start_reg_22 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  start_reg_23 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  start_reg_24 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  start_reg_25 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  start_reg_26 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  start_reg_27 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  start_reg_28 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  start_reg_29 = _RAND_149[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
