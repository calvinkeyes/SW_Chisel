module SWCell(
  input  [1:0]  io_q,
  input  [1:0]  io_r,
  input  [15:0] io_e_i,
  input  [15:0] io_f_i,
  input  [15:0] io_ve_i,
  input  [15:0] io_vf_i,
  input  [15:0] io_vv_i,
  output [15:0] io_e_o,
  output [15:0] io_f_o,
  output [15:0] io_v_o
);
  wire [15:0] _T_2 = $signed(io_ve_i) - 16'sh2; // @[SWChisel.scala 78:17]
  wire [15:0] _T_5 = $signed(io_e_i) - 16'sh1; // @[SWChisel.scala 78:39]
  wire [15:0] e_max = $signed(_T_2) >= $signed(_T_5) ? $signed(_T_2) : $signed(_T_5); // @[SWChisel.scala 78:51 79:11 81:11]
  wire [15:0] _T_9 = $signed(io_vf_i) - 16'sh2; // @[SWChisel.scala 85:17]
  wire [15:0] _T_12 = $signed(io_f_i) - 16'sh1; // @[SWChisel.scala 85:38]
  wire [15:0] f_max = $signed(_T_9) > $signed(_T_12) ? $signed(_T_9) : $signed(_T_12); // @[SWChisel.scala 85:50 86:11 88:11]
  wire [15:0] ef_temp = $signed(e_max) > $signed(f_max) ? $signed(e_max) : $signed(f_max); // @[SWChisel.scala 92:24 93:13 95:13]
  wire [15:0] _v_temp_T_2 = $signed(io_vv_i) + 16'sh2; // @[SWChisel.scala 100:23]
  wire [15:0] _v_temp_T_5 = $signed(io_vv_i) - 16'sh2; // @[SWChisel.scala 102:23]
  wire [15:0] v_temp = io_q == io_r ? $signed(_v_temp_T_2) : $signed(_v_temp_T_5); // @[SWChisel.scala 100:12 102:12 99:24]
  assign io_e_o = $signed(_T_2) >= $signed(_T_5) ? $signed(_T_2) : $signed(_T_5); // @[SWChisel.scala 78:51 79:11 81:11]
  assign io_f_o = $signed(_T_9) > $signed(_T_12) ? $signed(_T_9) : $signed(_T_12); // @[SWChisel.scala 85:50 86:11 88:11]
  assign io_v_o = $signed(v_temp) > $signed(ef_temp) ? $signed(v_temp) : $signed(ef_temp); // @[SWChisel.scala 106:27 107:11 109:11]
endmodule
module MyCounter(
  input        clock,
  input        reset,
  input        io_en,
  output [7:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] _io_out_T_2 = io_out + 8'h1; // @[SWChisel.scala 155:55]
  reg [7:0] io_out_r; // @[Reg.scala 35:20]
  assign io_out = io_out_r; // @[SWChisel.scala 155:12]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      io_out_r <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_out < 8'hc8) begin // @[SWChisel.scala 155:28]
        io_out_r <= _io_out_T_2;
      end else begin
        io_out_r <= 8'h0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_out_r = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MAX(
  input         clock,
  input         reset,
  input         io_start,
  input  [15:0] io_in,
  output        io_done,
  output [15:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] max; // @[SWChisel.scala 122:20]
  reg [7:0] counter; // @[SWChisel.scala 133:24]
  wire [7:0] _counter_T_1 = counter - 8'h1; // @[SWChisel.scala 135:24]
  assign io_done = counter == 8'h0; // @[SWChisel.scala 141:17]
  assign io_out = max; // @[SWChisel.scala 123:10]
  always @(posedge clock) begin
    if (reset) begin // @[SWChisel.scala 122:20]
      max <= 16'sh8000; // @[SWChisel.scala 122:20]
    end else if ($signed(io_in) > $signed(max)) begin // @[SWChisel.scala 126:22]
      max <= io_in; // @[SWChisel.scala 127:9]
    end
    if (reset) begin // @[SWChisel.scala 133:24]
      counter <= 8'hc9; // @[SWChisel.scala 133:24]
    end else if (counter == 8'h0) begin // @[SWChisel.scala 141:26]
      counter <= 8'h0; // @[SWChisel.scala 143:13]
    end else if (io_start) begin // @[SWChisel.scala 134:19]
      counter <= _counter_T_1; // @[SWChisel.scala 135:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  max = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  counter = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SW(
  input         clock,
  input         reset,
  input  [1:0]  io_q_0_b,
  input  [1:0]  io_q_1_b,
  input  [1:0]  io_q_2_b,
  input  [1:0]  io_q_3_b,
  input  [1:0]  io_q_4_b,
  input  [1:0]  io_q_5_b,
  input  [1:0]  io_q_6_b,
  input  [1:0]  io_q_7_b,
  input  [1:0]  io_q_8_b,
  input  [1:0]  io_q_9_b,
  input  [1:0]  io_q_10_b,
  input  [1:0]  io_q_11_b,
  input  [1:0]  io_q_12_b,
  input  [1:0]  io_q_13_b,
  input  [1:0]  io_q_14_b,
  input  [1:0]  io_q_15_b,
  input  [1:0]  io_q_16_b,
  input  [1:0]  io_q_17_b,
  input  [1:0]  io_q_18_b,
  input  [1:0]  io_q_19_b,
  input  [1:0]  io_q_20_b,
  input  [1:0]  io_q_21_b,
  input  [1:0]  io_q_22_b,
  input  [1:0]  io_q_23_b,
  input  [1:0]  io_q_24_b,
  input  [1:0]  io_q_25_b,
  input  [1:0]  io_q_26_b,
  input  [1:0]  io_q_27_b,
  input  [1:0]  io_q_28_b,
  input  [1:0]  io_q_29_b,
  input  [1:0]  io_q_30_b,
  input  [1:0]  io_q_31_b,
  input  [1:0]  io_q_32_b,
  input  [1:0]  io_q_33_b,
  input  [1:0]  io_q_34_b,
  input  [1:0]  io_q_35_b,
  input  [1:0]  io_q_36_b,
  input  [1:0]  io_q_37_b,
  input  [1:0]  io_q_38_b,
  input  [1:0]  io_q_39_b,
  input  [1:0]  io_q_40_b,
  input  [1:0]  io_q_41_b,
  input  [1:0]  io_q_42_b,
  input  [1:0]  io_q_43_b,
  input  [1:0]  io_q_44_b,
  input  [1:0]  io_q_45_b,
  input  [1:0]  io_q_46_b,
  input  [1:0]  io_q_47_b,
  input  [1:0]  io_q_48_b,
  input  [1:0]  io_q_49_b,
  input  [1:0]  io_q_50_b,
  input  [1:0]  io_q_51_b,
  input  [1:0]  io_q_52_b,
  input  [1:0]  io_q_53_b,
  input  [1:0]  io_q_54_b,
  input  [1:0]  io_q_55_b,
  input  [1:0]  io_q_56_b,
  input  [1:0]  io_q_57_b,
  input  [1:0]  io_q_58_b,
  input  [1:0]  io_q_59_b,
  input  [1:0]  io_q_60_b,
  input  [1:0]  io_q_61_b,
  input  [1:0]  io_q_62_b,
  input  [1:0]  io_q_63_b,
  input  [1:0]  io_q_64_b,
  input  [1:0]  io_q_65_b,
  input  [1:0]  io_q_66_b,
  input  [1:0]  io_q_67_b,
  input  [1:0]  io_q_68_b,
  input  [1:0]  io_q_69_b,
  input  [1:0]  io_q_70_b,
  input  [1:0]  io_q_71_b,
  input  [1:0]  io_q_72_b,
  input  [1:0]  io_q_73_b,
  input  [1:0]  io_q_74_b,
  input  [1:0]  io_q_75_b,
  input  [1:0]  io_q_76_b,
  input  [1:0]  io_q_77_b,
  input  [1:0]  io_q_78_b,
  input  [1:0]  io_q_79_b,
  input  [1:0]  io_q_80_b,
  input  [1:0]  io_q_81_b,
  input  [1:0]  io_q_82_b,
  input  [1:0]  io_q_83_b,
  input  [1:0]  io_q_84_b,
  input  [1:0]  io_q_85_b,
  input  [1:0]  io_q_86_b,
  input  [1:0]  io_q_87_b,
  input  [1:0]  io_q_88_b,
  input  [1:0]  io_q_89_b,
  input  [1:0]  io_q_90_b,
  input  [1:0]  io_q_91_b,
  input  [1:0]  io_q_92_b,
  input  [1:0]  io_q_93_b,
  input  [1:0]  io_q_94_b,
  input  [1:0]  io_q_95_b,
  input  [1:0]  io_q_96_b,
  input  [1:0]  io_q_97_b,
  input  [1:0]  io_q_98_b,
  input  [1:0]  io_q_99_b,
  input  [1:0]  io_r_0_b,
  input  [1:0]  io_r_1_b,
  input  [1:0]  io_r_2_b,
  input  [1:0]  io_r_3_b,
  input  [1:0]  io_r_4_b,
  input  [1:0]  io_r_5_b,
  input  [1:0]  io_r_6_b,
  input  [1:0]  io_r_7_b,
  input  [1:0]  io_r_8_b,
  input  [1:0]  io_r_9_b,
  input  [1:0]  io_r_10_b,
  input  [1:0]  io_r_11_b,
  input  [1:0]  io_r_12_b,
  input  [1:0]  io_r_13_b,
  input  [1:0]  io_r_14_b,
  input  [1:0]  io_r_15_b,
  input  [1:0]  io_r_16_b,
  input  [1:0]  io_r_17_b,
  input  [1:0]  io_r_18_b,
  input  [1:0]  io_r_19_b,
  input  [1:0]  io_r_20_b,
  input  [1:0]  io_r_21_b,
  input  [1:0]  io_r_22_b,
  input  [1:0]  io_r_23_b,
  input  [1:0]  io_r_24_b,
  input  [1:0]  io_r_25_b,
  input  [1:0]  io_r_26_b,
  input  [1:0]  io_r_27_b,
  input  [1:0]  io_r_28_b,
  input  [1:0]  io_r_29_b,
  input  [1:0]  io_r_30_b,
  input  [1:0]  io_r_31_b,
  input  [1:0]  io_r_32_b,
  input  [1:0]  io_r_33_b,
  input  [1:0]  io_r_34_b,
  input  [1:0]  io_r_35_b,
  input  [1:0]  io_r_36_b,
  input  [1:0]  io_r_37_b,
  input  [1:0]  io_r_38_b,
  input  [1:0]  io_r_39_b,
  input  [1:0]  io_r_40_b,
  input  [1:0]  io_r_41_b,
  input  [1:0]  io_r_42_b,
  input  [1:0]  io_r_43_b,
  input  [1:0]  io_r_44_b,
  input  [1:0]  io_r_45_b,
  input  [1:0]  io_r_46_b,
  input  [1:0]  io_r_47_b,
  input  [1:0]  io_r_48_b,
  input  [1:0]  io_r_49_b,
  input  [1:0]  io_r_50_b,
  input  [1:0]  io_r_51_b,
  input  [1:0]  io_r_52_b,
  input  [1:0]  io_r_53_b,
  input  [1:0]  io_r_54_b,
  input  [1:0]  io_r_55_b,
  input  [1:0]  io_r_56_b,
  input  [1:0]  io_r_57_b,
  input  [1:0]  io_r_58_b,
  input  [1:0]  io_r_59_b,
  input  [1:0]  io_r_60_b,
  input  [1:0]  io_r_61_b,
  input  [1:0]  io_r_62_b,
  input  [1:0]  io_r_63_b,
  input  [1:0]  io_r_64_b,
  input  [1:0]  io_r_65_b,
  input  [1:0]  io_r_66_b,
  input  [1:0]  io_r_67_b,
  input  [1:0]  io_r_68_b,
  input  [1:0]  io_r_69_b,
  input  [1:0]  io_r_70_b,
  input  [1:0]  io_r_71_b,
  input  [1:0]  io_r_72_b,
  input  [1:0]  io_r_73_b,
  input  [1:0]  io_r_74_b,
  input  [1:0]  io_r_75_b,
  input  [1:0]  io_r_76_b,
  input  [1:0]  io_r_77_b,
  input  [1:0]  io_r_78_b,
  input  [1:0]  io_r_79_b,
  input  [1:0]  io_r_80_b,
  input  [1:0]  io_r_81_b,
  input  [1:0]  io_r_82_b,
  input  [1:0]  io_r_83_b,
  input  [1:0]  io_r_84_b,
  input  [1:0]  io_r_85_b,
  input  [1:0]  io_r_86_b,
  input  [1:0]  io_r_87_b,
  input  [1:0]  io_r_88_b,
  input  [1:0]  io_r_89_b,
  input  [1:0]  io_r_90_b,
  input  [1:0]  io_r_91_b,
  input  [1:0]  io_r_92_b,
  input  [1:0]  io_r_93_b,
  input  [1:0]  io_r_94_b,
  input  [1:0]  io_r_95_b,
  input  [1:0]  io_r_96_b,
  input  [1:0]  io_r_97_b,
  input  [1:0]  io_r_98_b,
  input  [1:0]  io_r_99_b,
  input  [1:0]  io_r_100_b,
  input  [1:0]  io_r_101_b,
  input  [1:0]  io_r_102_b,
  input  [1:0]  io_r_103_b,
  input  [1:0]  io_r_104_b,
  input  [1:0]  io_r_105_b,
  input  [1:0]  io_r_106_b,
  input  [1:0]  io_r_107_b,
  input  [1:0]  io_r_108_b,
  input  [1:0]  io_r_109_b,
  input  [1:0]  io_r_110_b,
  input  [1:0]  io_r_111_b,
  input  [1:0]  io_r_112_b,
  input  [1:0]  io_r_113_b,
  input  [1:0]  io_r_114_b,
  input  [1:0]  io_r_115_b,
  input  [1:0]  io_r_116_b,
  input  [1:0]  io_r_117_b,
  input  [1:0]  io_r_118_b,
  input  [1:0]  io_r_119_b,
  input  [1:0]  io_r_120_b,
  input  [1:0]  io_r_121_b,
  input  [1:0]  io_r_122_b,
  input  [1:0]  io_r_123_b,
  input  [1:0]  io_r_124_b,
  input  [1:0]  io_r_125_b,
  input  [1:0]  io_r_126_b,
  input  [1:0]  io_r_127_b,
  input  [1:0]  io_r_128_b,
  input  [1:0]  io_r_129_b,
  input  [1:0]  io_r_130_b,
  input  [1:0]  io_r_131_b,
  input  [1:0]  io_r_132_b,
  input  [1:0]  io_r_133_b,
  input  [1:0]  io_r_134_b,
  input  [1:0]  io_r_135_b,
  input  [1:0]  io_r_136_b,
  input  [1:0]  io_r_137_b,
  input  [1:0]  io_r_138_b,
  input  [1:0]  io_r_139_b,
  input  [1:0]  io_r_140_b,
  input  [1:0]  io_r_141_b,
  input  [1:0]  io_r_142_b,
  input  [1:0]  io_r_143_b,
  input  [1:0]  io_r_144_b,
  input  [1:0]  io_r_145_b,
  input  [1:0]  io_r_146_b,
  input  [1:0]  io_r_147_b,
  input  [1:0]  io_r_148_b,
  input  [1:0]  io_r_149_b,
  input  [1:0]  io_r_150_b,
  input  [1:0]  io_r_151_b,
  input  [1:0]  io_r_152_b,
  input  [1:0]  io_r_153_b,
  input  [1:0]  io_r_154_b,
  input  [1:0]  io_r_155_b,
  input  [1:0]  io_r_156_b,
  input  [1:0]  io_r_157_b,
  input  [1:0]  io_r_158_b,
  input  [1:0]  io_r_159_b,
  input  [1:0]  io_r_160_b,
  input  [1:0]  io_r_161_b,
  input  [1:0]  io_r_162_b,
  input  [1:0]  io_r_163_b,
  input  [1:0]  io_r_164_b,
  input  [1:0]  io_r_165_b,
  input  [1:0]  io_r_166_b,
  input  [1:0]  io_r_167_b,
  input  [1:0]  io_r_168_b,
  input  [1:0]  io_r_169_b,
  input  [1:0]  io_r_170_b,
  input  [1:0]  io_r_171_b,
  input  [1:0]  io_r_172_b,
  input  [1:0]  io_r_173_b,
  input  [1:0]  io_r_174_b,
  input  [1:0]  io_r_175_b,
  input  [1:0]  io_r_176_b,
  input  [1:0]  io_r_177_b,
  input  [1:0]  io_r_178_b,
  input  [1:0]  io_r_179_b,
  input  [1:0]  io_r_180_b,
  input  [1:0]  io_r_181_b,
  input  [1:0]  io_r_182_b,
  input  [1:0]  io_r_183_b,
  input  [1:0]  io_r_184_b,
  input  [1:0]  io_r_185_b,
  input  [1:0]  io_r_186_b,
  input  [1:0]  io_r_187_b,
  input  [1:0]  io_r_188_b,
  input  [1:0]  io_r_189_b,
  input  [1:0]  io_r_190_b,
  input  [1:0]  io_r_191_b,
  input  [1:0]  io_r_192_b,
  input  [1:0]  io_r_193_b,
  input  [1:0]  io_r_194_b,
  input  [1:0]  io_r_195_b,
  input  [1:0]  io_r_196_b,
  input  [1:0]  io_r_197_b,
  input  [1:0]  io_r_198_b,
  input  [1:0]  io_r_199_b,
  input         io_start,
  output [15:0] io_result,
  output        io_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
`endif // RANDOMIZE_REG_INIT
  wire [1:0] array_0_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_0_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_1_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_1_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_2_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_2_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_3_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_3_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_4_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_4_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_5_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_5_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_6_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_6_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_7_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_7_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_8_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_8_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_9_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_9_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_10_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_10_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_11_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_11_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_12_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_12_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_13_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_13_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_14_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_14_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_15_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_15_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_16_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_16_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_17_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_17_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_18_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_18_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_19_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_19_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_20_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_20_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_21_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_21_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_22_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_22_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_23_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_23_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_24_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_24_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_25_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_25_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_26_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_26_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_27_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_27_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_28_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_28_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_29_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_29_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_30_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_30_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_31_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_31_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_32_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_32_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_33_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_33_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_34_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_34_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_35_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_35_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_36_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_36_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_37_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_37_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_38_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_38_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_39_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_39_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_40_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_40_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_41_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_41_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_42_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_42_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_43_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_43_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_44_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_44_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_45_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_45_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_46_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_46_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_47_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_47_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_48_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_48_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_49_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_49_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_50_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_50_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_50_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_50_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_50_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_50_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_50_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_50_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_50_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_50_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_51_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_51_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_51_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_51_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_51_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_51_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_51_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_51_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_51_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_51_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_52_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_52_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_52_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_52_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_52_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_52_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_52_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_52_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_52_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_52_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_53_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_53_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_53_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_53_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_53_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_53_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_53_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_53_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_53_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_53_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_54_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_54_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_54_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_54_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_54_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_54_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_54_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_54_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_54_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_54_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_55_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_55_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_55_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_55_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_55_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_55_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_55_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_55_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_55_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_55_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_56_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_56_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_56_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_56_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_56_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_56_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_56_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_56_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_56_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_56_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_57_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_57_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_57_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_57_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_57_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_57_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_57_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_57_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_57_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_57_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_58_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_58_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_58_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_58_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_58_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_58_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_58_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_58_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_58_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_58_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_59_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_59_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_59_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_59_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_59_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_59_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_59_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_59_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_59_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_59_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_60_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_60_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_60_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_60_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_60_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_60_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_60_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_60_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_60_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_60_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_61_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_61_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_61_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_61_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_61_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_61_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_61_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_61_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_61_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_61_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_62_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_62_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_62_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_62_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_62_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_62_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_62_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_62_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_62_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_62_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_63_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_63_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_63_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_63_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_63_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_63_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_63_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_63_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_63_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_63_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_64_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_64_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_64_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_64_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_64_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_64_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_64_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_64_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_64_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_64_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_65_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_65_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_65_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_65_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_65_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_65_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_65_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_65_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_65_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_65_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_66_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_66_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_66_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_66_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_66_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_66_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_66_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_66_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_66_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_66_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_67_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_67_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_67_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_67_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_67_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_67_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_67_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_67_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_67_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_67_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_68_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_68_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_68_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_68_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_68_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_68_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_68_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_68_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_68_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_68_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_69_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_69_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_69_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_69_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_69_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_69_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_69_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_69_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_69_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_69_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_70_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_70_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_70_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_70_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_70_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_70_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_70_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_70_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_70_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_70_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_71_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_71_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_71_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_71_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_71_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_71_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_71_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_71_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_71_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_71_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_72_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_72_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_72_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_72_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_72_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_72_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_72_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_72_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_72_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_72_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_73_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_73_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_73_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_73_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_73_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_73_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_73_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_73_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_73_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_73_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_74_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_74_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_74_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_74_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_74_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_74_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_74_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_74_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_74_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_74_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_75_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_75_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_75_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_75_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_75_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_75_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_75_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_75_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_75_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_75_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_76_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_76_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_76_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_76_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_76_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_76_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_76_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_76_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_76_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_76_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_77_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_77_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_77_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_77_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_77_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_77_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_77_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_77_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_77_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_77_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_78_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_78_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_78_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_78_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_78_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_78_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_78_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_78_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_78_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_78_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_79_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_79_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_79_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_79_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_79_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_79_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_79_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_79_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_79_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_79_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_80_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_80_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_80_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_80_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_80_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_80_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_80_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_80_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_80_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_80_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_81_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_81_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_81_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_81_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_81_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_81_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_81_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_81_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_81_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_81_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_82_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_82_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_82_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_82_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_82_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_82_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_82_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_82_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_82_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_82_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_83_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_83_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_83_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_83_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_83_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_83_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_83_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_83_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_83_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_83_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_84_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_84_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_84_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_84_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_84_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_84_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_84_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_84_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_84_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_84_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_85_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_85_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_85_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_85_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_85_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_85_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_85_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_85_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_85_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_85_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_86_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_86_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_86_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_86_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_86_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_86_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_86_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_86_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_86_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_86_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_87_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_87_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_87_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_87_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_87_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_87_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_87_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_87_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_87_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_87_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_88_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_88_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_88_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_88_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_88_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_88_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_88_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_88_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_88_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_88_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_89_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_89_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_89_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_89_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_89_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_89_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_89_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_89_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_89_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_89_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_90_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_90_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_90_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_90_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_90_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_90_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_90_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_90_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_90_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_90_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_91_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_91_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_91_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_91_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_91_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_91_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_91_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_91_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_91_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_91_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_92_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_92_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_92_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_92_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_92_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_92_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_92_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_92_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_92_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_92_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_93_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_93_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_93_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_93_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_93_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_93_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_93_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_93_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_93_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_93_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_94_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_94_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_94_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_94_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_94_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_94_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_94_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_94_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_94_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_94_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_95_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_95_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_95_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_95_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_95_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_95_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_95_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_95_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_95_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_95_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_96_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_96_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_96_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_96_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_96_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_96_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_96_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_96_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_96_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_96_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_97_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_97_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_97_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_97_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_97_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_97_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_97_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_97_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_97_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_97_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_98_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_98_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_98_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_98_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_98_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_98_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_98_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_98_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_98_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_98_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_99_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_99_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_99_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_99_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_99_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_99_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_99_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_99_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_99_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_99_io_v_o; // @[SWChisel.scala 170:39]
  wire  r_count_0_clock; // @[SWChisel.scala 171:41]
  wire  r_count_0_reset; // @[SWChisel.scala 171:41]
  wire  r_count_0_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_0_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_1_clock; // @[SWChisel.scala 171:41]
  wire  r_count_1_reset; // @[SWChisel.scala 171:41]
  wire  r_count_1_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_1_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_2_clock; // @[SWChisel.scala 171:41]
  wire  r_count_2_reset; // @[SWChisel.scala 171:41]
  wire  r_count_2_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_2_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_3_clock; // @[SWChisel.scala 171:41]
  wire  r_count_3_reset; // @[SWChisel.scala 171:41]
  wire  r_count_3_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_3_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_4_clock; // @[SWChisel.scala 171:41]
  wire  r_count_4_reset; // @[SWChisel.scala 171:41]
  wire  r_count_4_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_4_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_5_clock; // @[SWChisel.scala 171:41]
  wire  r_count_5_reset; // @[SWChisel.scala 171:41]
  wire  r_count_5_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_5_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_6_clock; // @[SWChisel.scala 171:41]
  wire  r_count_6_reset; // @[SWChisel.scala 171:41]
  wire  r_count_6_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_6_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_7_clock; // @[SWChisel.scala 171:41]
  wire  r_count_7_reset; // @[SWChisel.scala 171:41]
  wire  r_count_7_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_7_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_8_clock; // @[SWChisel.scala 171:41]
  wire  r_count_8_reset; // @[SWChisel.scala 171:41]
  wire  r_count_8_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_8_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_9_clock; // @[SWChisel.scala 171:41]
  wire  r_count_9_reset; // @[SWChisel.scala 171:41]
  wire  r_count_9_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_9_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_10_clock; // @[SWChisel.scala 171:41]
  wire  r_count_10_reset; // @[SWChisel.scala 171:41]
  wire  r_count_10_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_10_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_11_clock; // @[SWChisel.scala 171:41]
  wire  r_count_11_reset; // @[SWChisel.scala 171:41]
  wire  r_count_11_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_11_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_12_clock; // @[SWChisel.scala 171:41]
  wire  r_count_12_reset; // @[SWChisel.scala 171:41]
  wire  r_count_12_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_12_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_13_clock; // @[SWChisel.scala 171:41]
  wire  r_count_13_reset; // @[SWChisel.scala 171:41]
  wire  r_count_13_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_13_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_14_clock; // @[SWChisel.scala 171:41]
  wire  r_count_14_reset; // @[SWChisel.scala 171:41]
  wire  r_count_14_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_14_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_15_clock; // @[SWChisel.scala 171:41]
  wire  r_count_15_reset; // @[SWChisel.scala 171:41]
  wire  r_count_15_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_15_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_16_clock; // @[SWChisel.scala 171:41]
  wire  r_count_16_reset; // @[SWChisel.scala 171:41]
  wire  r_count_16_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_16_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_17_clock; // @[SWChisel.scala 171:41]
  wire  r_count_17_reset; // @[SWChisel.scala 171:41]
  wire  r_count_17_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_17_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_18_clock; // @[SWChisel.scala 171:41]
  wire  r_count_18_reset; // @[SWChisel.scala 171:41]
  wire  r_count_18_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_18_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_19_clock; // @[SWChisel.scala 171:41]
  wire  r_count_19_reset; // @[SWChisel.scala 171:41]
  wire  r_count_19_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_19_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_20_clock; // @[SWChisel.scala 171:41]
  wire  r_count_20_reset; // @[SWChisel.scala 171:41]
  wire  r_count_20_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_20_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_21_clock; // @[SWChisel.scala 171:41]
  wire  r_count_21_reset; // @[SWChisel.scala 171:41]
  wire  r_count_21_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_21_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_22_clock; // @[SWChisel.scala 171:41]
  wire  r_count_22_reset; // @[SWChisel.scala 171:41]
  wire  r_count_22_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_22_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_23_clock; // @[SWChisel.scala 171:41]
  wire  r_count_23_reset; // @[SWChisel.scala 171:41]
  wire  r_count_23_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_23_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_24_clock; // @[SWChisel.scala 171:41]
  wire  r_count_24_reset; // @[SWChisel.scala 171:41]
  wire  r_count_24_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_24_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_25_clock; // @[SWChisel.scala 171:41]
  wire  r_count_25_reset; // @[SWChisel.scala 171:41]
  wire  r_count_25_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_25_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_26_clock; // @[SWChisel.scala 171:41]
  wire  r_count_26_reset; // @[SWChisel.scala 171:41]
  wire  r_count_26_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_26_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_27_clock; // @[SWChisel.scala 171:41]
  wire  r_count_27_reset; // @[SWChisel.scala 171:41]
  wire  r_count_27_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_27_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_28_clock; // @[SWChisel.scala 171:41]
  wire  r_count_28_reset; // @[SWChisel.scala 171:41]
  wire  r_count_28_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_28_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_29_clock; // @[SWChisel.scala 171:41]
  wire  r_count_29_reset; // @[SWChisel.scala 171:41]
  wire  r_count_29_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_29_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_30_clock; // @[SWChisel.scala 171:41]
  wire  r_count_30_reset; // @[SWChisel.scala 171:41]
  wire  r_count_30_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_30_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_31_clock; // @[SWChisel.scala 171:41]
  wire  r_count_31_reset; // @[SWChisel.scala 171:41]
  wire  r_count_31_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_31_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_32_clock; // @[SWChisel.scala 171:41]
  wire  r_count_32_reset; // @[SWChisel.scala 171:41]
  wire  r_count_32_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_32_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_33_clock; // @[SWChisel.scala 171:41]
  wire  r_count_33_reset; // @[SWChisel.scala 171:41]
  wire  r_count_33_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_33_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_34_clock; // @[SWChisel.scala 171:41]
  wire  r_count_34_reset; // @[SWChisel.scala 171:41]
  wire  r_count_34_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_34_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_35_clock; // @[SWChisel.scala 171:41]
  wire  r_count_35_reset; // @[SWChisel.scala 171:41]
  wire  r_count_35_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_35_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_36_clock; // @[SWChisel.scala 171:41]
  wire  r_count_36_reset; // @[SWChisel.scala 171:41]
  wire  r_count_36_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_36_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_37_clock; // @[SWChisel.scala 171:41]
  wire  r_count_37_reset; // @[SWChisel.scala 171:41]
  wire  r_count_37_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_37_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_38_clock; // @[SWChisel.scala 171:41]
  wire  r_count_38_reset; // @[SWChisel.scala 171:41]
  wire  r_count_38_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_38_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_39_clock; // @[SWChisel.scala 171:41]
  wire  r_count_39_reset; // @[SWChisel.scala 171:41]
  wire  r_count_39_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_39_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_40_clock; // @[SWChisel.scala 171:41]
  wire  r_count_40_reset; // @[SWChisel.scala 171:41]
  wire  r_count_40_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_40_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_41_clock; // @[SWChisel.scala 171:41]
  wire  r_count_41_reset; // @[SWChisel.scala 171:41]
  wire  r_count_41_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_41_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_42_clock; // @[SWChisel.scala 171:41]
  wire  r_count_42_reset; // @[SWChisel.scala 171:41]
  wire  r_count_42_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_42_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_43_clock; // @[SWChisel.scala 171:41]
  wire  r_count_43_reset; // @[SWChisel.scala 171:41]
  wire  r_count_43_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_43_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_44_clock; // @[SWChisel.scala 171:41]
  wire  r_count_44_reset; // @[SWChisel.scala 171:41]
  wire  r_count_44_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_44_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_45_clock; // @[SWChisel.scala 171:41]
  wire  r_count_45_reset; // @[SWChisel.scala 171:41]
  wire  r_count_45_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_45_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_46_clock; // @[SWChisel.scala 171:41]
  wire  r_count_46_reset; // @[SWChisel.scala 171:41]
  wire  r_count_46_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_46_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_47_clock; // @[SWChisel.scala 171:41]
  wire  r_count_47_reset; // @[SWChisel.scala 171:41]
  wire  r_count_47_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_47_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_48_clock; // @[SWChisel.scala 171:41]
  wire  r_count_48_reset; // @[SWChisel.scala 171:41]
  wire  r_count_48_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_48_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_49_clock; // @[SWChisel.scala 171:41]
  wire  r_count_49_reset; // @[SWChisel.scala 171:41]
  wire  r_count_49_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_49_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_50_clock; // @[SWChisel.scala 171:41]
  wire  r_count_50_reset; // @[SWChisel.scala 171:41]
  wire  r_count_50_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_50_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_51_clock; // @[SWChisel.scala 171:41]
  wire  r_count_51_reset; // @[SWChisel.scala 171:41]
  wire  r_count_51_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_51_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_52_clock; // @[SWChisel.scala 171:41]
  wire  r_count_52_reset; // @[SWChisel.scala 171:41]
  wire  r_count_52_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_52_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_53_clock; // @[SWChisel.scala 171:41]
  wire  r_count_53_reset; // @[SWChisel.scala 171:41]
  wire  r_count_53_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_53_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_54_clock; // @[SWChisel.scala 171:41]
  wire  r_count_54_reset; // @[SWChisel.scala 171:41]
  wire  r_count_54_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_54_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_55_clock; // @[SWChisel.scala 171:41]
  wire  r_count_55_reset; // @[SWChisel.scala 171:41]
  wire  r_count_55_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_55_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_56_clock; // @[SWChisel.scala 171:41]
  wire  r_count_56_reset; // @[SWChisel.scala 171:41]
  wire  r_count_56_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_56_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_57_clock; // @[SWChisel.scala 171:41]
  wire  r_count_57_reset; // @[SWChisel.scala 171:41]
  wire  r_count_57_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_57_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_58_clock; // @[SWChisel.scala 171:41]
  wire  r_count_58_reset; // @[SWChisel.scala 171:41]
  wire  r_count_58_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_58_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_59_clock; // @[SWChisel.scala 171:41]
  wire  r_count_59_reset; // @[SWChisel.scala 171:41]
  wire  r_count_59_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_59_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_60_clock; // @[SWChisel.scala 171:41]
  wire  r_count_60_reset; // @[SWChisel.scala 171:41]
  wire  r_count_60_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_60_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_61_clock; // @[SWChisel.scala 171:41]
  wire  r_count_61_reset; // @[SWChisel.scala 171:41]
  wire  r_count_61_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_61_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_62_clock; // @[SWChisel.scala 171:41]
  wire  r_count_62_reset; // @[SWChisel.scala 171:41]
  wire  r_count_62_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_62_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_63_clock; // @[SWChisel.scala 171:41]
  wire  r_count_63_reset; // @[SWChisel.scala 171:41]
  wire  r_count_63_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_63_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_64_clock; // @[SWChisel.scala 171:41]
  wire  r_count_64_reset; // @[SWChisel.scala 171:41]
  wire  r_count_64_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_64_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_65_clock; // @[SWChisel.scala 171:41]
  wire  r_count_65_reset; // @[SWChisel.scala 171:41]
  wire  r_count_65_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_65_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_66_clock; // @[SWChisel.scala 171:41]
  wire  r_count_66_reset; // @[SWChisel.scala 171:41]
  wire  r_count_66_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_66_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_67_clock; // @[SWChisel.scala 171:41]
  wire  r_count_67_reset; // @[SWChisel.scala 171:41]
  wire  r_count_67_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_67_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_68_clock; // @[SWChisel.scala 171:41]
  wire  r_count_68_reset; // @[SWChisel.scala 171:41]
  wire  r_count_68_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_68_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_69_clock; // @[SWChisel.scala 171:41]
  wire  r_count_69_reset; // @[SWChisel.scala 171:41]
  wire  r_count_69_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_69_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_70_clock; // @[SWChisel.scala 171:41]
  wire  r_count_70_reset; // @[SWChisel.scala 171:41]
  wire  r_count_70_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_70_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_71_clock; // @[SWChisel.scala 171:41]
  wire  r_count_71_reset; // @[SWChisel.scala 171:41]
  wire  r_count_71_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_71_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_72_clock; // @[SWChisel.scala 171:41]
  wire  r_count_72_reset; // @[SWChisel.scala 171:41]
  wire  r_count_72_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_72_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_73_clock; // @[SWChisel.scala 171:41]
  wire  r_count_73_reset; // @[SWChisel.scala 171:41]
  wire  r_count_73_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_73_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_74_clock; // @[SWChisel.scala 171:41]
  wire  r_count_74_reset; // @[SWChisel.scala 171:41]
  wire  r_count_74_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_74_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_75_clock; // @[SWChisel.scala 171:41]
  wire  r_count_75_reset; // @[SWChisel.scala 171:41]
  wire  r_count_75_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_75_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_76_clock; // @[SWChisel.scala 171:41]
  wire  r_count_76_reset; // @[SWChisel.scala 171:41]
  wire  r_count_76_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_76_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_77_clock; // @[SWChisel.scala 171:41]
  wire  r_count_77_reset; // @[SWChisel.scala 171:41]
  wire  r_count_77_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_77_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_78_clock; // @[SWChisel.scala 171:41]
  wire  r_count_78_reset; // @[SWChisel.scala 171:41]
  wire  r_count_78_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_78_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_79_clock; // @[SWChisel.scala 171:41]
  wire  r_count_79_reset; // @[SWChisel.scala 171:41]
  wire  r_count_79_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_79_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_80_clock; // @[SWChisel.scala 171:41]
  wire  r_count_80_reset; // @[SWChisel.scala 171:41]
  wire  r_count_80_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_80_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_81_clock; // @[SWChisel.scala 171:41]
  wire  r_count_81_reset; // @[SWChisel.scala 171:41]
  wire  r_count_81_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_81_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_82_clock; // @[SWChisel.scala 171:41]
  wire  r_count_82_reset; // @[SWChisel.scala 171:41]
  wire  r_count_82_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_82_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_83_clock; // @[SWChisel.scala 171:41]
  wire  r_count_83_reset; // @[SWChisel.scala 171:41]
  wire  r_count_83_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_83_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_84_clock; // @[SWChisel.scala 171:41]
  wire  r_count_84_reset; // @[SWChisel.scala 171:41]
  wire  r_count_84_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_84_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_85_clock; // @[SWChisel.scala 171:41]
  wire  r_count_85_reset; // @[SWChisel.scala 171:41]
  wire  r_count_85_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_85_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_86_clock; // @[SWChisel.scala 171:41]
  wire  r_count_86_reset; // @[SWChisel.scala 171:41]
  wire  r_count_86_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_86_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_87_clock; // @[SWChisel.scala 171:41]
  wire  r_count_87_reset; // @[SWChisel.scala 171:41]
  wire  r_count_87_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_87_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_88_clock; // @[SWChisel.scala 171:41]
  wire  r_count_88_reset; // @[SWChisel.scala 171:41]
  wire  r_count_88_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_88_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_89_clock; // @[SWChisel.scala 171:41]
  wire  r_count_89_reset; // @[SWChisel.scala 171:41]
  wire  r_count_89_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_89_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_90_clock; // @[SWChisel.scala 171:41]
  wire  r_count_90_reset; // @[SWChisel.scala 171:41]
  wire  r_count_90_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_90_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_91_clock; // @[SWChisel.scala 171:41]
  wire  r_count_91_reset; // @[SWChisel.scala 171:41]
  wire  r_count_91_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_91_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_92_clock; // @[SWChisel.scala 171:41]
  wire  r_count_92_reset; // @[SWChisel.scala 171:41]
  wire  r_count_92_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_92_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_93_clock; // @[SWChisel.scala 171:41]
  wire  r_count_93_reset; // @[SWChisel.scala 171:41]
  wire  r_count_93_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_93_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_94_clock; // @[SWChisel.scala 171:41]
  wire  r_count_94_reset; // @[SWChisel.scala 171:41]
  wire  r_count_94_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_94_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_95_clock; // @[SWChisel.scala 171:41]
  wire  r_count_95_reset; // @[SWChisel.scala 171:41]
  wire  r_count_95_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_95_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_96_clock; // @[SWChisel.scala 171:41]
  wire  r_count_96_reset; // @[SWChisel.scala 171:41]
  wire  r_count_96_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_96_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_97_clock; // @[SWChisel.scala 171:41]
  wire  r_count_97_reset; // @[SWChisel.scala 171:41]
  wire  r_count_97_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_97_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_98_clock; // @[SWChisel.scala 171:41]
  wire  r_count_98_reset; // @[SWChisel.scala 171:41]
  wire  r_count_98_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_98_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_99_clock; // @[SWChisel.scala 171:41]
  wire  r_count_99_reset; // @[SWChisel.scala 171:41]
  wire  r_count_99_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_99_io_out; // @[SWChisel.scala 171:41]
  wire  max_clock; // @[SWChisel.scala 174:19]
  wire  max_reset; // @[SWChisel.scala 174:19]
  wire  max_io_start; // @[SWChisel.scala 174:19]
  wire [15:0] max_io_in; // @[SWChisel.scala 174:19]
  wire  max_io_done; // @[SWChisel.scala 174:19]
  wire [15:0] max_io_out; // @[SWChisel.scala 174:19]
  reg [15:0] E_0; // @[SWChisel.scala 162:18]
  reg [15:0] E_1; // @[SWChisel.scala 162:18]
  reg [15:0] E_2; // @[SWChisel.scala 162:18]
  reg [15:0] E_3; // @[SWChisel.scala 162:18]
  reg [15:0] E_4; // @[SWChisel.scala 162:18]
  reg [15:0] E_5; // @[SWChisel.scala 162:18]
  reg [15:0] E_6; // @[SWChisel.scala 162:18]
  reg [15:0] E_7; // @[SWChisel.scala 162:18]
  reg [15:0] E_8; // @[SWChisel.scala 162:18]
  reg [15:0] E_9; // @[SWChisel.scala 162:18]
  reg [15:0] E_10; // @[SWChisel.scala 162:18]
  reg [15:0] E_11; // @[SWChisel.scala 162:18]
  reg [15:0] E_12; // @[SWChisel.scala 162:18]
  reg [15:0] E_13; // @[SWChisel.scala 162:18]
  reg [15:0] E_14; // @[SWChisel.scala 162:18]
  reg [15:0] E_15; // @[SWChisel.scala 162:18]
  reg [15:0] E_16; // @[SWChisel.scala 162:18]
  reg [15:0] E_17; // @[SWChisel.scala 162:18]
  reg [15:0] E_18; // @[SWChisel.scala 162:18]
  reg [15:0] E_19; // @[SWChisel.scala 162:18]
  reg [15:0] E_20; // @[SWChisel.scala 162:18]
  reg [15:0] E_21; // @[SWChisel.scala 162:18]
  reg [15:0] E_22; // @[SWChisel.scala 162:18]
  reg [15:0] E_23; // @[SWChisel.scala 162:18]
  reg [15:0] E_24; // @[SWChisel.scala 162:18]
  reg [15:0] E_25; // @[SWChisel.scala 162:18]
  reg [15:0] E_26; // @[SWChisel.scala 162:18]
  reg [15:0] E_27; // @[SWChisel.scala 162:18]
  reg [15:0] E_28; // @[SWChisel.scala 162:18]
  reg [15:0] E_29; // @[SWChisel.scala 162:18]
  reg [15:0] E_30; // @[SWChisel.scala 162:18]
  reg [15:0] E_31; // @[SWChisel.scala 162:18]
  reg [15:0] E_32; // @[SWChisel.scala 162:18]
  reg [15:0] E_33; // @[SWChisel.scala 162:18]
  reg [15:0] E_34; // @[SWChisel.scala 162:18]
  reg [15:0] E_35; // @[SWChisel.scala 162:18]
  reg [15:0] E_36; // @[SWChisel.scala 162:18]
  reg [15:0] E_37; // @[SWChisel.scala 162:18]
  reg [15:0] E_38; // @[SWChisel.scala 162:18]
  reg [15:0] E_39; // @[SWChisel.scala 162:18]
  reg [15:0] E_40; // @[SWChisel.scala 162:18]
  reg [15:0] E_41; // @[SWChisel.scala 162:18]
  reg [15:0] E_42; // @[SWChisel.scala 162:18]
  reg [15:0] E_43; // @[SWChisel.scala 162:18]
  reg [15:0] E_44; // @[SWChisel.scala 162:18]
  reg [15:0] E_45; // @[SWChisel.scala 162:18]
  reg [15:0] E_46; // @[SWChisel.scala 162:18]
  reg [15:0] E_47; // @[SWChisel.scala 162:18]
  reg [15:0] E_48; // @[SWChisel.scala 162:18]
  reg [15:0] E_49; // @[SWChisel.scala 162:18]
  reg [15:0] E_50; // @[SWChisel.scala 162:18]
  reg [15:0] E_51; // @[SWChisel.scala 162:18]
  reg [15:0] E_52; // @[SWChisel.scala 162:18]
  reg [15:0] E_53; // @[SWChisel.scala 162:18]
  reg [15:0] E_54; // @[SWChisel.scala 162:18]
  reg [15:0] E_55; // @[SWChisel.scala 162:18]
  reg [15:0] E_56; // @[SWChisel.scala 162:18]
  reg [15:0] E_57; // @[SWChisel.scala 162:18]
  reg [15:0] E_58; // @[SWChisel.scala 162:18]
  reg [15:0] E_59; // @[SWChisel.scala 162:18]
  reg [15:0] E_60; // @[SWChisel.scala 162:18]
  reg [15:0] E_61; // @[SWChisel.scala 162:18]
  reg [15:0] E_62; // @[SWChisel.scala 162:18]
  reg [15:0] E_63; // @[SWChisel.scala 162:18]
  reg [15:0] E_64; // @[SWChisel.scala 162:18]
  reg [15:0] E_65; // @[SWChisel.scala 162:18]
  reg [15:0] E_66; // @[SWChisel.scala 162:18]
  reg [15:0] E_67; // @[SWChisel.scala 162:18]
  reg [15:0] E_68; // @[SWChisel.scala 162:18]
  reg [15:0] E_69; // @[SWChisel.scala 162:18]
  reg [15:0] E_70; // @[SWChisel.scala 162:18]
  reg [15:0] E_71; // @[SWChisel.scala 162:18]
  reg [15:0] E_72; // @[SWChisel.scala 162:18]
  reg [15:0] E_73; // @[SWChisel.scala 162:18]
  reg [15:0] E_74; // @[SWChisel.scala 162:18]
  reg [15:0] E_75; // @[SWChisel.scala 162:18]
  reg [15:0] E_76; // @[SWChisel.scala 162:18]
  reg [15:0] E_77; // @[SWChisel.scala 162:18]
  reg [15:0] E_78; // @[SWChisel.scala 162:18]
  reg [15:0] E_79; // @[SWChisel.scala 162:18]
  reg [15:0] E_80; // @[SWChisel.scala 162:18]
  reg [15:0] E_81; // @[SWChisel.scala 162:18]
  reg [15:0] E_82; // @[SWChisel.scala 162:18]
  reg [15:0] E_83; // @[SWChisel.scala 162:18]
  reg [15:0] E_84; // @[SWChisel.scala 162:18]
  reg [15:0] E_85; // @[SWChisel.scala 162:18]
  reg [15:0] E_86; // @[SWChisel.scala 162:18]
  reg [15:0] E_87; // @[SWChisel.scala 162:18]
  reg [15:0] E_88; // @[SWChisel.scala 162:18]
  reg [15:0] E_89; // @[SWChisel.scala 162:18]
  reg [15:0] E_90; // @[SWChisel.scala 162:18]
  reg [15:0] E_91; // @[SWChisel.scala 162:18]
  reg [15:0] E_92; // @[SWChisel.scala 162:18]
  reg [15:0] E_93; // @[SWChisel.scala 162:18]
  reg [15:0] E_94; // @[SWChisel.scala 162:18]
  reg [15:0] E_95; // @[SWChisel.scala 162:18]
  reg [15:0] E_96; // @[SWChisel.scala 162:18]
  reg [15:0] E_97; // @[SWChisel.scala 162:18]
  reg [15:0] E_98; // @[SWChisel.scala 162:18]
  reg [15:0] E_99; // @[SWChisel.scala 162:18]
  reg [15:0] F_1; // @[SWChisel.scala 163:18]
  reg [15:0] F_2; // @[SWChisel.scala 163:18]
  reg [15:0] F_3; // @[SWChisel.scala 163:18]
  reg [15:0] F_4; // @[SWChisel.scala 163:18]
  reg [15:0] F_5; // @[SWChisel.scala 163:18]
  reg [15:0] F_6; // @[SWChisel.scala 163:18]
  reg [15:0] F_7; // @[SWChisel.scala 163:18]
  reg [15:0] F_8; // @[SWChisel.scala 163:18]
  reg [15:0] F_9; // @[SWChisel.scala 163:18]
  reg [15:0] F_10; // @[SWChisel.scala 163:18]
  reg [15:0] F_11; // @[SWChisel.scala 163:18]
  reg [15:0] F_12; // @[SWChisel.scala 163:18]
  reg [15:0] F_13; // @[SWChisel.scala 163:18]
  reg [15:0] F_14; // @[SWChisel.scala 163:18]
  reg [15:0] F_15; // @[SWChisel.scala 163:18]
  reg [15:0] F_16; // @[SWChisel.scala 163:18]
  reg [15:0] F_17; // @[SWChisel.scala 163:18]
  reg [15:0] F_18; // @[SWChisel.scala 163:18]
  reg [15:0] F_19; // @[SWChisel.scala 163:18]
  reg [15:0] F_20; // @[SWChisel.scala 163:18]
  reg [15:0] F_21; // @[SWChisel.scala 163:18]
  reg [15:0] F_22; // @[SWChisel.scala 163:18]
  reg [15:0] F_23; // @[SWChisel.scala 163:18]
  reg [15:0] F_24; // @[SWChisel.scala 163:18]
  reg [15:0] F_25; // @[SWChisel.scala 163:18]
  reg [15:0] F_26; // @[SWChisel.scala 163:18]
  reg [15:0] F_27; // @[SWChisel.scala 163:18]
  reg [15:0] F_28; // @[SWChisel.scala 163:18]
  reg [15:0] F_29; // @[SWChisel.scala 163:18]
  reg [15:0] F_30; // @[SWChisel.scala 163:18]
  reg [15:0] F_31; // @[SWChisel.scala 163:18]
  reg [15:0] F_32; // @[SWChisel.scala 163:18]
  reg [15:0] F_33; // @[SWChisel.scala 163:18]
  reg [15:0] F_34; // @[SWChisel.scala 163:18]
  reg [15:0] F_35; // @[SWChisel.scala 163:18]
  reg [15:0] F_36; // @[SWChisel.scala 163:18]
  reg [15:0] F_37; // @[SWChisel.scala 163:18]
  reg [15:0] F_38; // @[SWChisel.scala 163:18]
  reg [15:0] F_39; // @[SWChisel.scala 163:18]
  reg [15:0] F_40; // @[SWChisel.scala 163:18]
  reg [15:0] F_41; // @[SWChisel.scala 163:18]
  reg [15:0] F_42; // @[SWChisel.scala 163:18]
  reg [15:0] F_43; // @[SWChisel.scala 163:18]
  reg [15:0] F_44; // @[SWChisel.scala 163:18]
  reg [15:0] F_45; // @[SWChisel.scala 163:18]
  reg [15:0] F_46; // @[SWChisel.scala 163:18]
  reg [15:0] F_47; // @[SWChisel.scala 163:18]
  reg [15:0] F_48; // @[SWChisel.scala 163:18]
  reg [15:0] F_49; // @[SWChisel.scala 163:18]
  reg [15:0] F_50; // @[SWChisel.scala 163:18]
  reg [15:0] F_51; // @[SWChisel.scala 163:18]
  reg [15:0] F_52; // @[SWChisel.scala 163:18]
  reg [15:0] F_53; // @[SWChisel.scala 163:18]
  reg [15:0] F_54; // @[SWChisel.scala 163:18]
  reg [15:0] F_55; // @[SWChisel.scala 163:18]
  reg [15:0] F_56; // @[SWChisel.scala 163:18]
  reg [15:0] F_57; // @[SWChisel.scala 163:18]
  reg [15:0] F_58; // @[SWChisel.scala 163:18]
  reg [15:0] F_59; // @[SWChisel.scala 163:18]
  reg [15:0] F_60; // @[SWChisel.scala 163:18]
  reg [15:0] F_61; // @[SWChisel.scala 163:18]
  reg [15:0] F_62; // @[SWChisel.scala 163:18]
  reg [15:0] F_63; // @[SWChisel.scala 163:18]
  reg [15:0] F_64; // @[SWChisel.scala 163:18]
  reg [15:0] F_65; // @[SWChisel.scala 163:18]
  reg [15:0] F_66; // @[SWChisel.scala 163:18]
  reg [15:0] F_67; // @[SWChisel.scala 163:18]
  reg [15:0] F_68; // @[SWChisel.scala 163:18]
  reg [15:0] F_69; // @[SWChisel.scala 163:18]
  reg [15:0] F_70; // @[SWChisel.scala 163:18]
  reg [15:0] F_71; // @[SWChisel.scala 163:18]
  reg [15:0] F_72; // @[SWChisel.scala 163:18]
  reg [15:0] F_73; // @[SWChisel.scala 163:18]
  reg [15:0] F_74; // @[SWChisel.scala 163:18]
  reg [15:0] F_75; // @[SWChisel.scala 163:18]
  reg [15:0] F_76; // @[SWChisel.scala 163:18]
  reg [15:0] F_77; // @[SWChisel.scala 163:18]
  reg [15:0] F_78; // @[SWChisel.scala 163:18]
  reg [15:0] F_79; // @[SWChisel.scala 163:18]
  reg [15:0] F_80; // @[SWChisel.scala 163:18]
  reg [15:0] F_81; // @[SWChisel.scala 163:18]
  reg [15:0] F_82; // @[SWChisel.scala 163:18]
  reg [15:0] F_83; // @[SWChisel.scala 163:18]
  reg [15:0] F_84; // @[SWChisel.scala 163:18]
  reg [15:0] F_85; // @[SWChisel.scala 163:18]
  reg [15:0] F_86; // @[SWChisel.scala 163:18]
  reg [15:0] F_87; // @[SWChisel.scala 163:18]
  reg [15:0] F_88; // @[SWChisel.scala 163:18]
  reg [15:0] F_89; // @[SWChisel.scala 163:18]
  reg [15:0] F_90; // @[SWChisel.scala 163:18]
  reg [15:0] F_91; // @[SWChisel.scala 163:18]
  reg [15:0] F_92; // @[SWChisel.scala 163:18]
  reg [15:0] F_93; // @[SWChisel.scala 163:18]
  reg [15:0] F_94; // @[SWChisel.scala 163:18]
  reg [15:0] F_95; // @[SWChisel.scala 163:18]
  reg [15:0] F_96; // @[SWChisel.scala 163:18]
  reg [15:0] F_97; // @[SWChisel.scala 163:18]
  reg [15:0] F_98; // @[SWChisel.scala 163:18]
  reg [15:0] F_99; // @[SWChisel.scala 163:18]
  reg [15:0] V1_0; // @[SWChisel.scala 164:19]
  reg [15:0] V1_1; // @[SWChisel.scala 164:19]
  reg [15:0] V1_2; // @[SWChisel.scala 164:19]
  reg [15:0] V1_3; // @[SWChisel.scala 164:19]
  reg [15:0] V1_4; // @[SWChisel.scala 164:19]
  reg [15:0] V1_5; // @[SWChisel.scala 164:19]
  reg [15:0] V1_6; // @[SWChisel.scala 164:19]
  reg [15:0] V1_7; // @[SWChisel.scala 164:19]
  reg [15:0] V1_8; // @[SWChisel.scala 164:19]
  reg [15:0] V1_9; // @[SWChisel.scala 164:19]
  reg [15:0] V1_10; // @[SWChisel.scala 164:19]
  reg [15:0] V1_11; // @[SWChisel.scala 164:19]
  reg [15:0] V1_12; // @[SWChisel.scala 164:19]
  reg [15:0] V1_13; // @[SWChisel.scala 164:19]
  reg [15:0] V1_14; // @[SWChisel.scala 164:19]
  reg [15:0] V1_15; // @[SWChisel.scala 164:19]
  reg [15:0] V1_16; // @[SWChisel.scala 164:19]
  reg [15:0] V1_17; // @[SWChisel.scala 164:19]
  reg [15:0] V1_18; // @[SWChisel.scala 164:19]
  reg [15:0] V1_19; // @[SWChisel.scala 164:19]
  reg [15:0] V1_20; // @[SWChisel.scala 164:19]
  reg [15:0] V1_21; // @[SWChisel.scala 164:19]
  reg [15:0] V1_22; // @[SWChisel.scala 164:19]
  reg [15:0] V1_23; // @[SWChisel.scala 164:19]
  reg [15:0] V1_24; // @[SWChisel.scala 164:19]
  reg [15:0] V1_25; // @[SWChisel.scala 164:19]
  reg [15:0] V1_26; // @[SWChisel.scala 164:19]
  reg [15:0] V1_27; // @[SWChisel.scala 164:19]
  reg [15:0] V1_28; // @[SWChisel.scala 164:19]
  reg [15:0] V1_29; // @[SWChisel.scala 164:19]
  reg [15:0] V1_30; // @[SWChisel.scala 164:19]
  reg [15:0] V1_31; // @[SWChisel.scala 164:19]
  reg [15:0] V1_32; // @[SWChisel.scala 164:19]
  reg [15:0] V1_33; // @[SWChisel.scala 164:19]
  reg [15:0] V1_34; // @[SWChisel.scala 164:19]
  reg [15:0] V1_35; // @[SWChisel.scala 164:19]
  reg [15:0] V1_36; // @[SWChisel.scala 164:19]
  reg [15:0] V1_37; // @[SWChisel.scala 164:19]
  reg [15:0] V1_38; // @[SWChisel.scala 164:19]
  reg [15:0] V1_39; // @[SWChisel.scala 164:19]
  reg [15:0] V1_40; // @[SWChisel.scala 164:19]
  reg [15:0] V1_41; // @[SWChisel.scala 164:19]
  reg [15:0] V1_42; // @[SWChisel.scala 164:19]
  reg [15:0] V1_43; // @[SWChisel.scala 164:19]
  reg [15:0] V1_44; // @[SWChisel.scala 164:19]
  reg [15:0] V1_45; // @[SWChisel.scala 164:19]
  reg [15:0] V1_46; // @[SWChisel.scala 164:19]
  reg [15:0] V1_47; // @[SWChisel.scala 164:19]
  reg [15:0] V1_48; // @[SWChisel.scala 164:19]
  reg [15:0] V1_49; // @[SWChisel.scala 164:19]
  reg [15:0] V1_50; // @[SWChisel.scala 164:19]
  reg [15:0] V1_51; // @[SWChisel.scala 164:19]
  reg [15:0] V1_52; // @[SWChisel.scala 164:19]
  reg [15:0] V1_53; // @[SWChisel.scala 164:19]
  reg [15:0] V1_54; // @[SWChisel.scala 164:19]
  reg [15:0] V1_55; // @[SWChisel.scala 164:19]
  reg [15:0] V1_56; // @[SWChisel.scala 164:19]
  reg [15:0] V1_57; // @[SWChisel.scala 164:19]
  reg [15:0] V1_58; // @[SWChisel.scala 164:19]
  reg [15:0] V1_59; // @[SWChisel.scala 164:19]
  reg [15:0] V1_60; // @[SWChisel.scala 164:19]
  reg [15:0] V1_61; // @[SWChisel.scala 164:19]
  reg [15:0] V1_62; // @[SWChisel.scala 164:19]
  reg [15:0] V1_63; // @[SWChisel.scala 164:19]
  reg [15:0] V1_64; // @[SWChisel.scala 164:19]
  reg [15:0] V1_65; // @[SWChisel.scala 164:19]
  reg [15:0] V1_66; // @[SWChisel.scala 164:19]
  reg [15:0] V1_67; // @[SWChisel.scala 164:19]
  reg [15:0] V1_68; // @[SWChisel.scala 164:19]
  reg [15:0] V1_69; // @[SWChisel.scala 164:19]
  reg [15:0] V1_70; // @[SWChisel.scala 164:19]
  reg [15:0] V1_71; // @[SWChisel.scala 164:19]
  reg [15:0] V1_72; // @[SWChisel.scala 164:19]
  reg [15:0] V1_73; // @[SWChisel.scala 164:19]
  reg [15:0] V1_74; // @[SWChisel.scala 164:19]
  reg [15:0] V1_75; // @[SWChisel.scala 164:19]
  reg [15:0] V1_76; // @[SWChisel.scala 164:19]
  reg [15:0] V1_77; // @[SWChisel.scala 164:19]
  reg [15:0] V1_78; // @[SWChisel.scala 164:19]
  reg [15:0] V1_79; // @[SWChisel.scala 164:19]
  reg [15:0] V1_80; // @[SWChisel.scala 164:19]
  reg [15:0] V1_81; // @[SWChisel.scala 164:19]
  reg [15:0] V1_82; // @[SWChisel.scala 164:19]
  reg [15:0] V1_83; // @[SWChisel.scala 164:19]
  reg [15:0] V1_84; // @[SWChisel.scala 164:19]
  reg [15:0] V1_85; // @[SWChisel.scala 164:19]
  reg [15:0] V1_86; // @[SWChisel.scala 164:19]
  reg [15:0] V1_87; // @[SWChisel.scala 164:19]
  reg [15:0] V1_88; // @[SWChisel.scala 164:19]
  reg [15:0] V1_89; // @[SWChisel.scala 164:19]
  reg [15:0] V1_90; // @[SWChisel.scala 164:19]
  reg [15:0] V1_91; // @[SWChisel.scala 164:19]
  reg [15:0] V1_92; // @[SWChisel.scala 164:19]
  reg [15:0] V1_93; // @[SWChisel.scala 164:19]
  reg [15:0] V1_94; // @[SWChisel.scala 164:19]
  reg [15:0] V1_95; // @[SWChisel.scala 164:19]
  reg [15:0] V1_96; // @[SWChisel.scala 164:19]
  reg [15:0] V1_97; // @[SWChisel.scala 164:19]
  reg [15:0] V1_98; // @[SWChisel.scala 164:19]
  reg [15:0] V1_99; // @[SWChisel.scala 164:19]
  reg [15:0] V1_100; // @[SWChisel.scala 164:19]
  reg [15:0] V2_0; // @[SWChisel.scala 166:19]
  reg [15:0] V2_1; // @[SWChisel.scala 166:19]
  reg [15:0] V2_2; // @[SWChisel.scala 166:19]
  reg [15:0] V2_3; // @[SWChisel.scala 166:19]
  reg [15:0] V2_4; // @[SWChisel.scala 166:19]
  reg [15:0] V2_5; // @[SWChisel.scala 166:19]
  reg [15:0] V2_6; // @[SWChisel.scala 166:19]
  reg [15:0] V2_7; // @[SWChisel.scala 166:19]
  reg [15:0] V2_8; // @[SWChisel.scala 166:19]
  reg [15:0] V2_9; // @[SWChisel.scala 166:19]
  reg [15:0] V2_10; // @[SWChisel.scala 166:19]
  reg [15:0] V2_11; // @[SWChisel.scala 166:19]
  reg [15:0] V2_12; // @[SWChisel.scala 166:19]
  reg [15:0] V2_13; // @[SWChisel.scala 166:19]
  reg [15:0] V2_14; // @[SWChisel.scala 166:19]
  reg [15:0] V2_15; // @[SWChisel.scala 166:19]
  reg [15:0] V2_16; // @[SWChisel.scala 166:19]
  reg [15:0] V2_17; // @[SWChisel.scala 166:19]
  reg [15:0] V2_18; // @[SWChisel.scala 166:19]
  reg [15:0] V2_19; // @[SWChisel.scala 166:19]
  reg [15:0] V2_20; // @[SWChisel.scala 166:19]
  reg [15:0] V2_21; // @[SWChisel.scala 166:19]
  reg [15:0] V2_22; // @[SWChisel.scala 166:19]
  reg [15:0] V2_23; // @[SWChisel.scala 166:19]
  reg [15:0] V2_24; // @[SWChisel.scala 166:19]
  reg [15:0] V2_25; // @[SWChisel.scala 166:19]
  reg [15:0] V2_26; // @[SWChisel.scala 166:19]
  reg [15:0] V2_27; // @[SWChisel.scala 166:19]
  reg [15:0] V2_28; // @[SWChisel.scala 166:19]
  reg [15:0] V2_29; // @[SWChisel.scala 166:19]
  reg [15:0] V2_30; // @[SWChisel.scala 166:19]
  reg [15:0] V2_31; // @[SWChisel.scala 166:19]
  reg [15:0] V2_32; // @[SWChisel.scala 166:19]
  reg [15:0] V2_33; // @[SWChisel.scala 166:19]
  reg [15:0] V2_34; // @[SWChisel.scala 166:19]
  reg [15:0] V2_35; // @[SWChisel.scala 166:19]
  reg [15:0] V2_36; // @[SWChisel.scala 166:19]
  reg [15:0] V2_37; // @[SWChisel.scala 166:19]
  reg [15:0] V2_38; // @[SWChisel.scala 166:19]
  reg [15:0] V2_39; // @[SWChisel.scala 166:19]
  reg [15:0] V2_40; // @[SWChisel.scala 166:19]
  reg [15:0] V2_41; // @[SWChisel.scala 166:19]
  reg [15:0] V2_42; // @[SWChisel.scala 166:19]
  reg [15:0] V2_43; // @[SWChisel.scala 166:19]
  reg [15:0] V2_44; // @[SWChisel.scala 166:19]
  reg [15:0] V2_45; // @[SWChisel.scala 166:19]
  reg [15:0] V2_46; // @[SWChisel.scala 166:19]
  reg [15:0] V2_47; // @[SWChisel.scala 166:19]
  reg [15:0] V2_48; // @[SWChisel.scala 166:19]
  reg [15:0] V2_49; // @[SWChisel.scala 166:19]
  reg [15:0] V2_50; // @[SWChisel.scala 166:19]
  reg [15:0] V2_51; // @[SWChisel.scala 166:19]
  reg [15:0] V2_52; // @[SWChisel.scala 166:19]
  reg [15:0] V2_53; // @[SWChisel.scala 166:19]
  reg [15:0] V2_54; // @[SWChisel.scala 166:19]
  reg [15:0] V2_55; // @[SWChisel.scala 166:19]
  reg [15:0] V2_56; // @[SWChisel.scala 166:19]
  reg [15:0] V2_57; // @[SWChisel.scala 166:19]
  reg [15:0] V2_58; // @[SWChisel.scala 166:19]
  reg [15:0] V2_59; // @[SWChisel.scala 166:19]
  reg [15:0] V2_60; // @[SWChisel.scala 166:19]
  reg [15:0] V2_61; // @[SWChisel.scala 166:19]
  reg [15:0] V2_62; // @[SWChisel.scala 166:19]
  reg [15:0] V2_63; // @[SWChisel.scala 166:19]
  reg [15:0] V2_64; // @[SWChisel.scala 166:19]
  reg [15:0] V2_65; // @[SWChisel.scala 166:19]
  reg [15:0] V2_66; // @[SWChisel.scala 166:19]
  reg [15:0] V2_67; // @[SWChisel.scala 166:19]
  reg [15:0] V2_68; // @[SWChisel.scala 166:19]
  reg [15:0] V2_69; // @[SWChisel.scala 166:19]
  reg [15:0] V2_70; // @[SWChisel.scala 166:19]
  reg [15:0] V2_71; // @[SWChisel.scala 166:19]
  reg [15:0] V2_72; // @[SWChisel.scala 166:19]
  reg [15:0] V2_73; // @[SWChisel.scala 166:19]
  reg [15:0] V2_74; // @[SWChisel.scala 166:19]
  reg [15:0] V2_75; // @[SWChisel.scala 166:19]
  reg [15:0] V2_76; // @[SWChisel.scala 166:19]
  reg [15:0] V2_77; // @[SWChisel.scala 166:19]
  reg [15:0] V2_78; // @[SWChisel.scala 166:19]
  reg [15:0] V2_79; // @[SWChisel.scala 166:19]
  reg [15:0] V2_80; // @[SWChisel.scala 166:19]
  reg [15:0] V2_81; // @[SWChisel.scala 166:19]
  reg [15:0] V2_82; // @[SWChisel.scala 166:19]
  reg [15:0] V2_83; // @[SWChisel.scala 166:19]
  reg [15:0] V2_84; // @[SWChisel.scala 166:19]
  reg [15:0] V2_85; // @[SWChisel.scala 166:19]
  reg [15:0] V2_86; // @[SWChisel.scala 166:19]
  reg [15:0] V2_87; // @[SWChisel.scala 166:19]
  reg [15:0] V2_88; // @[SWChisel.scala 166:19]
  reg [15:0] V2_89; // @[SWChisel.scala 166:19]
  reg [15:0] V2_90; // @[SWChisel.scala 166:19]
  reg [15:0] V2_91; // @[SWChisel.scala 166:19]
  reg [15:0] V2_92; // @[SWChisel.scala 166:19]
  reg [15:0] V2_93; // @[SWChisel.scala 166:19]
  reg [15:0] V2_94; // @[SWChisel.scala 166:19]
  reg [15:0] V2_95; // @[SWChisel.scala 166:19]
  reg [15:0] V2_96; // @[SWChisel.scala 166:19]
  reg [15:0] V2_97; // @[SWChisel.scala 166:19]
  reg [15:0] V2_98; // @[SWChisel.scala 166:19]
  reg [15:0] V2_99; // @[SWChisel.scala 166:19]
  reg  start_reg_0; // @[SWChisel.scala 167:26]
  reg  start_reg_1; // @[SWChisel.scala 167:26]
  reg  start_reg_2; // @[SWChisel.scala 167:26]
  reg  start_reg_3; // @[SWChisel.scala 167:26]
  reg  start_reg_4; // @[SWChisel.scala 167:26]
  reg  start_reg_5; // @[SWChisel.scala 167:26]
  reg  start_reg_6; // @[SWChisel.scala 167:26]
  reg  start_reg_7; // @[SWChisel.scala 167:26]
  reg  start_reg_8; // @[SWChisel.scala 167:26]
  reg  start_reg_9; // @[SWChisel.scala 167:26]
  reg  start_reg_10; // @[SWChisel.scala 167:26]
  reg  start_reg_11; // @[SWChisel.scala 167:26]
  reg  start_reg_12; // @[SWChisel.scala 167:26]
  reg  start_reg_13; // @[SWChisel.scala 167:26]
  reg  start_reg_14; // @[SWChisel.scala 167:26]
  reg  start_reg_15; // @[SWChisel.scala 167:26]
  reg  start_reg_16; // @[SWChisel.scala 167:26]
  reg  start_reg_17; // @[SWChisel.scala 167:26]
  reg  start_reg_18; // @[SWChisel.scala 167:26]
  reg  start_reg_19; // @[SWChisel.scala 167:26]
  reg  start_reg_20; // @[SWChisel.scala 167:26]
  reg  start_reg_21; // @[SWChisel.scala 167:26]
  reg  start_reg_22; // @[SWChisel.scala 167:26]
  reg  start_reg_23; // @[SWChisel.scala 167:26]
  reg  start_reg_24; // @[SWChisel.scala 167:26]
  reg  start_reg_25; // @[SWChisel.scala 167:26]
  reg  start_reg_26; // @[SWChisel.scala 167:26]
  reg  start_reg_27; // @[SWChisel.scala 167:26]
  reg  start_reg_28; // @[SWChisel.scala 167:26]
  reg  start_reg_29; // @[SWChisel.scala 167:26]
  reg  start_reg_30; // @[SWChisel.scala 167:26]
  reg  start_reg_31; // @[SWChisel.scala 167:26]
  reg  start_reg_32; // @[SWChisel.scala 167:26]
  reg  start_reg_33; // @[SWChisel.scala 167:26]
  reg  start_reg_34; // @[SWChisel.scala 167:26]
  reg  start_reg_35; // @[SWChisel.scala 167:26]
  reg  start_reg_36; // @[SWChisel.scala 167:26]
  reg  start_reg_37; // @[SWChisel.scala 167:26]
  reg  start_reg_38; // @[SWChisel.scala 167:26]
  reg  start_reg_39; // @[SWChisel.scala 167:26]
  reg  start_reg_40; // @[SWChisel.scala 167:26]
  reg  start_reg_41; // @[SWChisel.scala 167:26]
  reg  start_reg_42; // @[SWChisel.scala 167:26]
  reg  start_reg_43; // @[SWChisel.scala 167:26]
  reg  start_reg_44; // @[SWChisel.scala 167:26]
  reg  start_reg_45; // @[SWChisel.scala 167:26]
  reg  start_reg_46; // @[SWChisel.scala 167:26]
  reg  start_reg_47; // @[SWChisel.scala 167:26]
  reg  start_reg_48; // @[SWChisel.scala 167:26]
  reg  start_reg_49; // @[SWChisel.scala 167:26]
  reg  start_reg_50; // @[SWChisel.scala 167:26]
  reg  start_reg_51; // @[SWChisel.scala 167:26]
  reg  start_reg_52; // @[SWChisel.scala 167:26]
  reg  start_reg_53; // @[SWChisel.scala 167:26]
  reg  start_reg_54; // @[SWChisel.scala 167:26]
  reg  start_reg_55; // @[SWChisel.scala 167:26]
  reg  start_reg_56; // @[SWChisel.scala 167:26]
  reg  start_reg_57; // @[SWChisel.scala 167:26]
  reg  start_reg_58; // @[SWChisel.scala 167:26]
  reg  start_reg_59; // @[SWChisel.scala 167:26]
  reg  start_reg_60; // @[SWChisel.scala 167:26]
  reg  start_reg_61; // @[SWChisel.scala 167:26]
  reg  start_reg_62; // @[SWChisel.scala 167:26]
  reg  start_reg_63; // @[SWChisel.scala 167:26]
  reg  start_reg_64; // @[SWChisel.scala 167:26]
  reg  start_reg_65; // @[SWChisel.scala 167:26]
  reg  start_reg_66; // @[SWChisel.scala 167:26]
  reg  start_reg_67; // @[SWChisel.scala 167:26]
  reg  start_reg_68; // @[SWChisel.scala 167:26]
  reg  start_reg_69; // @[SWChisel.scala 167:26]
  reg  start_reg_70; // @[SWChisel.scala 167:26]
  reg  start_reg_71; // @[SWChisel.scala 167:26]
  reg  start_reg_72; // @[SWChisel.scala 167:26]
  reg  start_reg_73; // @[SWChisel.scala 167:26]
  reg  start_reg_74; // @[SWChisel.scala 167:26]
  reg  start_reg_75; // @[SWChisel.scala 167:26]
  reg  start_reg_76; // @[SWChisel.scala 167:26]
  reg  start_reg_77; // @[SWChisel.scala 167:26]
  reg  start_reg_78; // @[SWChisel.scala 167:26]
  reg  start_reg_79; // @[SWChisel.scala 167:26]
  reg  start_reg_80; // @[SWChisel.scala 167:26]
  reg  start_reg_81; // @[SWChisel.scala 167:26]
  reg  start_reg_82; // @[SWChisel.scala 167:26]
  reg  start_reg_83; // @[SWChisel.scala 167:26]
  reg  start_reg_84; // @[SWChisel.scala 167:26]
  reg  start_reg_85; // @[SWChisel.scala 167:26]
  reg  start_reg_86; // @[SWChisel.scala 167:26]
  reg  start_reg_87; // @[SWChisel.scala 167:26]
  reg  start_reg_88; // @[SWChisel.scala 167:26]
  reg  start_reg_89; // @[SWChisel.scala 167:26]
  reg  start_reg_90; // @[SWChisel.scala 167:26]
  reg  start_reg_91; // @[SWChisel.scala 167:26]
  reg  start_reg_92; // @[SWChisel.scala 167:26]
  reg  start_reg_93; // @[SWChisel.scala 167:26]
  reg  start_reg_94; // @[SWChisel.scala 167:26]
  reg  start_reg_95; // @[SWChisel.scala 167:26]
  reg  start_reg_96; // @[SWChisel.scala 167:26]
  reg  start_reg_97; // @[SWChisel.scala 167:26]
  reg  start_reg_98; // @[SWChisel.scala 167:26]
  reg  start_reg_99; // @[SWChisel.scala 167:26]
  wire [1:0] _GEN_301 = 8'h1 == r_count_0_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_302 = 8'h2 == r_count_0_io_out ? io_r_2_b : _GEN_301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_303 = 8'h3 == r_count_0_io_out ? io_r_3_b : _GEN_302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_304 = 8'h4 == r_count_0_io_out ? io_r_4_b : _GEN_303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_305 = 8'h5 == r_count_0_io_out ? io_r_5_b : _GEN_304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_306 = 8'h6 == r_count_0_io_out ? io_r_6_b : _GEN_305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_307 = 8'h7 == r_count_0_io_out ? io_r_7_b : _GEN_306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_308 = 8'h8 == r_count_0_io_out ? io_r_8_b : _GEN_307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_309 = 8'h9 == r_count_0_io_out ? io_r_9_b : _GEN_308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_310 = 8'ha == r_count_0_io_out ? io_r_10_b : _GEN_309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_311 = 8'hb == r_count_0_io_out ? io_r_11_b : _GEN_310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_312 = 8'hc == r_count_0_io_out ? io_r_12_b : _GEN_311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_313 = 8'hd == r_count_0_io_out ? io_r_13_b : _GEN_312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_314 = 8'he == r_count_0_io_out ? io_r_14_b : _GEN_313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_315 = 8'hf == r_count_0_io_out ? io_r_15_b : _GEN_314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_316 = 8'h10 == r_count_0_io_out ? io_r_16_b : _GEN_315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_317 = 8'h11 == r_count_0_io_out ? io_r_17_b : _GEN_316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_318 = 8'h12 == r_count_0_io_out ? io_r_18_b : _GEN_317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_319 = 8'h13 == r_count_0_io_out ? io_r_19_b : _GEN_318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_320 = 8'h14 == r_count_0_io_out ? io_r_20_b : _GEN_319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_321 = 8'h15 == r_count_0_io_out ? io_r_21_b : _GEN_320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_322 = 8'h16 == r_count_0_io_out ? io_r_22_b : _GEN_321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_323 = 8'h17 == r_count_0_io_out ? io_r_23_b : _GEN_322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_324 = 8'h18 == r_count_0_io_out ? io_r_24_b : _GEN_323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_325 = 8'h19 == r_count_0_io_out ? io_r_25_b : _GEN_324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_326 = 8'h1a == r_count_0_io_out ? io_r_26_b : _GEN_325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_327 = 8'h1b == r_count_0_io_out ? io_r_27_b : _GEN_326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_328 = 8'h1c == r_count_0_io_out ? io_r_28_b : _GEN_327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_329 = 8'h1d == r_count_0_io_out ? io_r_29_b : _GEN_328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_330 = 8'h1e == r_count_0_io_out ? io_r_30_b : _GEN_329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_331 = 8'h1f == r_count_0_io_out ? io_r_31_b : _GEN_330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_332 = 8'h20 == r_count_0_io_out ? io_r_32_b : _GEN_331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_333 = 8'h21 == r_count_0_io_out ? io_r_33_b : _GEN_332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_334 = 8'h22 == r_count_0_io_out ? io_r_34_b : _GEN_333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_335 = 8'h23 == r_count_0_io_out ? io_r_35_b : _GEN_334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_336 = 8'h24 == r_count_0_io_out ? io_r_36_b : _GEN_335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_337 = 8'h25 == r_count_0_io_out ? io_r_37_b : _GEN_336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_338 = 8'h26 == r_count_0_io_out ? io_r_38_b : _GEN_337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_339 = 8'h27 == r_count_0_io_out ? io_r_39_b : _GEN_338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_340 = 8'h28 == r_count_0_io_out ? io_r_40_b : _GEN_339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_341 = 8'h29 == r_count_0_io_out ? io_r_41_b : _GEN_340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_342 = 8'h2a == r_count_0_io_out ? io_r_42_b : _GEN_341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_343 = 8'h2b == r_count_0_io_out ? io_r_43_b : _GEN_342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_344 = 8'h2c == r_count_0_io_out ? io_r_44_b : _GEN_343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_345 = 8'h2d == r_count_0_io_out ? io_r_45_b : _GEN_344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_346 = 8'h2e == r_count_0_io_out ? io_r_46_b : _GEN_345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_347 = 8'h2f == r_count_0_io_out ? io_r_47_b : _GEN_346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_348 = 8'h30 == r_count_0_io_out ? io_r_48_b : _GEN_347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_349 = 8'h31 == r_count_0_io_out ? io_r_49_b : _GEN_348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_350 = 8'h32 == r_count_0_io_out ? io_r_50_b : _GEN_349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_351 = 8'h33 == r_count_0_io_out ? io_r_51_b : _GEN_350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_352 = 8'h34 == r_count_0_io_out ? io_r_52_b : _GEN_351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_353 = 8'h35 == r_count_0_io_out ? io_r_53_b : _GEN_352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_354 = 8'h36 == r_count_0_io_out ? io_r_54_b : _GEN_353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_355 = 8'h37 == r_count_0_io_out ? io_r_55_b : _GEN_354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_356 = 8'h38 == r_count_0_io_out ? io_r_56_b : _GEN_355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_357 = 8'h39 == r_count_0_io_out ? io_r_57_b : _GEN_356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_358 = 8'h3a == r_count_0_io_out ? io_r_58_b : _GEN_357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_359 = 8'h3b == r_count_0_io_out ? io_r_59_b : _GEN_358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_360 = 8'h3c == r_count_0_io_out ? io_r_60_b : _GEN_359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_361 = 8'h3d == r_count_0_io_out ? io_r_61_b : _GEN_360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_362 = 8'h3e == r_count_0_io_out ? io_r_62_b : _GEN_361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_363 = 8'h3f == r_count_0_io_out ? io_r_63_b : _GEN_362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_364 = 8'h40 == r_count_0_io_out ? io_r_64_b : _GEN_363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_365 = 8'h41 == r_count_0_io_out ? io_r_65_b : _GEN_364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_366 = 8'h42 == r_count_0_io_out ? io_r_66_b : _GEN_365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_367 = 8'h43 == r_count_0_io_out ? io_r_67_b : _GEN_366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_368 = 8'h44 == r_count_0_io_out ? io_r_68_b : _GEN_367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_369 = 8'h45 == r_count_0_io_out ? io_r_69_b : _GEN_368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_370 = 8'h46 == r_count_0_io_out ? io_r_70_b : _GEN_369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_371 = 8'h47 == r_count_0_io_out ? io_r_71_b : _GEN_370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_372 = 8'h48 == r_count_0_io_out ? io_r_72_b : _GEN_371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_373 = 8'h49 == r_count_0_io_out ? io_r_73_b : _GEN_372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_374 = 8'h4a == r_count_0_io_out ? io_r_74_b : _GEN_373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_375 = 8'h4b == r_count_0_io_out ? io_r_75_b : _GEN_374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_376 = 8'h4c == r_count_0_io_out ? io_r_76_b : _GEN_375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_377 = 8'h4d == r_count_0_io_out ? io_r_77_b : _GEN_376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_378 = 8'h4e == r_count_0_io_out ? io_r_78_b : _GEN_377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_379 = 8'h4f == r_count_0_io_out ? io_r_79_b : _GEN_378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_380 = 8'h50 == r_count_0_io_out ? io_r_80_b : _GEN_379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_381 = 8'h51 == r_count_0_io_out ? io_r_81_b : _GEN_380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_382 = 8'h52 == r_count_0_io_out ? io_r_82_b : _GEN_381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_383 = 8'h53 == r_count_0_io_out ? io_r_83_b : _GEN_382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_384 = 8'h54 == r_count_0_io_out ? io_r_84_b : _GEN_383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_385 = 8'h55 == r_count_0_io_out ? io_r_85_b : _GEN_384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_386 = 8'h56 == r_count_0_io_out ? io_r_86_b : _GEN_385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_387 = 8'h57 == r_count_0_io_out ? io_r_87_b : _GEN_386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_388 = 8'h58 == r_count_0_io_out ? io_r_88_b : _GEN_387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_389 = 8'h59 == r_count_0_io_out ? io_r_89_b : _GEN_388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_390 = 8'h5a == r_count_0_io_out ? io_r_90_b : _GEN_389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_391 = 8'h5b == r_count_0_io_out ? io_r_91_b : _GEN_390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_392 = 8'h5c == r_count_0_io_out ? io_r_92_b : _GEN_391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_393 = 8'h5d == r_count_0_io_out ? io_r_93_b : _GEN_392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_394 = 8'h5e == r_count_0_io_out ? io_r_94_b : _GEN_393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_395 = 8'h5f == r_count_0_io_out ? io_r_95_b : _GEN_394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_396 = 8'h60 == r_count_0_io_out ? io_r_96_b : _GEN_395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_397 = 8'h61 == r_count_0_io_out ? io_r_97_b : _GEN_396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_398 = 8'h62 == r_count_0_io_out ? io_r_98_b : _GEN_397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_399 = 8'h63 == r_count_0_io_out ? io_r_99_b : _GEN_398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_400 = 8'h64 == r_count_0_io_out ? io_r_100_b : _GEN_399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_401 = 8'h65 == r_count_0_io_out ? io_r_101_b : _GEN_400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_402 = 8'h66 == r_count_0_io_out ? io_r_102_b : _GEN_401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_403 = 8'h67 == r_count_0_io_out ? io_r_103_b : _GEN_402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_404 = 8'h68 == r_count_0_io_out ? io_r_104_b : _GEN_403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_405 = 8'h69 == r_count_0_io_out ? io_r_105_b : _GEN_404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_406 = 8'h6a == r_count_0_io_out ? io_r_106_b : _GEN_405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_407 = 8'h6b == r_count_0_io_out ? io_r_107_b : _GEN_406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_408 = 8'h6c == r_count_0_io_out ? io_r_108_b : _GEN_407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_409 = 8'h6d == r_count_0_io_out ? io_r_109_b : _GEN_408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_410 = 8'h6e == r_count_0_io_out ? io_r_110_b : _GEN_409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_411 = 8'h6f == r_count_0_io_out ? io_r_111_b : _GEN_410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_412 = 8'h70 == r_count_0_io_out ? io_r_112_b : _GEN_411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_413 = 8'h71 == r_count_0_io_out ? io_r_113_b : _GEN_412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_414 = 8'h72 == r_count_0_io_out ? io_r_114_b : _GEN_413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_415 = 8'h73 == r_count_0_io_out ? io_r_115_b : _GEN_414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_416 = 8'h74 == r_count_0_io_out ? io_r_116_b : _GEN_415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_417 = 8'h75 == r_count_0_io_out ? io_r_117_b : _GEN_416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_418 = 8'h76 == r_count_0_io_out ? io_r_118_b : _GEN_417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_419 = 8'h77 == r_count_0_io_out ? io_r_119_b : _GEN_418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_420 = 8'h78 == r_count_0_io_out ? io_r_120_b : _GEN_419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_421 = 8'h79 == r_count_0_io_out ? io_r_121_b : _GEN_420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_422 = 8'h7a == r_count_0_io_out ? io_r_122_b : _GEN_421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_423 = 8'h7b == r_count_0_io_out ? io_r_123_b : _GEN_422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_424 = 8'h7c == r_count_0_io_out ? io_r_124_b : _GEN_423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_425 = 8'h7d == r_count_0_io_out ? io_r_125_b : _GEN_424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_426 = 8'h7e == r_count_0_io_out ? io_r_126_b : _GEN_425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_427 = 8'h7f == r_count_0_io_out ? io_r_127_b : _GEN_426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_428 = 8'h80 == r_count_0_io_out ? io_r_128_b : _GEN_427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_429 = 8'h81 == r_count_0_io_out ? io_r_129_b : _GEN_428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_430 = 8'h82 == r_count_0_io_out ? io_r_130_b : _GEN_429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_431 = 8'h83 == r_count_0_io_out ? io_r_131_b : _GEN_430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_432 = 8'h84 == r_count_0_io_out ? io_r_132_b : _GEN_431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_433 = 8'h85 == r_count_0_io_out ? io_r_133_b : _GEN_432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_434 = 8'h86 == r_count_0_io_out ? io_r_134_b : _GEN_433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_435 = 8'h87 == r_count_0_io_out ? io_r_135_b : _GEN_434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_436 = 8'h88 == r_count_0_io_out ? io_r_136_b : _GEN_435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_437 = 8'h89 == r_count_0_io_out ? io_r_137_b : _GEN_436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_438 = 8'h8a == r_count_0_io_out ? io_r_138_b : _GEN_437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_439 = 8'h8b == r_count_0_io_out ? io_r_139_b : _GEN_438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_440 = 8'h8c == r_count_0_io_out ? io_r_140_b : _GEN_439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_441 = 8'h8d == r_count_0_io_out ? io_r_141_b : _GEN_440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_442 = 8'h8e == r_count_0_io_out ? io_r_142_b : _GEN_441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_443 = 8'h8f == r_count_0_io_out ? io_r_143_b : _GEN_442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_444 = 8'h90 == r_count_0_io_out ? io_r_144_b : _GEN_443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_445 = 8'h91 == r_count_0_io_out ? io_r_145_b : _GEN_444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_446 = 8'h92 == r_count_0_io_out ? io_r_146_b : _GEN_445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_447 = 8'h93 == r_count_0_io_out ? io_r_147_b : _GEN_446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_448 = 8'h94 == r_count_0_io_out ? io_r_148_b : _GEN_447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_449 = 8'h95 == r_count_0_io_out ? io_r_149_b : _GEN_448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_450 = 8'h96 == r_count_0_io_out ? io_r_150_b : _GEN_449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_451 = 8'h97 == r_count_0_io_out ? io_r_151_b : _GEN_450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_452 = 8'h98 == r_count_0_io_out ? io_r_152_b : _GEN_451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_453 = 8'h99 == r_count_0_io_out ? io_r_153_b : _GEN_452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_454 = 8'h9a == r_count_0_io_out ? io_r_154_b : _GEN_453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_455 = 8'h9b == r_count_0_io_out ? io_r_155_b : _GEN_454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_456 = 8'h9c == r_count_0_io_out ? io_r_156_b : _GEN_455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_457 = 8'h9d == r_count_0_io_out ? io_r_157_b : _GEN_456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_458 = 8'h9e == r_count_0_io_out ? io_r_158_b : _GEN_457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_459 = 8'h9f == r_count_0_io_out ? io_r_159_b : _GEN_458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_460 = 8'ha0 == r_count_0_io_out ? io_r_160_b : _GEN_459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_461 = 8'ha1 == r_count_0_io_out ? io_r_161_b : _GEN_460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_462 = 8'ha2 == r_count_0_io_out ? io_r_162_b : _GEN_461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_463 = 8'ha3 == r_count_0_io_out ? io_r_163_b : _GEN_462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_464 = 8'ha4 == r_count_0_io_out ? io_r_164_b : _GEN_463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_465 = 8'ha5 == r_count_0_io_out ? io_r_165_b : _GEN_464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_466 = 8'ha6 == r_count_0_io_out ? io_r_166_b : _GEN_465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_467 = 8'ha7 == r_count_0_io_out ? io_r_167_b : _GEN_466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_468 = 8'ha8 == r_count_0_io_out ? io_r_168_b : _GEN_467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_469 = 8'ha9 == r_count_0_io_out ? io_r_169_b : _GEN_468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_470 = 8'haa == r_count_0_io_out ? io_r_170_b : _GEN_469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_471 = 8'hab == r_count_0_io_out ? io_r_171_b : _GEN_470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_472 = 8'hac == r_count_0_io_out ? io_r_172_b : _GEN_471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_473 = 8'had == r_count_0_io_out ? io_r_173_b : _GEN_472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_474 = 8'hae == r_count_0_io_out ? io_r_174_b : _GEN_473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_475 = 8'haf == r_count_0_io_out ? io_r_175_b : _GEN_474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_476 = 8'hb0 == r_count_0_io_out ? io_r_176_b : _GEN_475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_477 = 8'hb1 == r_count_0_io_out ? io_r_177_b : _GEN_476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_478 = 8'hb2 == r_count_0_io_out ? io_r_178_b : _GEN_477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_479 = 8'hb3 == r_count_0_io_out ? io_r_179_b : _GEN_478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_480 = 8'hb4 == r_count_0_io_out ? io_r_180_b : _GEN_479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_481 = 8'hb5 == r_count_0_io_out ? io_r_181_b : _GEN_480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_482 = 8'hb6 == r_count_0_io_out ? io_r_182_b : _GEN_481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_483 = 8'hb7 == r_count_0_io_out ? io_r_183_b : _GEN_482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_484 = 8'hb8 == r_count_0_io_out ? io_r_184_b : _GEN_483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_485 = 8'hb9 == r_count_0_io_out ? io_r_185_b : _GEN_484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_486 = 8'hba == r_count_0_io_out ? io_r_186_b : _GEN_485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_487 = 8'hbb == r_count_0_io_out ? io_r_187_b : _GEN_486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_488 = 8'hbc == r_count_0_io_out ? io_r_188_b : _GEN_487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_489 = 8'hbd == r_count_0_io_out ? io_r_189_b : _GEN_488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_490 = 8'hbe == r_count_0_io_out ? io_r_190_b : _GEN_489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_491 = 8'hbf == r_count_0_io_out ? io_r_191_b : _GEN_490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_492 = 8'hc0 == r_count_0_io_out ? io_r_192_b : _GEN_491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_493 = 8'hc1 == r_count_0_io_out ? io_r_193_b : _GEN_492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_494 = 8'hc2 == r_count_0_io_out ? io_r_194_b : _GEN_493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_495 = 8'hc3 == r_count_0_io_out ? io_r_195_b : _GEN_494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_496 = 8'hc4 == r_count_0_io_out ? io_r_196_b : _GEN_495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_497 = 8'hc5 == r_count_0_io_out ? io_r_197_b : _GEN_496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_498 = 8'hc6 == r_count_0_io_out ? io_r_198_b : _GEN_497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_501 = 8'h1 == r_count_1_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_502 = 8'h2 == r_count_1_io_out ? io_r_2_b : _GEN_501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_503 = 8'h3 == r_count_1_io_out ? io_r_3_b : _GEN_502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_504 = 8'h4 == r_count_1_io_out ? io_r_4_b : _GEN_503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_505 = 8'h5 == r_count_1_io_out ? io_r_5_b : _GEN_504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_506 = 8'h6 == r_count_1_io_out ? io_r_6_b : _GEN_505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_507 = 8'h7 == r_count_1_io_out ? io_r_7_b : _GEN_506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_508 = 8'h8 == r_count_1_io_out ? io_r_8_b : _GEN_507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_509 = 8'h9 == r_count_1_io_out ? io_r_9_b : _GEN_508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_510 = 8'ha == r_count_1_io_out ? io_r_10_b : _GEN_509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_511 = 8'hb == r_count_1_io_out ? io_r_11_b : _GEN_510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_512 = 8'hc == r_count_1_io_out ? io_r_12_b : _GEN_511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_513 = 8'hd == r_count_1_io_out ? io_r_13_b : _GEN_512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_514 = 8'he == r_count_1_io_out ? io_r_14_b : _GEN_513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_515 = 8'hf == r_count_1_io_out ? io_r_15_b : _GEN_514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_516 = 8'h10 == r_count_1_io_out ? io_r_16_b : _GEN_515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_517 = 8'h11 == r_count_1_io_out ? io_r_17_b : _GEN_516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_518 = 8'h12 == r_count_1_io_out ? io_r_18_b : _GEN_517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_519 = 8'h13 == r_count_1_io_out ? io_r_19_b : _GEN_518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_520 = 8'h14 == r_count_1_io_out ? io_r_20_b : _GEN_519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_521 = 8'h15 == r_count_1_io_out ? io_r_21_b : _GEN_520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_522 = 8'h16 == r_count_1_io_out ? io_r_22_b : _GEN_521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_523 = 8'h17 == r_count_1_io_out ? io_r_23_b : _GEN_522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_524 = 8'h18 == r_count_1_io_out ? io_r_24_b : _GEN_523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_525 = 8'h19 == r_count_1_io_out ? io_r_25_b : _GEN_524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_526 = 8'h1a == r_count_1_io_out ? io_r_26_b : _GEN_525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_527 = 8'h1b == r_count_1_io_out ? io_r_27_b : _GEN_526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_528 = 8'h1c == r_count_1_io_out ? io_r_28_b : _GEN_527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_529 = 8'h1d == r_count_1_io_out ? io_r_29_b : _GEN_528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_530 = 8'h1e == r_count_1_io_out ? io_r_30_b : _GEN_529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_531 = 8'h1f == r_count_1_io_out ? io_r_31_b : _GEN_530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_532 = 8'h20 == r_count_1_io_out ? io_r_32_b : _GEN_531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_533 = 8'h21 == r_count_1_io_out ? io_r_33_b : _GEN_532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_534 = 8'h22 == r_count_1_io_out ? io_r_34_b : _GEN_533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_535 = 8'h23 == r_count_1_io_out ? io_r_35_b : _GEN_534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_536 = 8'h24 == r_count_1_io_out ? io_r_36_b : _GEN_535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_537 = 8'h25 == r_count_1_io_out ? io_r_37_b : _GEN_536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_538 = 8'h26 == r_count_1_io_out ? io_r_38_b : _GEN_537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_539 = 8'h27 == r_count_1_io_out ? io_r_39_b : _GEN_538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_540 = 8'h28 == r_count_1_io_out ? io_r_40_b : _GEN_539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_541 = 8'h29 == r_count_1_io_out ? io_r_41_b : _GEN_540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_542 = 8'h2a == r_count_1_io_out ? io_r_42_b : _GEN_541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_543 = 8'h2b == r_count_1_io_out ? io_r_43_b : _GEN_542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_544 = 8'h2c == r_count_1_io_out ? io_r_44_b : _GEN_543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_545 = 8'h2d == r_count_1_io_out ? io_r_45_b : _GEN_544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_546 = 8'h2e == r_count_1_io_out ? io_r_46_b : _GEN_545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_547 = 8'h2f == r_count_1_io_out ? io_r_47_b : _GEN_546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_548 = 8'h30 == r_count_1_io_out ? io_r_48_b : _GEN_547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_549 = 8'h31 == r_count_1_io_out ? io_r_49_b : _GEN_548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_550 = 8'h32 == r_count_1_io_out ? io_r_50_b : _GEN_549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_551 = 8'h33 == r_count_1_io_out ? io_r_51_b : _GEN_550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_552 = 8'h34 == r_count_1_io_out ? io_r_52_b : _GEN_551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_553 = 8'h35 == r_count_1_io_out ? io_r_53_b : _GEN_552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_554 = 8'h36 == r_count_1_io_out ? io_r_54_b : _GEN_553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_555 = 8'h37 == r_count_1_io_out ? io_r_55_b : _GEN_554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_556 = 8'h38 == r_count_1_io_out ? io_r_56_b : _GEN_555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_557 = 8'h39 == r_count_1_io_out ? io_r_57_b : _GEN_556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_558 = 8'h3a == r_count_1_io_out ? io_r_58_b : _GEN_557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_559 = 8'h3b == r_count_1_io_out ? io_r_59_b : _GEN_558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_560 = 8'h3c == r_count_1_io_out ? io_r_60_b : _GEN_559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_561 = 8'h3d == r_count_1_io_out ? io_r_61_b : _GEN_560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_562 = 8'h3e == r_count_1_io_out ? io_r_62_b : _GEN_561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_563 = 8'h3f == r_count_1_io_out ? io_r_63_b : _GEN_562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_564 = 8'h40 == r_count_1_io_out ? io_r_64_b : _GEN_563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_565 = 8'h41 == r_count_1_io_out ? io_r_65_b : _GEN_564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_566 = 8'h42 == r_count_1_io_out ? io_r_66_b : _GEN_565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_567 = 8'h43 == r_count_1_io_out ? io_r_67_b : _GEN_566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_568 = 8'h44 == r_count_1_io_out ? io_r_68_b : _GEN_567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_569 = 8'h45 == r_count_1_io_out ? io_r_69_b : _GEN_568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_570 = 8'h46 == r_count_1_io_out ? io_r_70_b : _GEN_569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_571 = 8'h47 == r_count_1_io_out ? io_r_71_b : _GEN_570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_572 = 8'h48 == r_count_1_io_out ? io_r_72_b : _GEN_571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_573 = 8'h49 == r_count_1_io_out ? io_r_73_b : _GEN_572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_574 = 8'h4a == r_count_1_io_out ? io_r_74_b : _GEN_573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_575 = 8'h4b == r_count_1_io_out ? io_r_75_b : _GEN_574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_576 = 8'h4c == r_count_1_io_out ? io_r_76_b : _GEN_575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_577 = 8'h4d == r_count_1_io_out ? io_r_77_b : _GEN_576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_578 = 8'h4e == r_count_1_io_out ? io_r_78_b : _GEN_577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_579 = 8'h4f == r_count_1_io_out ? io_r_79_b : _GEN_578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_580 = 8'h50 == r_count_1_io_out ? io_r_80_b : _GEN_579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_581 = 8'h51 == r_count_1_io_out ? io_r_81_b : _GEN_580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_582 = 8'h52 == r_count_1_io_out ? io_r_82_b : _GEN_581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_583 = 8'h53 == r_count_1_io_out ? io_r_83_b : _GEN_582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_584 = 8'h54 == r_count_1_io_out ? io_r_84_b : _GEN_583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_585 = 8'h55 == r_count_1_io_out ? io_r_85_b : _GEN_584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_586 = 8'h56 == r_count_1_io_out ? io_r_86_b : _GEN_585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_587 = 8'h57 == r_count_1_io_out ? io_r_87_b : _GEN_586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_588 = 8'h58 == r_count_1_io_out ? io_r_88_b : _GEN_587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_589 = 8'h59 == r_count_1_io_out ? io_r_89_b : _GEN_588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_590 = 8'h5a == r_count_1_io_out ? io_r_90_b : _GEN_589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_591 = 8'h5b == r_count_1_io_out ? io_r_91_b : _GEN_590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_592 = 8'h5c == r_count_1_io_out ? io_r_92_b : _GEN_591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_593 = 8'h5d == r_count_1_io_out ? io_r_93_b : _GEN_592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_594 = 8'h5e == r_count_1_io_out ? io_r_94_b : _GEN_593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_595 = 8'h5f == r_count_1_io_out ? io_r_95_b : _GEN_594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_596 = 8'h60 == r_count_1_io_out ? io_r_96_b : _GEN_595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_597 = 8'h61 == r_count_1_io_out ? io_r_97_b : _GEN_596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_598 = 8'h62 == r_count_1_io_out ? io_r_98_b : _GEN_597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_599 = 8'h63 == r_count_1_io_out ? io_r_99_b : _GEN_598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_600 = 8'h64 == r_count_1_io_out ? io_r_100_b : _GEN_599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_601 = 8'h65 == r_count_1_io_out ? io_r_101_b : _GEN_600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_602 = 8'h66 == r_count_1_io_out ? io_r_102_b : _GEN_601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_603 = 8'h67 == r_count_1_io_out ? io_r_103_b : _GEN_602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_604 = 8'h68 == r_count_1_io_out ? io_r_104_b : _GEN_603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_605 = 8'h69 == r_count_1_io_out ? io_r_105_b : _GEN_604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_606 = 8'h6a == r_count_1_io_out ? io_r_106_b : _GEN_605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_607 = 8'h6b == r_count_1_io_out ? io_r_107_b : _GEN_606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_608 = 8'h6c == r_count_1_io_out ? io_r_108_b : _GEN_607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_609 = 8'h6d == r_count_1_io_out ? io_r_109_b : _GEN_608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_610 = 8'h6e == r_count_1_io_out ? io_r_110_b : _GEN_609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_611 = 8'h6f == r_count_1_io_out ? io_r_111_b : _GEN_610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_612 = 8'h70 == r_count_1_io_out ? io_r_112_b : _GEN_611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_613 = 8'h71 == r_count_1_io_out ? io_r_113_b : _GEN_612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_614 = 8'h72 == r_count_1_io_out ? io_r_114_b : _GEN_613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_615 = 8'h73 == r_count_1_io_out ? io_r_115_b : _GEN_614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_616 = 8'h74 == r_count_1_io_out ? io_r_116_b : _GEN_615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_617 = 8'h75 == r_count_1_io_out ? io_r_117_b : _GEN_616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_618 = 8'h76 == r_count_1_io_out ? io_r_118_b : _GEN_617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_619 = 8'h77 == r_count_1_io_out ? io_r_119_b : _GEN_618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_620 = 8'h78 == r_count_1_io_out ? io_r_120_b : _GEN_619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_621 = 8'h79 == r_count_1_io_out ? io_r_121_b : _GEN_620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_622 = 8'h7a == r_count_1_io_out ? io_r_122_b : _GEN_621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_623 = 8'h7b == r_count_1_io_out ? io_r_123_b : _GEN_622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_624 = 8'h7c == r_count_1_io_out ? io_r_124_b : _GEN_623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_625 = 8'h7d == r_count_1_io_out ? io_r_125_b : _GEN_624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_626 = 8'h7e == r_count_1_io_out ? io_r_126_b : _GEN_625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_627 = 8'h7f == r_count_1_io_out ? io_r_127_b : _GEN_626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_628 = 8'h80 == r_count_1_io_out ? io_r_128_b : _GEN_627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_629 = 8'h81 == r_count_1_io_out ? io_r_129_b : _GEN_628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_630 = 8'h82 == r_count_1_io_out ? io_r_130_b : _GEN_629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_631 = 8'h83 == r_count_1_io_out ? io_r_131_b : _GEN_630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_632 = 8'h84 == r_count_1_io_out ? io_r_132_b : _GEN_631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_633 = 8'h85 == r_count_1_io_out ? io_r_133_b : _GEN_632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_634 = 8'h86 == r_count_1_io_out ? io_r_134_b : _GEN_633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_635 = 8'h87 == r_count_1_io_out ? io_r_135_b : _GEN_634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_636 = 8'h88 == r_count_1_io_out ? io_r_136_b : _GEN_635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_637 = 8'h89 == r_count_1_io_out ? io_r_137_b : _GEN_636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_638 = 8'h8a == r_count_1_io_out ? io_r_138_b : _GEN_637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_639 = 8'h8b == r_count_1_io_out ? io_r_139_b : _GEN_638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_640 = 8'h8c == r_count_1_io_out ? io_r_140_b : _GEN_639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_641 = 8'h8d == r_count_1_io_out ? io_r_141_b : _GEN_640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_642 = 8'h8e == r_count_1_io_out ? io_r_142_b : _GEN_641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_643 = 8'h8f == r_count_1_io_out ? io_r_143_b : _GEN_642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_644 = 8'h90 == r_count_1_io_out ? io_r_144_b : _GEN_643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_645 = 8'h91 == r_count_1_io_out ? io_r_145_b : _GEN_644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_646 = 8'h92 == r_count_1_io_out ? io_r_146_b : _GEN_645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_647 = 8'h93 == r_count_1_io_out ? io_r_147_b : _GEN_646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_648 = 8'h94 == r_count_1_io_out ? io_r_148_b : _GEN_647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_649 = 8'h95 == r_count_1_io_out ? io_r_149_b : _GEN_648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_650 = 8'h96 == r_count_1_io_out ? io_r_150_b : _GEN_649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_651 = 8'h97 == r_count_1_io_out ? io_r_151_b : _GEN_650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_652 = 8'h98 == r_count_1_io_out ? io_r_152_b : _GEN_651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_653 = 8'h99 == r_count_1_io_out ? io_r_153_b : _GEN_652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_654 = 8'h9a == r_count_1_io_out ? io_r_154_b : _GEN_653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_655 = 8'h9b == r_count_1_io_out ? io_r_155_b : _GEN_654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_656 = 8'h9c == r_count_1_io_out ? io_r_156_b : _GEN_655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_657 = 8'h9d == r_count_1_io_out ? io_r_157_b : _GEN_656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_658 = 8'h9e == r_count_1_io_out ? io_r_158_b : _GEN_657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_659 = 8'h9f == r_count_1_io_out ? io_r_159_b : _GEN_658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_660 = 8'ha0 == r_count_1_io_out ? io_r_160_b : _GEN_659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_661 = 8'ha1 == r_count_1_io_out ? io_r_161_b : _GEN_660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_662 = 8'ha2 == r_count_1_io_out ? io_r_162_b : _GEN_661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_663 = 8'ha3 == r_count_1_io_out ? io_r_163_b : _GEN_662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_664 = 8'ha4 == r_count_1_io_out ? io_r_164_b : _GEN_663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_665 = 8'ha5 == r_count_1_io_out ? io_r_165_b : _GEN_664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_666 = 8'ha6 == r_count_1_io_out ? io_r_166_b : _GEN_665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_667 = 8'ha7 == r_count_1_io_out ? io_r_167_b : _GEN_666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_668 = 8'ha8 == r_count_1_io_out ? io_r_168_b : _GEN_667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_669 = 8'ha9 == r_count_1_io_out ? io_r_169_b : _GEN_668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_670 = 8'haa == r_count_1_io_out ? io_r_170_b : _GEN_669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_671 = 8'hab == r_count_1_io_out ? io_r_171_b : _GEN_670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_672 = 8'hac == r_count_1_io_out ? io_r_172_b : _GEN_671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_673 = 8'had == r_count_1_io_out ? io_r_173_b : _GEN_672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_674 = 8'hae == r_count_1_io_out ? io_r_174_b : _GEN_673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_675 = 8'haf == r_count_1_io_out ? io_r_175_b : _GEN_674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_676 = 8'hb0 == r_count_1_io_out ? io_r_176_b : _GEN_675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_677 = 8'hb1 == r_count_1_io_out ? io_r_177_b : _GEN_676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_678 = 8'hb2 == r_count_1_io_out ? io_r_178_b : _GEN_677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_679 = 8'hb3 == r_count_1_io_out ? io_r_179_b : _GEN_678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_680 = 8'hb4 == r_count_1_io_out ? io_r_180_b : _GEN_679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_681 = 8'hb5 == r_count_1_io_out ? io_r_181_b : _GEN_680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_682 = 8'hb6 == r_count_1_io_out ? io_r_182_b : _GEN_681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_683 = 8'hb7 == r_count_1_io_out ? io_r_183_b : _GEN_682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_684 = 8'hb8 == r_count_1_io_out ? io_r_184_b : _GEN_683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_685 = 8'hb9 == r_count_1_io_out ? io_r_185_b : _GEN_684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_686 = 8'hba == r_count_1_io_out ? io_r_186_b : _GEN_685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_687 = 8'hbb == r_count_1_io_out ? io_r_187_b : _GEN_686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_688 = 8'hbc == r_count_1_io_out ? io_r_188_b : _GEN_687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_689 = 8'hbd == r_count_1_io_out ? io_r_189_b : _GEN_688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_690 = 8'hbe == r_count_1_io_out ? io_r_190_b : _GEN_689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_691 = 8'hbf == r_count_1_io_out ? io_r_191_b : _GEN_690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_692 = 8'hc0 == r_count_1_io_out ? io_r_192_b : _GEN_691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_693 = 8'hc1 == r_count_1_io_out ? io_r_193_b : _GEN_692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_694 = 8'hc2 == r_count_1_io_out ? io_r_194_b : _GEN_693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_695 = 8'hc3 == r_count_1_io_out ? io_r_195_b : _GEN_694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_696 = 8'hc4 == r_count_1_io_out ? io_r_196_b : _GEN_695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_697 = 8'hc5 == r_count_1_io_out ? io_r_197_b : _GEN_696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_698 = 8'hc6 == r_count_1_io_out ? io_r_198_b : _GEN_697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_701 = 8'h1 == r_count_2_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_702 = 8'h2 == r_count_2_io_out ? io_r_2_b : _GEN_701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_703 = 8'h3 == r_count_2_io_out ? io_r_3_b : _GEN_702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_704 = 8'h4 == r_count_2_io_out ? io_r_4_b : _GEN_703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_705 = 8'h5 == r_count_2_io_out ? io_r_5_b : _GEN_704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_706 = 8'h6 == r_count_2_io_out ? io_r_6_b : _GEN_705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_707 = 8'h7 == r_count_2_io_out ? io_r_7_b : _GEN_706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_708 = 8'h8 == r_count_2_io_out ? io_r_8_b : _GEN_707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_709 = 8'h9 == r_count_2_io_out ? io_r_9_b : _GEN_708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_710 = 8'ha == r_count_2_io_out ? io_r_10_b : _GEN_709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_711 = 8'hb == r_count_2_io_out ? io_r_11_b : _GEN_710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_712 = 8'hc == r_count_2_io_out ? io_r_12_b : _GEN_711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_713 = 8'hd == r_count_2_io_out ? io_r_13_b : _GEN_712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_714 = 8'he == r_count_2_io_out ? io_r_14_b : _GEN_713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_715 = 8'hf == r_count_2_io_out ? io_r_15_b : _GEN_714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_716 = 8'h10 == r_count_2_io_out ? io_r_16_b : _GEN_715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_717 = 8'h11 == r_count_2_io_out ? io_r_17_b : _GEN_716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_718 = 8'h12 == r_count_2_io_out ? io_r_18_b : _GEN_717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_719 = 8'h13 == r_count_2_io_out ? io_r_19_b : _GEN_718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_720 = 8'h14 == r_count_2_io_out ? io_r_20_b : _GEN_719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_721 = 8'h15 == r_count_2_io_out ? io_r_21_b : _GEN_720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_722 = 8'h16 == r_count_2_io_out ? io_r_22_b : _GEN_721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_723 = 8'h17 == r_count_2_io_out ? io_r_23_b : _GEN_722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_724 = 8'h18 == r_count_2_io_out ? io_r_24_b : _GEN_723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_725 = 8'h19 == r_count_2_io_out ? io_r_25_b : _GEN_724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_726 = 8'h1a == r_count_2_io_out ? io_r_26_b : _GEN_725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_727 = 8'h1b == r_count_2_io_out ? io_r_27_b : _GEN_726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_728 = 8'h1c == r_count_2_io_out ? io_r_28_b : _GEN_727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_729 = 8'h1d == r_count_2_io_out ? io_r_29_b : _GEN_728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_730 = 8'h1e == r_count_2_io_out ? io_r_30_b : _GEN_729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_731 = 8'h1f == r_count_2_io_out ? io_r_31_b : _GEN_730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_732 = 8'h20 == r_count_2_io_out ? io_r_32_b : _GEN_731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_733 = 8'h21 == r_count_2_io_out ? io_r_33_b : _GEN_732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_734 = 8'h22 == r_count_2_io_out ? io_r_34_b : _GEN_733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_735 = 8'h23 == r_count_2_io_out ? io_r_35_b : _GEN_734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_736 = 8'h24 == r_count_2_io_out ? io_r_36_b : _GEN_735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_737 = 8'h25 == r_count_2_io_out ? io_r_37_b : _GEN_736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_738 = 8'h26 == r_count_2_io_out ? io_r_38_b : _GEN_737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_739 = 8'h27 == r_count_2_io_out ? io_r_39_b : _GEN_738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_740 = 8'h28 == r_count_2_io_out ? io_r_40_b : _GEN_739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_741 = 8'h29 == r_count_2_io_out ? io_r_41_b : _GEN_740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_742 = 8'h2a == r_count_2_io_out ? io_r_42_b : _GEN_741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_743 = 8'h2b == r_count_2_io_out ? io_r_43_b : _GEN_742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_744 = 8'h2c == r_count_2_io_out ? io_r_44_b : _GEN_743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_745 = 8'h2d == r_count_2_io_out ? io_r_45_b : _GEN_744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_746 = 8'h2e == r_count_2_io_out ? io_r_46_b : _GEN_745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_747 = 8'h2f == r_count_2_io_out ? io_r_47_b : _GEN_746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_748 = 8'h30 == r_count_2_io_out ? io_r_48_b : _GEN_747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_749 = 8'h31 == r_count_2_io_out ? io_r_49_b : _GEN_748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_750 = 8'h32 == r_count_2_io_out ? io_r_50_b : _GEN_749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_751 = 8'h33 == r_count_2_io_out ? io_r_51_b : _GEN_750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_752 = 8'h34 == r_count_2_io_out ? io_r_52_b : _GEN_751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_753 = 8'h35 == r_count_2_io_out ? io_r_53_b : _GEN_752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_754 = 8'h36 == r_count_2_io_out ? io_r_54_b : _GEN_753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_755 = 8'h37 == r_count_2_io_out ? io_r_55_b : _GEN_754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_756 = 8'h38 == r_count_2_io_out ? io_r_56_b : _GEN_755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_757 = 8'h39 == r_count_2_io_out ? io_r_57_b : _GEN_756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_758 = 8'h3a == r_count_2_io_out ? io_r_58_b : _GEN_757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_759 = 8'h3b == r_count_2_io_out ? io_r_59_b : _GEN_758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_760 = 8'h3c == r_count_2_io_out ? io_r_60_b : _GEN_759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_761 = 8'h3d == r_count_2_io_out ? io_r_61_b : _GEN_760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_762 = 8'h3e == r_count_2_io_out ? io_r_62_b : _GEN_761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_763 = 8'h3f == r_count_2_io_out ? io_r_63_b : _GEN_762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_764 = 8'h40 == r_count_2_io_out ? io_r_64_b : _GEN_763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_765 = 8'h41 == r_count_2_io_out ? io_r_65_b : _GEN_764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_766 = 8'h42 == r_count_2_io_out ? io_r_66_b : _GEN_765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_767 = 8'h43 == r_count_2_io_out ? io_r_67_b : _GEN_766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_768 = 8'h44 == r_count_2_io_out ? io_r_68_b : _GEN_767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_769 = 8'h45 == r_count_2_io_out ? io_r_69_b : _GEN_768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_770 = 8'h46 == r_count_2_io_out ? io_r_70_b : _GEN_769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_771 = 8'h47 == r_count_2_io_out ? io_r_71_b : _GEN_770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_772 = 8'h48 == r_count_2_io_out ? io_r_72_b : _GEN_771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_773 = 8'h49 == r_count_2_io_out ? io_r_73_b : _GEN_772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_774 = 8'h4a == r_count_2_io_out ? io_r_74_b : _GEN_773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_775 = 8'h4b == r_count_2_io_out ? io_r_75_b : _GEN_774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_776 = 8'h4c == r_count_2_io_out ? io_r_76_b : _GEN_775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_777 = 8'h4d == r_count_2_io_out ? io_r_77_b : _GEN_776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_778 = 8'h4e == r_count_2_io_out ? io_r_78_b : _GEN_777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_779 = 8'h4f == r_count_2_io_out ? io_r_79_b : _GEN_778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_780 = 8'h50 == r_count_2_io_out ? io_r_80_b : _GEN_779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_781 = 8'h51 == r_count_2_io_out ? io_r_81_b : _GEN_780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_782 = 8'h52 == r_count_2_io_out ? io_r_82_b : _GEN_781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_783 = 8'h53 == r_count_2_io_out ? io_r_83_b : _GEN_782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_784 = 8'h54 == r_count_2_io_out ? io_r_84_b : _GEN_783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_785 = 8'h55 == r_count_2_io_out ? io_r_85_b : _GEN_784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_786 = 8'h56 == r_count_2_io_out ? io_r_86_b : _GEN_785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_787 = 8'h57 == r_count_2_io_out ? io_r_87_b : _GEN_786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_788 = 8'h58 == r_count_2_io_out ? io_r_88_b : _GEN_787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_789 = 8'h59 == r_count_2_io_out ? io_r_89_b : _GEN_788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_790 = 8'h5a == r_count_2_io_out ? io_r_90_b : _GEN_789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_791 = 8'h5b == r_count_2_io_out ? io_r_91_b : _GEN_790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_792 = 8'h5c == r_count_2_io_out ? io_r_92_b : _GEN_791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_793 = 8'h5d == r_count_2_io_out ? io_r_93_b : _GEN_792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_794 = 8'h5e == r_count_2_io_out ? io_r_94_b : _GEN_793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_795 = 8'h5f == r_count_2_io_out ? io_r_95_b : _GEN_794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_796 = 8'h60 == r_count_2_io_out ? io_r_96_b : _GEN_795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_797 = 8'h61 == r_count_2_io_out ? io_r_97_b : _GEN_796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_798 = 8'h62 == r_count_2_io_out ? io_r_98_b : _GEN_797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_799 = 8'h63 == r_count_2_io_out ? io_r_99_b : _GEN_798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_800 = 8'h64 == r_count_2_io_out ? io_r_100_b : _GEN_799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_801 = 8'h65 == r_count_2_io_out ? io_r_101_b : _GEN_800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_802 = 8'h66 == r_count_2_io_out ? io_r_102_b : _GEN_801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_803 = 8'h67 == r_count_2_io_out ? io_r_103_b : _GEN_802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_804 = 8'h68 == r_count_2_io_out ? io_r_104_b : _GEN_803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_805 = 8'h69 == r_count_2_io_out ? io_r_105_b : _GEN_804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_806 = 8'h6a == r_count_2_io_out ? io_r_106_b : _GEN_805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_807 = 8'h6b == r_count_2_io_out ? io_r_107_b : _GEN_806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_808 = 8'h6c == r_count_2_io_out ? io_r_108_b : _GEN_807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_809 = 8'h6d == r_count_2_io_out ? io_r_109_b : _GEN_808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_810 = 8'h6e == r_count_2_io_out ? io_r_110_b : _GEN_809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_811 = 8'h6f == r_count_2_io_out ? io_r_111_b : _GEN_810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_812 = 8'h70 == r_count_2_io_out ? io_r_112_b : _GEN_811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_813 = 8'h71 == r_count_2_io_out ? io_r_113_b : _GEN_812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_814 = 8'h72 == r_count_2_io_out ? io_r_114_b : _GEN_813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_815 = 8'h73 == r_count_2_io_out ? io_r_115_b : _GEN_814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_816 = 8'h74 == r_count_2_io_out ? io_r_116_b : _GEN_815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_817 = 8'h75 == r_count_2_io_out ? io_r_117_b : _GEN_816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_818 = 8'h76 == r_count_2_io_out ? io_r_118_b : _GEN_817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_819 = 8'h77 == r_count_2_io_out ? io_r_119_b : _GEN_818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_820 = 8'h78 == r_count_2_io_out ? io_r_120_b : _GEN_819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_821 = 8'h79 == r_count_2_io_out ? io_r_121_b : _GEN_820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_822 = 8'h7a == r_count_2_io_out ? io_r_122_b : _GEN_821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_823 = 8'h7b == r_count_2_io_out ? io_r_123_b : _GEN_822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_824 = 8'h7c == r_count_2_io_out ? io_r_124_b : _GEN_823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_825 = 8'h7d == r_count_2_io_out ? io_r_125_b : _GEN_824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_826 = 8'h7e == r_count_2_io_out ? io_r_126_b : _GEN_825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_827 = 8'h7f == r_count_2_io_out ? io_r_127_b : _GEN_826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_828 = 8'h80 == r_count_2_io_out ? io_r_128_b : _GEN_827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_829 = 8'h81 == r_count_2_io_out ? io_r_129_b : _GEN_828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_830 = 8'h82 == r_count_2_io_out ? io_r_130_b : _GEN_829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_831 = 8'h83 == r_count_2_io_out ? io_r_131_b : _GEN_830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_832 = 8'h84 == r_count_2_io_out ? io_r_132_b : _GEN_831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_833 = 8'h85 == r_count_2_io_out ? io_r_133_b : _GEN_832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_834 = 8'h86 == r_count_2_io_out ? io_r_134_b : _GEN_833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_835 = 8'h87 == r_count_2_io_out ? io_r_135_b : _GEN_834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_836 = 8'h88 == r_count_2_io_out ? io_r_136_b : _GEN_835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_837 = 8'h89 == r_count_2_io_out ? io_r_137_b : _GEN_836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_838 = 8'h8a == r_count_2_io_out ? io_r_138_b : _GEN_837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_839 = 8'h8b == r_count_2_io_out ? io_r_139_b : _GEN_838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_840 = 8'h8c == r_count_2_io_out ? io_r_140_b : _GEN_839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_841 = 8'h8d == r_count_2_io_out ? io_r_141_b : _GEN_840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_842 = 8'h8e == r_count_2_io_out ? io_r_142_b : _GEN_841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_843 = 8'h8f == r_count_2_io_out ? io_r_143_b : _GEN_842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_844 = 8'h90 == r_count_2_io_out ? io_r_144_b : _GEN_843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_845 = 8'h91 == r_count_2_io_out ? io_r_145_b : _GEN_844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_846 = 8'h92 == r_count_2_io_out ? io_r_146_b : _GEN_845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_847 = 8'h93 == r_count_2_io_out ? io_r_147_b : _GEN_846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_848 = 8'h94 == r_count_2_io_out ? io_r_148_b : _GEN_847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_849 = 8'h95 == r_count_2_io_out ? io_r_149_b : _GEN_848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_850 = 8'h96 == r_count_2_io_out ? io_r_150_b : _GEN_849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_851 = 8'h97 == r_count_2_io_out ? io_r_151_b : _GEN_850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_852 = 8'h98 == r_count_2_io_out ? io_r_152_b : _GEN_851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_853 = 8'h99 == r_count_2_io_out ? io_r_153_b : _GEN_852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_854 = 8'h9a == r_count_2_io_out ? io_r_154_b : _GEN_853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_855 = 8'h9b == r_count_2_io_out ? io_r_155_b : _GEN_854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_856 = 8'h9c == r_count_2_io_out ? io_r_156_b : _GEN_855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_857 = 8'h9d == r_count_2_io_out ? io_r_157_b : _GEN_856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_858 = 8'h9e == r_count_2_io_out ? io_r_158_b : _GEN_857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_859 = 8'h9f == r_count_2_io_out ? io_r_159_b : _GEN_858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_860 = 8'ha0 == r_count_2_io_out ? io_r_160_b : _GEN_859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_861 = 8'ha1 == r_count_2_io_out ? io_r_161_b : _GEN_860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_862 = 8'ha2 == r_count_2_io_out ? io_r_162_b : _GEN_861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_863 = 8'ha3 == r_count_2_io_out ? io_r_163_b : _GEN_862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_864 = 8'ha4 == r_count_2_io_out ? io_r_164_b : _GEN_863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_865 = 8'ha5 == r_count_2_io_out ? io_r_165_b : _GEN_864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_866 = 8'ha6 == r_count_2_io_out ? io_r_166_b : _GEN_865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_867 = 8'ha7 == r_count_2_io_out ? io_r_167_b : _GEN_866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_868 = 8'ha8 == r_count_2_io_out ? io_r_168_b : _GEN_867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_869 = 8'ha9 == r_count_2_io_out ? io_r_169_b : _GEN_868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_870 = 8'haa == r_count_2_io_out ? io_r_170_b : _GEN_869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_871 = 8'hab == r_count_2_io_out ? io_r_171_b : _GEN_870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_872 = 8'hac == r_count_2_io_out ? io_r_172_b : _GEN_871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_873 = 8'had == r_count_2_io_out ? io_r_173_b : _GEN_872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_874 = 8'hae == r_count_2_io_out ? io_r_174_b : _GEN_873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_875 = 8'haf == r_count_2_io_out ? io_r_175_b : _GEN_874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_876 = 8'hb0 == r_count_2_io_out ? io_r_176_b : _GEN_875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_877 = 8'hb1 == r_count_2_io_out ? io_r_177_b : _GEN_876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_878 = 8'hb2 == r_count_2_io_out ? io_r_178_b : _GEN_877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_879 = 8'hb3 == r_count_2_io_out ? io_r_179_b : _GEN_878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_880 = 8'hb4 == r_count_2_io_out ? io_r_180_b : _GEN_879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_881 = 8'hb5 == r_count_2_io_out ? io_r_181_b : _GEN_880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_882 = 8'hb6 == r_count_2_io_out ? io_r_182_b : _GEN_881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_883 = 8'hb7 == r_count_2_io_out ? io_r_183_b : _GEN_882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_884 = 8'hb8 == r_count_2_io_out ? io_r_184_b : _GEN_883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_885 = 8'hb9 == r_count_2_io_out ? io_r_185_b : _GEN_884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_886 = 8'hba == r_count_2_io_out ? io_r_186_b : _GEN_885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_887 = 8'hbb == r_count_2_io_out ? io_r_187_b : _GEN_886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_888 = 8'hbc == r_count_2_io_out ? io_r_188_b : _GEN_887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_889 = 8'hbd == r_count_2_io_out ? io_r_189_b : _GEN_888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_890 = 8'hbe == r_count_2_io_out ? io_r_190_b : _GEN_889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_891 = 8'hbf == r_count_2_io_out ? io_r_191_b : _GEN_890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_892 = 8'hc0 == r_count_2_io_out ? io_r_192_b : _GEN_891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_893 = 8'hc1 == r_count_2_io_out ? io_r_193_b : _GEN_892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_894 = 8'hc2 == r_count_2_io_out ? io_r_194_b : _GEN_893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_895 = 8'hc3 == r_count_2_io_out ? io_r_195_b : _GEN_894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_896 = 8'hc4 == r_count_2_io_out ? io_r_196_b : _GEN_895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_897 = 8'hc5 == r_count_2_io_out ? io_r_197_b : _GEN_896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_898 = 8'hc6 == r_count_2_io_out ? io_r_198_b : _GEN_897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_901 = 8'h1 == r_count_3_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_902 = 8'h2 == r_count_3_io_out ? io_r_2_b : _GEN_901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_903 = 8'h3 == r_count_3_io_out ? io_r_3_b : _GEN_902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_904 = 8'h4 == r_count_3_io_out ? io_r_4_b : _GEN_903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_905 = 8'h5 == r_count_3_io_out ? io_r_5_b : _GEN_904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_906 = 8'h6 == r_count_3_io_out ? io_r_6_b : _GEN_905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_907 = 8'h7 == r_count_3_io_out ? io_r_7_b : _GEN_906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_908 = 8'h8 == r_count_3_io_out ? io_r_8_b : _GEN_907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_909 = 8'h9 == r_count_3_io_out ? io_r_9_b : _GEN_908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_910 = 8'ha == r_count_3_io_out ? io_r_10_b : _GEN_909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_911 = 8'hb == r_count_3_io_out ? io_r_11_b : _GEN_910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_912 = 8'hc == r_count_3_io_out ? io_r_12_b : _GEN_911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_913 = 8'hd == r_count_3_io_out ? io_r_13_b : _GEN_912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_914 = 8'he == r_count_3_io_out ? io_r_14_b : _GEN_913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_915 = 8'hf == r_count_3_io_out ? io_r_15_b : _GEN_914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_916 = 8'h10 == r_count_3_io_out ? io_r_16_b : _GEN_915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_917 = 8'h11 == r_count_3_io_out ? io_r_17_b : _GEN_916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_918 = 8'h12 == r_count_3_io_out ? io_r_18_b : _GEN_917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_919 = 8'h13 == r_count_3_io_out ? io_r_19_b : _GEN_918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_920 = 8'h14 == r_count_3_io_out ? io_r_20_b : _GEN_919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_921 = 8'h15 == r_count_3_io_out ? io_r_21_b : _GEN_920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_922 = 8'h16 == r_count_3_io_out ? io_r_22_b : _GEN_921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_923 = 8'h17 == r_count_3_io_out ? io_r_23_b : _GEN_922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_924 = 8'h18 == r_count_3_io_out ? io_r_24_b : _GEN_923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_925 = 8'h19 == r_count_3_io_out ? io_r_25_b : _GEN_924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_926 = 8'h1a == r_count_3_io_out ? io_r_26_b : _GEN_925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_927 = 8'h1b == r_count_3_io_out ? io_r_27_b : _GEN_926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_928 = 8'h1c == r_count_3_io_out ? io_r_28_b : _GEN_927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_929 = 8'h1d == r_count_3_io_out ? io_r_29_b : _GEN_928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_930 = 8'h1e == r_count_3_io_out ? io_r_30_b : _GEN_929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_931 = 8'h1f == r_count_3_io_out ? io_r_31_b : _GEN_930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_932 = 8'h20 == r_count_3_io_out ? io_r_32_b : _GEN_931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_933 = 8'h21 == r_count_3_io_out ? io_r_33_b : _GEN_932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_934 = 8'h22 == r_count_3_io_out ? io_r_34_b : _GEN_933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_935 = 8'h23 == r_count_3_io_out ? io_r_35_b : _GEN_934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_936 = 8'h24 == r_count_3_io_out ? io_r_36_b : _GEN_935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_937 = 8'h25 == r_count_3_io_out ? io_r_37_b : _GEN_936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_938 = 8'h26 == r_count_3_io_out ? io_r_38_b : _GEN_937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_939 = 8'h27 == r_count_3_io_out ? io_r_39_b : _GEN_938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_940 = 8'h28 == r_count_3_io_out ? io_r_40_b : _GEN_939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_941 = 8'h29 == r_count_3_io_out ? io_r_41_b : _GEN_940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_942 = 8'h2a == r_count_3_io_out ? io_r_42_b : _GEN_941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_943 = 8'h2b == r_count_3_io_out ? io_r_43_b : _GEN_942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_944 = 8'h2c == r_count_3_io_out ? io_r_44_b : _GEN_943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_945 = 8'h2d == r_count_3_io_out ? io_r_45_b : _GEN_944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_946 = 8'h2e == r_count_3_io_out ? io_r_46_b : _GEN_945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_947 = 8'h2f == r_count_3_io_out ? io_r_47_b : _GEN_946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_948 = 8'h30 == r_count_3_io_out ? io_r_48_b : _GEN_947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_949 = 8'h31 == r_count_3_io_out ? io_r_49_b : _GEN_948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_950 = 8'h32 == r_count_3_io_out ? io_r_50_b : _GEN_949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_951 = 8'h33 == r_count_3_io_out ? io_r_51_b : _GEN_950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_952 = 8'h34 == r_count_3_io_out ? io_r_52_b : _GEN_951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_953 = 8'h35 == r_count_3_io_out ? io_r_53_b : _GEN_952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_954 = 8'h36 == r_count_3_io_out ? io_r_54_b : _GEN_953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_955 = 8'h37 == r_count_3_io_out ? io_r_55_b : _GEN_954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_956 = 8'h38 == r_count_3_io_out ? io_r_56_b : _GEN_955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_957 = 8'h39 == r_count_3_io_out ? io_r_57_b : _GEN_956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_958 = 8'h3a == r_count_3_io_out ? io_r_58_b : _GEN_957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_959 = 8'h3b == r_count_3_io_out ? io_r_59_b : _GEN_958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_960 = 8'h3c == r_count_3_io_out ? io_r_60_b : _GEN_959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_961 = 8'h3d == r_count_3_io_out ? io_r_61_b : _GEN_960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_962 = 8'h3e == r_count_3_io_out ? io_r_62_b : _GEN_961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_963 = 8'h3f == r_count_3_io_out ? io_r_63_b : _GEN_962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_964 = 8'h40 == r_count_3_io_out ? io_r_64_b : _GEN_963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_965 = 8'h41 == r_count_3_io_out ? io_r_65_b : _GEN_964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_966 = 8'h42 == r_count_3_io_out ? io_r_66_b : _GEN_965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_967 = 8'h43 == r_count_3_io_out ? io_r_67_b : _GEN_966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_968 = 8'h44 == r_count_3_io_out ? io_r_68_b : _GEN_967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_969 = 8'h45 == r_count_3_io_out ? io_r_69_b : _GEN_968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_970 = 8'h46 == r_count_3_io_out ? io_r_70_b : _GEN_969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_971 = 8'h47 == r_count_3_io_out ? io_r_71_b : _GEN_970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_972 = 8'h48 == r_count_3_io_out ? io_r_72_b : _GEN_971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_973 = 8'h49 == r_count_3_io_out ? io_r_73_b : _GEN_972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_974 = 8'h4a == r_count_3_io_out ? io_r_74_b : _GEN_973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_975 = 8'h4b == r_count_3_io_out ? io_r_75_b : _GEN_974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_976 = 8'h4c == r_count_3_io_out ? io_r_76_b : _GEN_975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_977 = 8'h4d == r_count_3_io_out ? io_r_77_b : _GEN_976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_978 = 8'h4e == r_count_3_io_out ? io_r_78_b : _GEN_977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_979 = 8'h4f == r_count_3_io_out ? io_r_79_b : _GEN_978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_980 = 8'h50 == r_count_3_io_out ? io_r_80_b : _GEN_979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_981 = 8'h51 == r_count_3_io_out ? io_r_81_b : _GEN_980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_982 = 8'h52 == r_count_3_io_out ? io_r_82_b : _GEN_981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_983 = 8'h53 == r_count_3_io_out ? io_r_83_b : _GEN_982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_984 = 8'h54 == r_count_3_io_out ? io_r_84_b : _GEN_983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_985 = 8'h55 == r_count_3_io_out ? io_r_85_b : _GEN_984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_986 = 8'h56 == r_count_3_io_out ? io_r_86_b : _GEN_985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_987 = 8'h57 == r_count_3_io_out ? io_r_87_b : _GEN_986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_988 = 8'h58 == r_count_3_io_out ? io_r_88_b : _GEN_987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_989 = 8'h59 == r_count_3_io_out ? io_r_89_b : _GEN_988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_990 = 8'h5a == r_count_3_io_out ? io_r_90_b : _GEN_989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_991 = 8'h5b == r_count_3_io_out ? io_r_91_b : _GEN_990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_992 = 8'h5c == r_count_3_io_out ? io_r_92_b : _GEN_991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_993 = 8'h5d == r_count_3_io_out ? io_r_93_b : _GEN_992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_994 = 8'h5e == r_count_3_io_out ? io_r_94_b : _GEN_993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_995 = 8'h5f == r_count_3_io_out ? io_r_95_b : _GEN_994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_996 = 8'h60 == r_count_3_io_out ? io_r_96_b : _GEN_995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_997 = 8'h61 == r_count_3_io_out ? io_r_97_b : _GEN_996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_998 = 8'h62 == r_count_3_io_out ? io_r_98_b : _GEN_997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_999 = 8'h63 == r_count_3_io_out ? io_r_99_b : _GEN_998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1000 = 8'h64 == r_count_3_io_out ? io_r_100_b : _GEN_999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1001 = 8'h65 == r_count_3_io_out ? io_r_101_b : _GEN_1000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1002 = 8'h66 == r_count_3_io_out ? io_r_102_b : _GEN_1001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1003 = 8'h67 == r_count_3_io_out ? io_r_103_b : _GEN_1002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1004 = 8'h68 == r_count_3_io_out ? io_r_104_b : _GEN_1003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1005 = 8'h69 == r_count_3_io_out ? io_r_105_b : _GEN_1004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1006 = 8'h6a == r_count_3_io_out ? io_r_106_b : _GEN_1005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1007 = 8'h6b == r_count_3_io_out ? io_r_107_b : _GEN_1006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1008 = 8'h6c == r_count_3_io_out ? io_r_108_b : _GEN_1007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1009 = 8'h6d == r_count_3_io_out ? io_r_109_b : _GEN_1008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1010 = 8'h6e == r_count_3_io_out ? io_r_110_b : _GEN_1009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1011 = 8'h6f == r_count_3_io_out ? io_r_111_b : _GEN_1010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1012 = 8'h70 == r_count_3_io_out ? io_r_112_b : _GEN_1011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1013 = 8'h71 == r_count_3_io_out ? io_r_113_b : _GEN_1012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1014 = 8'h72 == r_count_3_io_out ? io_r_114_b : _GEN_1013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1015 = 8'h73 == r_count_3_io_out ? io_r_115_b : _GEN_1014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1016 = 8'h74 == r_count_3_io_out ? io_r_116_b : _GEN_1015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1017 = 8'h75 == r_count_3_io_out ? io_r_117_b : _GEN_1016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1018 = 8'h76 == r_count_3_io_out ? io_r_118_b : _GEN_1017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1019 = 8'h77 == r_count_3_io_out ? io_r_119_b : _GEN_1018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1020 = 8'h78 == r_count_3_io_out ? io_r_120_b : _GEN_1019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1021 = 8'h79 == r_count_3_io_out ? io_r_121_b : _GEN_1020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1022 = 8'h7a == r_count_3_io_out ? io_r_122_b : _GEN_1021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1023 = 8'h7b == r_count_3_io_out ? io_r_123_b : _GEN_1022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1024 = 8'h7c == r_count_3_io_out ? io_r_124_b : _GEN_1023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1025 = 8'h7d == r_count_3_io_out ? io_r_125_b : _GEN_1024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1026 = 8'h7e == r_count_3_io_out ? io_r_126_b : _GEN_1025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1027 = 8'h7f == r_count_3_io_out ? io_r_127_b : _GEN_1026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1028 = 8'h80 == r_count_3_io_out ? io_r_128_b : _GEN_1027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1029 = 8'h81 == r_count_3_io_out ? io_r_129_b : _GEN_1028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1030 = 8'h82 == r_count_3_io_out ? io_r_130_b : _GEN_1029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1031 = 8'h83 == r_count_3_io_out ? io_r_131_b : _GEN_1030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1032 = 8'h84 == r_count_3_io_out ? io_r_132_b : _GEN_1031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1033 = 8'h85 == r_count_3_io_out ? io_r_133_b : _GEN_1032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1034 = 8'h86 == r_count_3_io_out ? io_r_134_b : _GEN_1033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1035 = 8'h87 == r_count_3_io_out ? io_r_135_b : _GEN_1034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1036 = 8'h88 == r_count_3_io_out ? io_r_136_b : _GEN_1035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1037 = 8'h89 == r_count_3_io_out ? io_r_137_b : _GEN_1036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1038 = 8'h8a == r_count_3_io_out ? io_r_138_b : _GEN_1037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1039 = 8'h8b == r_count_3_io_out ? io_r_139_b : _GEN_1038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1040 = 8'h8c == r_count_3_io_out ? io_r_140_b : _GEN_1039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1041 = 8'h8d == r_count_3_io_out ? io_r_141_b : _GEN_1040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1042 = 8'h8e == r_count_3_io_out ? io_r_142_b : _GEN_1041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1043 = 8'h8f == r_count_3_io_out ? io_r_143_b : _GEN_1042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1044 = 8'h90 == r_count_3_io_out ? io_r_144_b : _GEN_1043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1045 = 8'h91 == r_count_3_io_out ? io_r_145_b : _GEN_1044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1046 = 8'h92 == r_count_3_io_out ? io_r_146_b : _GEN_1045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1047 = 8'h93 == r_count_3_io_out ? io_r_147_b : _GEN_1046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1048 = 8'h94 == r_count_3_io_out ? io_r_148_b : _GEN_1047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1049 = 8'h95 == r_count_3_io_out ? io_r_149_b : _GEN_1048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1050 = 8'h96 == r_count_3_io_out ? io_r_150_b : _GEN_1049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1051 = 8'h97 == r_count_3_io_out ? io_r_151_b : _GEN_1050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1052 = 8'h98 == r_count_3_io_out ? io_r_152_b : _GEN_1051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1053 = 8'h99 == r_count_3_io_out ? io_r_153_b : _GEN_1052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1054 = 8'h9a == r_count_3_io_out ? io_r_154_b : _GEN_1053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1055 = 8'h9b == r_count_3_io_out ? io_r_155_b : _GEN_1054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1056 = 8'h9c == r_count_3_io_out ? io_r_156_b : _GEN_1055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1057 = 8'h9d == r_count_3_io_out ? io_r_157_b : _GEN_1056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1058 = 8'h9e == r_count_3_io_out ? io_r_158_b : _GEN_1057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1059 = 8'h9f == r_count_3_io_out ? io_r_159_b : _GEN_1058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1060 = 8'ha0 == r_count_3_io_out ? io_r_160_b : _GEN_1059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1061 = 8'ha1 == r_count_3_io_out ? io_r_161_b : _GEN_1060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1062 = 8'ha2 == r_count_3_io_out ? io_r_162_b : _GEN_1061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1063 = 8'ha3 == r_count_3_io_out ? io_r_163_b : _GEN_1062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1064 = 8'ha4 == r_count_3_io_out ? io_r_164_b : _GEN_1063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1065 = 8'ha5 == r_count_3_io_out ? io_r_165_b : _GEN_1064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1066 = 8'ha6 == r_count_3_io_out ? io_r_166_b : _GEN_1065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1067 = 8'ha7 == r_count_3_io_out ? io_r_167_b : _GEN_1066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1068 = 8'ha8 == r_count_3_io_out ? io_r_168_b : _GEN_1067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1069 = 8'ha9 == r_count_3_io_out ? io_r_169_b : _GEN_1068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1070 = 8'haa == r_count_3_io_out ? io_r_170_b : _GEN_1069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1071 = 8'hab == r_count_3_io_out ? io_r_171_b : _GEN_1070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1072 = 8'hac == r_count_3_io_out ? io_r_172_b : _GEN_1071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1073 = 8'had == r_count_3_io_out ? io_r_173_b : _GEN_1072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1074 = 8'hae == r_count_3_io_out ? io_r_174_b : _GEN_1073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1075 = 8'haf == r_count_3_io_out ? io_r_175_b : _GEN_1074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1076 = 8'hb0 == r_count_3_io_out ? io_r_176_b : _GEN_1075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1077 = 8'hb1 == r_count_3_io_out ? io_r_177_b : _GEN_1076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1078 = 8'hb2 == r_count_3_io_out ? io_r_178_b : _GEN_1077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1079 = 8'hb3 == r_count_3_io_out ? io_r_179_b : _GEN_1078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1080 = 8'hb4 == r_count_3_io_out ? io_r_180_b : _GEN_1079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1081 = 8'hb5 == r_count_3_io_out ? io_r_181_b : _GEN_1080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1082 = 8'hb6 == r_count_3_io_out ? io_r_182_b : _GEN_1081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1083 = 8'hb7 == r_count_3_io_out ? io_r_183_b : _GEN_1082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1084 = 8'hb8 == r_count_3_io_out ? io_r_184_b : _GEN_1083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1085 = 8'hb9 == r_count_3_io_out ? io_r_185_b : _GEN_1084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1086 = 8'hba == r_count_3_io_out ? io_r_186_b : _GEN_1085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1087 = 8'hbb == r_count_3_io_out ? io_r_187_b : _GEN_1086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1088 = 8'hbc == r_count_3_io_out ? io_r_188_b : _GEN_1087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1089 = 8'hbd == r_count_3_io_out ? io_r_189_b : _GEN_1088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1090 = 8'hbe == r_count_3_io_out ? io_r_190_b : _GEN_1089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1091 = 8'hbf == r_count_3_io_out ? io_r_191_b : _GEN_1090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1092 = 8'hc0 == r_count_3_io_out ? io_r_192_b : _GEN_1091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1093 = 8'hc1 == r_count_3_io_out ? io_r_193_b : _GEN_1092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1094 = 8'hc2 == r_count_3_io_out ? io_r_194_b : _GEN_1093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1095 = 8'hc3 == r_count_3_io_out ? io_r_195_b : _GEN_1094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1096 = 8'hc4 == r_count_3_io_out ? io_r_196_b : _GEN_1095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1097 = 8'hc5 == r_count_3_io_out ? io_r_197_b : _GEN_1096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1098 = 8'hc6 == r_count_3_io_out ? io_r_198_b : _GEN_1097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1101 = 8'h1 == r_count_4_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1102 = 8'h2 == r_count_4_io_out ? io_r_2_b : _GEN_1101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1103 = 8'h3 == r_count_4_io_out ? io_r_3_b : _GEN_1102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1104 = 8'h4 == r_count_4_io_out ? io_r_4_b : _GEN_1103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1105 = 8'h5 == r_count_4_io_out ? io_r_5_b : _GEN_1104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1106 = 8'h6 == r_count_4_io_out ? io_r_6_b : _GEN_1105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1107 = 8'h7 == r_count_4_io_out ? io_r_7_b : _GEN_1106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1108 = 8'h8 == r_count_4_io_out ? io_r_8_b : _GEN_1107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1109 = 8'h9 == r_count_4_io_out ? io_r_9_b : _GEN_1108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1110 = 8'ha == r_count_4_io_out ? io_r_10_b : _GEN_1109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1111 = 8'hb == r_count_4_io_out ? io_r_11_b : _GEN_1110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1112 = 8'hc == r_count_4_io_out ? io_r_12_b : _GEN_1111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1113 = 8'hd == r_count_4_io_out ? io_r_13_b : _GEN_1112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1114 = 8'he == r_count_4_io_out ? io_r_14_b : _GEN_1113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1115 = 8'hf == r_count_4_io_out ? io_r_15_b : _GEN_1114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1116 = 8'h10 == r_count_4_io_out ? io_r_16_b : _GEN_1115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1117 = 8'h11 == r_count_4_io_out ? io_r_17_b : _GEN_1116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1118 = 8'h12 == r_count_4_io_out ? io_r_18_b : _GEN_1117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1119 = 8'h13 == r_count_4_io_out ? io_r_19_b : _GEN_1118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1120 = 8'h14 == r_count_4_io_out ? io_r_20_b : _GEN_1119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1121 = 8'h15 == r_count_4_io_out ? io_r_21_b : _GEN_1120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1122 = 8'h16 == r_count_4_io_out ? io_r_22_b : _GEN_1121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1123 = 8'h17 == r_count_4_io_out ? io_r_23_b : _GEN_1122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1124 = 8'h18 == r_count_4_io_out ? io_r_24_b : _GEN_1123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1125 = 8'h19 == r_count_4_io_out ? io_r_25_b : _GEN_1124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1126 = 8'h1a == r_count_4_io_out ? io_r_26_b : _GEN_1125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1127 = 8'h1b == r_count_4_io_out ? io_r_27_b : _GEN_1126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1128 = 8'h1c == r_count_4_io_out ? io_r_28_b : _GEN_1127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1129 = 8'h1d == r_count_4_io_out ? io_r_29_b : _GEN_1128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1130 = 8'h1e == r_count_4_io_out ? io_r_30_b : _GEN_1129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1131 = 8'h1f == r_count_4_io_out ? io_r_31_b : _GEN_1130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1132 = 8'h20 == r_count_4_io_out ? io_r_32_b : _GEN_1131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1133 = 8'h21 == r_count_4_io_out ? io_r_33_b : _GEN_1132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1134 = 8'h22 == r_count_4_io_out ? io_r_34_b : _GEN_1133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1135 = 8'h23 == r_count_4_io_out ? io_r_35_b : _GEN_1134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1136 = 8'h24 == r_count_4_io_out ? io_r_36_b : _GEN_1135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1137 = 8'h25 == r_count_4_io_out ? io_r_37_b : _GEN_1136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1138 = 8'h26 == r_count_4_io_out ? io_r_38_b : _GEN_1137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1139 = 8'h27 == r_count_4_io_out ? io_r_39_b : _GEN_1138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1140 = 8'h28 == r_count_4_io_out ? io_r_40_b : _GEN_1139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1141 = 8'h29 == r_count_4_io_out ? io_r_41_b : _GEN_1140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1142 = 8'h2a == r_count_4_io_out ? io_r_42_b : _GEN_1141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1143 = 8'h2b == r_count_4_io_out ? io_r_43_b : _GEN_1142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1144 = 8'h2c == r_count_4_io_out ? io_r_44_b : _GEN_1143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1145 = 8'h2d == r_count_4_io_out ? io_r_45_b : _GEN_1144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1146 = 8'h2e == r_count_4_io_out ? io_r_46_b : _GEN_1145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1147 = 8'h2f == r_count_4_io_out ? io_r_47_b : _GEN_1146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1148 = 8'h30 == r_count_4_io_out ? io_r_48_b : _GEN_1147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1149 = 8'h31 == r_count_4_io_out ? io_r_49_b : _GEN_1148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1150 = 8'h32 == r_count_4_io_out ? io_r_50_b : _GEN_1149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1151 = 8'h33 == r_count_4_io_out ? io_r_51_b : _GEN_1150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1152 = 8'h34 == r_count_4_io_out ? io_r_52_b : _GEN_1151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1153 = 8'h35 == r_count_4_io_out ? io_r_53_b : _GEN_1152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1154 = 8'h36 == r_count_4_io_out ? io_r_54_b : _GEN_1153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1155 = 8'h37 == r_count_4_io_out ? io_r_55_b : _GEN_1154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1156 = 8'h38 == r_count_4_io_out ? io_r_56_b : _GEN_1155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1157 = 8'h39 == r_count_4_io_out ? io_r_57_b : _GEN_1156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1158 = 8'h3a == r_count_4_io_out ? io_r_58_b : _GEN_1157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1159 = 8'h3b == r_count_4_io_out ? io_r_59_b : _GEN_1158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1160 = 8'h3c == r_count_4_io_out ? io_r_60_b : _GEN_1159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1161 = 8'h3d == r_count_4_io_out ? io_r_61_b : _GEN_1160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1162 = 8'h3e == r_count_4_io_out ? io_r_62_b : _GEN_1161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1163 = 8'h3f == r_count_4_io_out ? io_r_63_b : _GEN_1162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1164 = 8'h40 == r_count_4_io_out ? io_r_64_b : _GEN_1163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1165 = 8'h41 == r_count_4_io_out ? io_r_65_b : _GEN_1164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1166 = 8'h42 == r_count_4_io_out ? io_r_66_b : _GEN_1165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1167 = 8'h43 == r_count_4_io_out ? io_r_67_b : _GEN_1166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1168 = 8'h44 == r_count_4_io_out ? io_r_68_b : _GEN_1167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1169 = 8'h45 == r_count_4_io_out ? io_r_69_b : _GEN_1168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1170 = 8'h46 == r_count_4_io_out ? io_r_70_b : _GEN_1169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1171 = 8'h47 == r_count_4_io_out ? io_r_71_b : _GEN_1170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1172 = 8'h48 == r_count_4_io_out ? io_r_72_b : _GEN_1171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1173 = 8'h49 == r_count_4_io_out ? io_r_73_b : _GEN_1172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1174 = 8'h4a == r_count_4_io_out ? io_r_74_b : _GEN_1173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1175 = 8'h4b == r_count_4_io_out ? io_r_75_b : _GEN_1174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1176 = 8'h4c == r_count_4_io_out ? io_r_76_b : _GEN_1175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1177 = 8'h4d == r_count_4_io_out ? io_r_77_b : _GEN_1176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1178 = 8'h4e == r_count_4_io_out ? io_r_78_b : _GEN_1177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1179 = 8'h4f == r_count_4_io_out ? io_r_79_b : _GEN_1178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1180 = 8'h50 == r_count_4_io_out ? io_r_80_b : _GEN_1179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1181 = 8'h51 == r_count_4_io_out ? io_r_81_b : _GEN_1180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1182 = 8'h52 == r_count_4_io_out ? io_r_82_b : _GEN_1181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1183 = 8'h53 == r_count_4_io_out ? io_r_83_b : _GEN_1182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1184 = 8'h54 == r_count_4_io_out ? io_r_84_b : _GEN_1183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1185 = 8'h55 == r_count_4_io_out ? io_r_85_b : _GEN_1184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1186 = 8'h56 == r_count_4_io_out ? io_r_86_b : _GEN_1185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1187 = 8'h57 == r_count_4_io_out ? io_r_87_b : _GEN_1186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1188 = 8'h58 == r_count_4_io_out ? io_r_88_b : _GEN_1187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1189 = 8'h59 == r_count_4_io_out ? io_r_89_b : _GEN_1188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1190 = 8'h5a == r_count_4_io_out ? io_r_90_b : _GEN_1189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1191 = 8'h5b == r_count_4_io_out ? io_r_91_b : _GEN_1190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1192 = 8'h5c == r_count_4_io_out ? io_r_92_b : _GEN_1191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1193 = 8'h5d == r_count_4_io_out ? io_r_93_b : _GEN_1192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1194 = 8'h5e == r_count_4_io_out ? io_r_94_b : _GEN_1193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1195 = 8'h5f == r_count_4_io_out ? io_r_95_b : _GEN_1194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1196 = 8'h60 == r_count_4_io_out ? io_r_96_b : _GEN_1195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1197 = 8'h61 == r_count_4_io_out ? io_r_97_b : _GEN_1196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1198 = 8'h62 == r_count_4_io_out ? io_r_98_b : _GEN_1197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1199 = 8'h63 == r_count_4_io_out ? io_r_99_b : _GEN_1198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1200 = 8'h64 == r_count_4_io_out ? io_r_100_b : _GEN_1199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1201 = 8'h65 == r_count_4_io_out ? io_r_101_b : _GEN_1200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1202 = 8'h66 == r_count_4_io_out ? io_r_102_b : _GEN_1201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1203 = 8'h67 == r_count_4_io_out ? io_r_103_b : _GEN_1202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1204 = 8'h68 == r_count_4_io_out ? io_r_104_b : _GEN_1203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1205 = 8'h69 == r_count_4_io_out ? io_r_105_b : _GEN_1204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1206 = 8'h6a == r_count_4_io_out ? io_r_106_b : _GEN_1205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1207 = 8'h6b == r_count_4_io_out ? io_r_107_b : _GEN_1206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1208 = 8'h6c == r_count_4_io_out ? io_r_108_b : _GEN_1207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1209 = 8'h6d == r_count_4_io_out ? io_r_109_b : _GEN_1208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1210 = 8'h6e == r_count_4_io_out ? io_r_110_b : _GEN_1209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1211 = 8'h6f == r_count_4_io_out ? io_r_111_b : _GEN_1210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1212 = 8'h70 == r_count_4_io_out ? io_r_112_b : _GEN_1211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1213 = 8'h71 == r_count_4_io_out ? io_r_113_b : _GEN_1212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1214 = 8'h72 == r_count_4_io_out ? io_r_114_b : _GEN_1213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1215 = 8'h73 == r_count_4_io_out ? io_r_115_b : _GEN_1214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1216 = 8'h74 == r_count_4_io_out ? io_r_116_b : _GEN_1215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1217 = 8'h75 == r_count_4_io_out ? io_r_117_b : _GEN_1216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1218 = 8'h76 == r_count_4_io_out ? io_r_118_b : _GEN_1217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1219 = 8'h77 == r_count_4_io_out ? io_r_119_b : _GEN_1218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1220 = 8'h78 == r_count_4_io_out ? io_r_120_b : _GEN_1219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1221 = 8'h79 == r_count_4_io_out ? io_r_121_b : _GEN_1220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1222 = 8'h7a == r_count_4_io_out ? io_r_122_b : _GEN_1221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1223 = 8'h7b == r_count_4_io_out ? io_r_123_b : _GEN_1222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1224 = 8'h7c == r_count_4_io_out ? io_r_124_b : _GEN_1223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1225 = 8'h7d == r_count_4_io_out ? io_r_125_b : _GEN_1224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1226 = 8'h7e == r_count_4_io_out ? io_r_126_b : _GEN_1225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1227 = 8'h7f == r_count_4_io_out ? io_r_127_b : _GEN_1226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1228 = 8'h80 == r_count_4_io_out ? io_r_128_b : _GEN_1227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1229 = 8'h81 == r_count_4_io_out ? io_r_129_b : _GEN_1228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1230 = 8'h82 == r_count_4_io_out ? io_r_130_b : _GEN_1229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1231 = 8'h83 == r_count_4_io_out ? io_r_131_b : _GEN_1230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1232 = 8'h84 == r_count_4_io_out ? io_r_132_b : _GEN_1231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1233 = 8'h85 == r_count_4_io_out ? io_r_133_b : _GEN_1232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1234 = 8'h86 == r_count_4_io_out ? io_r_134_b : _GEN_1233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1235 = 8'h87 == r_count_4_io_out ? io_r_135_b : _GEN_1234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1236 = 8'h88 == r_count_4_io_out ? io_r_136_b : _GEN_1235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1237 = 8'h89 == r_count_4_io_out ? io_r_137_b : _GEN_1236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1238 = 8'h8a == r_count_4_io_out ? io_r_138_b : _GEN_1237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1239 = 8'h8b == r_count_4_io_out ? io_r_139_b : _GEN_1238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1240 = 8'h8c == r_count_4_io_out ? io_r_140_b : _GEN_1239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1241 = 8'h8d == r_count_4_io_out ? io_r_141_b : _GEN_1240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1242 = 8'h8e == r_count_4_io_out ? io_r_142_b : _GEN_1241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1243 = 8'h8f == r_count_4_io_out ? io_r_143_b : _GEN_1242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1244 = 8'h90 == r_count_4_io_out ? io_r_144_b : _GEN_1243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1245 = 8'h91 == r_count_4_io_out ? io_r_145_b : _GEN_1244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1246 = 8'h92 == r_count_4_io_out ? io_r_146_b : _GEN_1245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1247 = 8'h93 == r_count_4_io_out ? io_r_147_b : _GEN_1246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1248 = 8'h94 == r_count_4_io_out ? io_r_148_b : _GEN_1247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1249 = 8'h95 == r_count_4_io_out ? io_r_149_b : _GEN_1248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1250 = 8'h96 == r_count_4_io_out ? io_r_150_b : _GEN_1249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1251 = 8'h97 == r_count_4_io_out ? io_r_151_b : _GEN_1250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1252 = 8'h98 == r_count_4_io_out ? io_r_152_b : _GEN_1251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1253 = 8'h99 == r_count_4_io_out ? io_r_153_b : _GEN_1252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1254 = 8'h9a == r_count_4_io_out ? io_r_154_b : _GEN_1253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1255 = 8'h9b == r_count_4_io_out ? io_r_155_b : _GEN_1254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1256 = 8'h9c == r_count_4_io_out ? io_r_156_b : _GEN_1255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1257 = 8'h9d == r_count_4_io_out ? io_r_157_b : _GEN_1256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1258 = 8'h9e == r_count_4_io_out ? io_r_158_b : _GEN_1257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1259 = 8'h9f == r_count_4_io_out ? io_r_159_b : _GEN_1258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1260 = 8'ha0 == r_count_4_io_out ? io_r_160_b : _GEN_1259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1261 = 8'ha1 == r_count_4_io_out ? io_r_161_b : _GEN_1260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1262 = 8'ha2 == r_count_4_io_out ? io_r_162_b : _GEN_1261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1263 = 8'ha3 == r_count_4_io_out ? io_r_163_b : _GEN_1262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1264 = 8'ha4 == r_count_4_io_out ? io_r_164_b : _GEN_1263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1265 = 8'ha5 == r_count_4_io_out ? io_r_165_b : _GEN_1264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1266 = 8'ha6 == r_count_4_io_out ? io_r_166_b : _GEN_1265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1267 = 8'ha7 == r_count_4_io_out ? io_r_167_b : _GEN_1266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1268 = 8'ha8 == r_count_4_io_out ? io_r_168_b : _GEN_1267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1269 = 8'ha9 == r_count_4_io_out ? io_r_169_b : _GEN_1268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1270 = 8'haa == r_count_4_io_out ? io_r_170_b : _GEN_1269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1271 = 8'hab == r_count_4_io_out ? io_r_171_b : _GEN_1270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1272 = 8'hac == r_count_4_io_out ? io_r_172_b : _GEN_1271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1273 = 8'had == r_count_4_io_out ? io_r_173_b : _GEN_1272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1274 = 8'hae == r_count_4_io_out ? io_r_174_b : _GEN_1273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1275 = 8'haf == r_count_4_io_out ? io_r_175_b : _GEN_1274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1276 = 8'hb0 == r_count_4_io_out ? io_r_176_b : _GEN_1275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1277 = 8'hb1 == r_count_4_io_out ? io_r_177_b : _GEN_1276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1278 = 8'hb2 == r_count_4_io_out ? io_r_178_b : _GEN_1277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1279 = 8'hb3 == r_count_4_io_out ? io_r_179_b : _GEN_1278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1280 = 8'hb4 == r_count_4_io_out ? io_r_180_b : _GEN_1279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1281 = 8'hb5 == r_count_4_io_out ? io_r_181_b : _GEN_1280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1282 = 8'hb6 == r_count_4_io_out ? io_r_182_b : _GEN_1281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1283 = 8'hb7 == r_count_4_io_out ? io_r_183_b : _GEN_1282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1284 = 8'hb8 == r_count_4_io_out ? io_r_184_b : _GEN_1283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1285 = 8'hb9 == r_count_4_io_out ? io_r_185_b : _GEN_1284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1286 = 8'hba == r_count_4_io_out ? io_r_186_b : _GEN_1285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1287 = 8'hbb == r_count_4_io_out ? io_r_187_b : _GEN_1286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1288 = 8'hbc == r_count_4_io_out ? io_r_188_b : _GEN_1287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1289 = 8'hbd == r_count_4_io_out ? io_r_189_b : _GEN_1288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1290 = 8'hbe == r_count_4_io_out ? io_r_190_b : _GEN_1289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1291 = 8'hbf == r_count_4_io_out ? io_r_191_b : _GEN_1290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1292 = 8'hc0 == r_count_4_io_out ? io_r_192_b : _GEN_1291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1293 = 8'hc1 == r_count_4_io_out ? io_r_193_b : _GEN_1292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1294 = 8'hc2 == r_count_4_io_out ? io_r_194_b : _GEN_1293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1295 = 8'hc3 == r_count_4_io_out ? io_r_195_b : _GEN_1294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1296 = 8'hc4 == r_count_4_io_out ? io_r_196_b : _GEN_1295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1297 = 8'hc5 == r_count_4_io_out ? io_r_197_b : _GEN_1296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1298 = 8'hc6 == r_count_4_io_out ? io_r_198_b : _GEN_1297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1301 = 8'h1 == r_count_5_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1302 = 8'h2 == r_count_5_io_out ? io_r_2_b : _GEN_1301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1303 = 8'h3 == r_count_5_io_out ? io_r_3_b : _GEN_1302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1304 = 8'h4 == r_count_5_io_out ? io_r_4_b : _GEN_1303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1305 = 8'h5 == r_count_5_io_out ? io_r_5_b : _GEN_1304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1306 = 8'h6 == r_count_5_io_out ? io_r_6_b : _GEN_1305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1307 = 8'h7 == r_count_5_io_out ? io_r_7_b : _GEN_1306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1308 = 8'h8 == r_count_5_io_out ? io_r_8_b : _GEN_1307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1309 = 8'h9 == r_count_5_io_out ? io_r_9_b : _GEN_1308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1310 = 8'ha == r_count_5_io_out ? io_r_10_b : _GEN_1309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1311 = 8'hb == r_count_5_io_out ? io_r_11_b : _GEN_1310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1312 = 8'hc == r_count_5_io_out ? io_r_12_b : _GEN_1311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1313 = 8'hd == r_count_5_io_out ? io_r_13_b : _GEN_1312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1314 = 8'he == r_count_5_io_out ? io_r_14_b : _GEN_1313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1315 = 8'hf == r_count_5_io_out ? io_r_15_b : _GEN_1314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1316 = 8'h10 == r_count_5_io_out ? io_r_16_b : _GEN_1315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1317 = 8'h11 == r_count_5_io_out ? io_r_17_b : _GEN_1316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1318 = 8'h12 == r_count_5_io_out ? io_r_18_b : _GEN_1317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1319 = 8'h13 == r_count_5_io_out ? io_r_19_b : _GEN_1318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1320 = 8'h14 == r_count_5_io_out ? io_r_20_b : _GEN_1319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1321 = 8'h15 == r_count_5_io_out ? io_r_21_b : _GEN_1320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1322 = 8'h16 == r_count_5_io_out ? io_r_22_b : _GEN_1321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1323 = 8'h17 == r_count_5_io_out ? io_r_23_b : _GEN_1322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1324 = 8'h18 == r_count_5_io_out ? io_r_24_b : _GEN_1323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1325 = 8'h19 == r_count_5_io_out ? io_r_25_b : _GEN_1324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1326 = 8'h1a == r_count_5_io_out ? io_r_26_b : _GEN_1325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1327 = 8'h1b == r_count_5_io_out ? io_r_27_b : _GEN_1326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1328 = 8'h1c == r_count_5_io_out ? io_r_28_b : _GEN_1327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1329 = 8'h1d == r_count_5_io_out ? io_r_29_b : _GEN_1328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1330 = 8'h1e == r_count_5_io_out ? io_r_30_b : _GEN_1329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1331 = 8'h1f == r_count_5_io_out ? io_r_31_b : _GEN_1330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1332 = 8'h20 == r_count_5_io_out ? io_r_32_b : _GEN_1331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1333 = 8'h21 == r_count_5_io_out ? io_r_33_b : _GEN_1332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1334 = 8'h22 == r_count_5_io_out ? io_r_34_b : _GEN_1333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1335 = 8'h23 == r_count_5_io_out ? io_r_35_b : _GEN_1334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1336 = 8'h24 == r_count_5_io_out ? io_r_36_b : _GEN_1335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1337 = 8'h25 == r_count_5_io_out ? io_r_37_b : _GEN_1336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1338 = 8'h26 == r_count_5_io_out ? io_r_38_b : _GEN_1337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1339 = 8'h27 == r_count_5_io_out ? io_r_39_b : _GEN_1338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1340 = 8'h28 == r_count_5_io_out ? io_r_40_b : _GEN_1339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1341 = 8'h29 == r_count_5_io_out ? io_r_41_b : _GEN_1340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1342 = 8'h2a == r_count_5_io_out ? io_r_42_b : _GEN_1341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1343 = 8'h2b == r_count_5_io_out ? io_r_43_b : _GEN_1342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1344 = 8'h2c == r_count_5_io_out ? io_r_44_b : _GEN_1343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1345 = 8'h2d == r_count_5_io_out ? io_r_45_b : _GEN_1344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1346 = 8'h2e == r_count_5_io_out ? io_r_46_b : _GEN_1345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1347 = 8'h2f == r_count_5_io_out ? io_r_47_b : _GEN_1346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1348 = 8'h30 == r_count_5_io_out ? io_r_48_b : _GEN_1347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1349 = 8'h31 == r_count_5_io_out ? io_r_49_b : _GEN_1348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1350 = 8'h32 == r_count_5_io_out ? io_r_50_b : _GEN_1349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1351 = 8'h33 == r_count_5_io_out ? io_r_51_b : _GEN_1350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1352 = 8'h34 == r_count_5_io_out ? io_r_52_b : _GEN_1351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1353 = 8'h35 == r_count_5_io_out ? io_r_53_b : _GEN_1352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1354 = 8'h36 == r_count_5_io_out ? io_r_54_b : _GEN_1353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1355 = 8'h37 == r_count_5_io_out ? io_r_55_b : _GEN_1354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1356 = 8'h38 == r_count_5_io_out ? io_r_56_b : _GEN_1355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1357 = 8'h39 == r_count_5_io_out ? io_r_57_b : _GEN_1356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1358 = 8'h3a == r_count_5_io_out ? io_r_58_b : _GEN_1357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1359 = 8'h3b == r_count_5_io_out ? io_r_59_b : _GEN_1358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1360 = 8'h3c == r_count_5_io_out ? io_r_60_b : _GEN_1359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1361 = 8'h3d == r_count_5_io_out ? io_r_61_b : _GEN_1360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1362 = 8'h3e == r_count_5_io_out ? io_r_62_b : _GEN_1361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1363 = 8'h3f == r_count_5_io_out ? io_r_63_b : _GEN_1362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1364 = 8'h40 == r_count_5_io_out ? io_r_64_b : _GEN_1363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1365 = 8'h41 == r_count_5_io_out ? io_r_65_b : _GEN_1364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1366 = 8'h42 == r_count_5_io_out ? io_r_66_b : _GEN_1365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1367 = 8'h43 == r_count_5_io_out ? io_r_67_b : _GEN_1366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1368 = 8'h44 == r_count_5_io_out ? io_r_68_b : _GEN_1367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1369 = 8'h45 == r_count_5_io_out ? io_r_69_b : _GEN_1368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1370 = 8'h46 == r_count_5_io_out ? io_r_70_b : _GEN_1369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1371 = 8'h47 == r_count_5_io_out ? io_r_71_b : _GEN_1370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1372 = 8'h48 == r_count_5_io_out ? io_r_72_b : _GEN_1371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1373 = 8'h49 == r_count_5_io_out ? io_r_73_b : _GEN_1372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1374 = 8'h4a == r_count_5_io_out ? io_r_74_b : _GEN_1373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1375 = 8'h4b == r_count_5_io_out ? io_r_75_b : _GEN_1374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1376 = 8'h4c == r_count_5_io_out ? io_r_76_b : _GEN_1375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1377 = 8'h4d == r_count_5_io_out ? io_r_77_b : _GEN_1376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1378 = 8'h4e == r_count_5_io_out ? io_r_78_b : _GEN_1377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1379 = 8'h4f == r_count_5_io_out ? io_r_79_b : _GEN_1378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1380 = 8'h50 == r_count_5_io_out ? io_r_80_b : _GEN_1379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1381 = 8'h51 == r_count_5_io_out ? io_r_81_b : _GEN_1380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1382 = 8'h52 == r_count_5_io_out ? io_r_82_b : _GEN_1381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1383 = 8'h53 == r_count_5_io_out ? io_r_83_b : _GEN_1382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1384 = 8'h54 == r_count_5_io_out ? io_r_84_b : _GEN_1383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1385 = 8'h55 == r_count_5_io_out ? io_r_85_b : _GEN_1384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1386 = 8'h56 == r_count_5_io_out ? io_r_86_b : _GEN_1385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1387 = 8'h57 == r_count_5_io_out ? io_r_87_b : _GEN_1386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1388 = 8'h58 == r_count_5_io_out ? io_r_88_b : _GEN_1387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1389 = 8'h59 == r_count_5_io_out ? io_r_89_b : _GEN_1388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1390 = 8'h5a == r_count_5_io_out ? io_r_90_b : _GEN_1389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1391 = 8'h5b == r_count_5_io_out ? io_r_91_b : _GEN_1390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1392 = 8'h5c == r_count_5_io_out ? io_r_92_b : _GEN_1391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1393 = 8'h5d == r_count_5_io_out ? io_r_93_b : _GEN_1392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1394 = 8'h5e == r_count_5_io_out ? io_r_94_b : _GEN_1393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1395 = 8'h5f == r_count_5_io_out ? io_r_95_b : _GEN_1394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1396 = 8'h60 == r_count_5_io_out ? io_r_96_b : _GEN_1395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1397 = 8'h61 == r_count_5_io_out ? io_r_97_b : _GEN_1396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1398 = 8'h62 == r_count_5_io_out ? io_r_98_b : _GEN_1397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1399 = 8'h63 == r_count_5_io_out ? io_r_99_b : _GEN_1398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1400 = 8'h64 == r_count_5_io_out ? io_r_100_b : _GEN_1399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1401 = 8'h65 == r_count_5_io_out ? io_r_101_b : _GEN_1400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1402 = 8'h66 == r_count_5_io_out ? io_r_102_b : _GEN_1401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1403 = 8'h67 == r_count_5_io_out ? io_r_103_b : _GEN_1402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1404 = 8'h68 == r_count_5_io_out ? io_r_104_b : _GEN_1403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1405 = 8'h69 == r_count_5_io_out ? io_r_105_b : _GEN_1404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1406 = 8'h6a == r_count_5_io_out ? io_r_106_b : _GEN_1405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1407 = 8'h6b == r_count_5_io_out ? io_r_107_b : _GEN_1406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1408 = 8'h6c == r_count_5_io_out ? io_r_108_b : _GEN_1407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1409 = 8'h6d == r_count_5_io_out ? io_r_109_b : _GEN_1408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1410 = 8'h6e == r_count_5_io_out ? io_r_110_b : _GEN_1409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1411 = 8'h6f == r_count_5_io_out ? io_r_111_b : _GEN_1410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1412 = 8'h70 == r_count_5_io_out ? io_r_112_b : _GEN_1411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1413 = 8'h71 == r_count_5_io_out ? io_r_113_b : _GEN_1412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1414 = 8'h72 == r_count_5_io_out ? io_r_114_b : _GEN_1413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1415 = 8'h73 == r_count_5_io_out ? io_r_115_b : _GEN_1414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1416 = 8'h74 == r_count_5_io_out ? io_r_116_b : _GEN_1415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1417 = 8'h75 == r_count_5_io_out ? io_r_117_b : _GEN_1416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1418 = 8'h76 == r_count_5_io_out ? io_r_118_b : _GEN_1417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1419 = 8'h77 == r_count_5_io_out ? io_r_119_b : _GEN_1418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1420 = 8'h78 == r_count_5_io_out ? io_r_120_b : _GEN_1419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1421 = 8'h79 == r_count_5_io_out ? io_r_121_b : _GEN_1420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1422 = 8'h7a == r_count_5_io_out ? io_r_122_b : _GEN_1421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1423 = 8'h7b == r_count_5_io_out ? io_r_123_b : _GEN_1422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1424 = 8'h7c == r_count_5_io_out ? io_r_124_b : _GEN_1423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1425 = 8'h7d == r_count_5_io_out ? io_r_125_b : _GEN_1424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1426 = 8'h7e == r_count_5_io_out ? io_r_126_b : _GEN_1425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1427 = 8'h7f == r_count_5_io_out ? io_r_127_b : _GEN_1426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1428 = 8'h80 == r_count_5_io_out ? io_r_128_b : _GEN_1427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1429 = 8'h81 == r_count_5_io_out ? io_r_129_b : _GEN_1428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1430 = 8'h82 == r_count_5_io_out ? io_r_130_b : _GEN_1429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1431 = 8'h83 == r_count_5_io_out ? io_r_131_b : _GEN_1430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1432 = 8'h84 == r_count_5_io_out ? io_r_132_b : _GEN_1431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1433 = 8'h85 == r_count_5_io_out ? io_r_133_b : _GEN_1432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1434 = 8'h86 == r_count_5_io_out ? io_r_134_b : _GEN_1433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1435 = 8'h87 == r_count_5_io_out ? io_r_135_b : _GEN_1434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1436 = 8'h88 == r_count_5_io_out ? io_r_136_b : _GEN_1435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1437 = 8'h89 == r_count_5_io_out ? io_r_137_b : _GEN_1436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1438 = 8'h8a == r_count_5_io_out ? io_r_138_b : _GEN_1437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1439 = 8'h8b == r_count_5_io_out ? io_r_139_b : _GEN_1438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1440 = 8'h8c == r_count_5_io_out ? io_r_140_b : _GEN_1439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1441 = 8'h8d == r_count_5_io_out ? io_r_141_b : _GEN_1440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1442 = 8'h8e == r_count_5_io_out ? io_r_142_b : _GEN_1441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1443 = 8'h8f == r_count_5_io_out ? io_r_143_b : _GEN_1442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1444 = 8'h90 == r_count_5_io_out ? io_r_144_b : _GEN_1443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1445 = 8'h91 == r_count_5_io_out ? io_r_145_b : _GEN_1444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1446 = 8'h92 == r_count_5_io_out ? io_r_146_b : _GEN_1445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1447 = 8'h93 == r_count_5_io_out ? io_r_147_b : _GEN_1446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1448 = 8'h94 == r_count_5_io_out ? io_r_148_b : _GEN_1447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1449 = 8'h95 == r_count_5_io_out ? io_r_149_b : _GEN_1448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1450 = 8'h96 == r_count_5_io_out ? io_r_150_b : _GEN_1449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1451 = 8'h97 == r_count_5_io_out ? io_r_151_b : _GEN_1450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1452 = 8'h98 == r_count_5_io_out ? io_r_152_b : _GEN_1451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1453 = 8'h99 == r_count_5_io_out ? io_r_153_b : _GEN_1452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1454 = 8'h9a == r_count_5_io_out ? io_r_154_b : _GEN_1453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1455 = 8'h9b == r_count_5_io_out ? io_r_155_b : _GEN_1454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1456 = 8'h9c == r_count_5_io_out ? io_r_156_b : _GEN_1455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1457 = 8'h9d == r_count_5_io_out ? io_r_157_b : _GEN_1456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1458 = 8'h9e == r_count_5_io_out ? io_r_158_b : _GEN_1457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1459 = 8'h9f == r_count_5_io_out ? io_r_159_b : _GEN_1458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1460 = 8'ha0 == r_count_5_io_out ? io_r_160_b : _GEN_1459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1461 = 8'ha1 == r_count_5_io_out ? io_r_161_b : _GEN_1460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1462 = 8'ha2 == r_count_5_io_out ? io_r_162_b : _GEN_1461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1463 = 8'ha3 == r_count_5_io_out ? io_r_163_b : _GEN_1462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1464 = 8'ha4 == r_count_5_io_out ? io_r_164_b : _GEN_1463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1465 = 8'ha5 == r_count_5_io_out ? io_r_165_b : _GEN_1464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1466 = 8'ha6 == r_count_5_io_out ? io_r_166_b : _GEN_1465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1467 = 8'ha7 == r_count_5_io_out ? io_r_167_b : _GEN_1466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1468 = 8'ha8 == r_count_5_io_out ? io_r_168_b : _GEN_1467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1469 = 8'ha9 == r_count_5_io_out ? io_r_169_b : _GEN_1468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1470 = 8'haa == r_count_5_io_out ? io_r_170_b : _GEN_1469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1471 = 8'hab == r_count_5_io_out ? io_r_171_b : _GEN_1470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1472 = 8'hac == r_count_5_io_out ? io_r_172_b : _GEN_1471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1473 = 8'had == r_count_5_io_out ? io_r_173_b : _GEN_1472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1474 = 8'hae == r_count_5_io_out ? io_r_174_b : _GEN_1473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1475 = 8'haf == r_count_5_io_out ? io_r_175_b : _GEN_1474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1476 = 8'hb0 == r_count_5_io_out ? io_r_176_b : _GEN_1475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1477 = 8'hb1 == r_count_5_io_out ? io_r_177_b : _GEN_1476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1478 = 8'hb2 == r_count_5_io_out ? io_r_178_b : _GEN_1477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1479 = 8'hb3 == r_count_5_io_out ? io_r_179_b : _GEN_1478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1480 = 8'hb4 == r_count_5_io_out ? io_r_180_b : _GEN_1479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1481 = 8'hb5 == r_count_5_io_out ? io_r_181_b : _GEN_1480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1482 = 8'hb6 == r_count_5_io_out ? io_r_182_b : _GEN_1481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1483 = 8'hb7 == r_count_5_io_out ? io_r_183_b : _GEN_1482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1484 = 8'hb8 == r_count_5_io_out ? io_r_184_b : _GEN_1483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1485 = 8'hb9 == r_count_5_io_out ? io_r_185_b : _GEN_1484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1486 = 8'hba == r_count_5_io_out ? io_r_186_b : _GEN_1485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1487 = 8'hbb == r_count_5_io_out ? io_r_187_b : _GEN_1486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1488 = 8'hbc == r_count_5_io_out ? io_r_188_b : _GEN_1487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1489 = 8'hbd == r_count_5_io_out ? io_r_189_b : _GEN_1488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1490 = 8'hbe == r_count_5_io_out ? io_r_190_b : _GEN_1489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1491 = 8'hbf == r_count_5_io_out ? io_r_191_b : _GEN_1490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1492 = 8'hc0 == r_count_5_io_out ? io_r_192_b : _GEN_1491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1493 = 8'hc1 == r_count_5_io_out ? io_r_193_b : _GEN_1492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1494 = 8'hc2 == r_count_5_io_out ? io_r_194_b : _GEN_1493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1495 = 8'hc3 == r_count_5_io_out ? io_r_195_b : _GEN_1494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1496 = 8'hc4 == r_count_5_io_out ? io_r_196_b : _GEN_1495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1497 = 8'hc5 == r_count_5_io_out ? io_r_197_b : _GEN_1496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1498 = 8'hc6 == r_count_5_io_out ? io_r_198_b : _GEN_1497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1501 = 8'h1 == r_count_6_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1502 = 8'h2 == r_count_6_io_out ? io_r_2_b : _GEN_1501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1503 = 8'h3 == r_count_6_io_out ? io_r_3_b : _GEN_1502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1504 = 8'h4 == r_count_6_io_out ? io_r_4_b : _GEN_1503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1505 = 8'h5 == r_count_6_io_out ? io_r_5_b : _GEN_1504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1506 = 8'h6 == r_count_6_io_out ? io_r_6_b : _GEN_1505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1507 = 8'h7 == r_count_6_io_out ? io_r_7_b : _GEN_1506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1508 = 8'h8 == r_count_6_io_out ? io_r_8_b : _GEN_1507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1509 = 8'h9 == r_count_6_io_out ? io_r_9_b : _GEN_1508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1510 = 8'ha == r_count_6_io_out ? io_r_10_b : _GEN_1509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1511 = 8'hb == r_count_6_io_out ? io_r_11_b : _GEN_1510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1512 = 8'hc == r_count_6_io_out ? io_r_12_b : _GEN_1511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1513 = 8'hd == r_count_6_io_out ? io_r_13_b : _GEN_1512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1514 = 8'he == r_count_6_io_out ? io_r_14_b : _GEN_1513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1515 = 8'hf == r_count_6_io_out ? io_r_15_b : _GEN_1514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1516 = 8'h10 == r_count_6_io_out ? io_r_16_b : _GEN_1515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1517 = 8'h11 == r_count_6_io_out ? io_r_17_b : _GEN_1516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1518 = 8'h12 == r_count_6_io_out ? io_r_18_b : _GEN_1517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1519 = 8'h13 == r_count_6_io_out ? io_r_19_b : _GEN_1518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1520 = 8'h14 == r_count_6_io_out ? io_r_20_b : _GEN_1519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1521 = 8'h15 == r_count_6_io_out ? io_r_21_b : _GEN_1520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1522 = 8'h16 == r_count_6_io_out ? io_r_22_b : _GEN_1521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1523 = 8'h17 == r_count_6_io_out ? io_r_23_b : _GEN_1522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1524 = 8'h18 == r_count_6_io_out ? io_r_24_b : _GEN_1523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1525 = 8'h19 == r_count_6_io_out ? io_r_25_b : _GEN_1524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1526 = 8'h1a == r_count_6_io_out ? io_r_26_b : _GEN_1525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1527 = 8'h1b == r_count_6_io_out ? io_r_27_b : _GEN_1526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1528 = 8'h1c == r_count_6_io_out ? io_r_28_b : _GEN_1527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1529 = 8'h1d == r_count_6_io_out ? io_r_29_b : _GEN_1528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1530 = 8'h1e == r_count_6_io_out ? io_r_30_b : _GEN_1529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1531 = 8'h1f == r_count_6_io_out ? io_r_31_b : _GEN_1530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1532 = 8'h20 == r_count_6_io_out ? io_r_32_b : _GEN_1531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1533 = 8'h21 == r_count_6_io_out ? io_r_33_b : _GEN_1532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1534 = 8'h22 == r_count_6_io_out ? io_r_34_b : _GEN_1533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1535 = 8'h23 == r_count_6_io_out ? io_r_35_b : _GEN_1534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1536 = 8'h24 == r_count_6_io_out ? io_r_36_b : _GEN_1535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1537 = 8'h25 == r_count_6_io_out ? io_r_37_b : _GEN_1536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1538 = 8'h26 == r_count_6_io_out ? io_r_38_b : _GEN_1537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1539 = 8'h27 == r_count_6_io_out ? io_r_39_b : _GEN_1538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1540 = 8'h28 == r_count_6_io_out ? io_r_40_b : _GEN_1539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1541 = 8'h29 == r_count_6_io_out ? io_r_41_b : _GEN_1540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1542 = 8'h2a == r_count_6_io_out ? io_r_42_b : _GEN_1541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1543 = 8'h2b == r_count_6_io_out ? io_r_43_b : _GEN_1542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1544 = 8'h2c == r_count_6_io_out ? io_r_44_b : _GEN_1543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1545 = 8'h2d == r_count_6_io_out ? io_r_45_b : _GEN_1544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1546 = 8'h2e == r_count_6_io_out ? io_r_46_b : _GEN_1545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1547 = 8'h2f == r_count_6_io_out ? io_r_47_b : _GEN_1546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1548 = 8'h30 == r_count_6_io_out ? io_r_48_b : _GEN_1547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1549 = 8'h31 == r_count_6_io_out ? io_r_49_b : _GEN_1548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1550 = 8'h32 == r_count_6_io_out ? io_r_50_b : _GEN_1549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1551 = 8'h33 == r_count_6_io_out ? io_r_51_b : _GEN_1550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1552 = 8'h34 == r_count_6_io_out ? io_r_52_b : _GEN_1551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1553 = 8'h35 == r_count_6_io_out ? io_r_53_b : _GEN_1552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1554 = 8'h36 == r_count_6_io_out ? io_r_54_b : _GEN_1553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1555 = 8'h37 == r_count_6_io_out ? io_r_55_b : _GEN_1554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1556 = 8'h38 == r_count_6_io_out ? io_r_56_b : _GEN_1555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1557 = 8'h39 == r_count_6_io_out ? io_r_57_b : _GEN_1556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1558 = 8'h3a == r_count_6_io_out ? io_r_58_b : _GEN_1557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1559 = 8'h3b == r_count_6_io_out ? io_r_59_b : _GEN_1558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1560 = 8'h3c == r_count_6_io_out ? io_r_60_b : _GEN_1559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1561 = 8'h3d == r_count_6_io_out ? io_r_61_b : _GEN_1560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1562 = 8'h3e == r_count_6_io_out ? io_r_62_b : _GEN_1561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1563 = 8'h3f == r_count_6_io_out ? io_r_63_b : _GEN_1562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1564 = 8'h40 == r_count_6_io_out ? io_r_64_b : _GEN_1563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1565 = 8'h41 == r_count_6_io_out ? io_r_65_b : _GEN_1564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1566 = 8'h42 == r_count_6_io_out ? io_r_66_b : _GEN_1565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1567 = 8'h43 == r_count_6_io_out ? io_r_67_b : _GEN_1566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1568 = 8'h44 == r_count_6_io_out ? io_r_68_b : _GEN_1567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1569 = 8'h45 == r_count_6_io_out ? io_r_69_b : _GEN_1568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1570 = 8'h46 == r_count_6_io_out ? io_r_70_b : _GEN_1569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1571 = 8'h47 == r_count_6_io_out ? io_r_71_b : _GEN_1570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1572 = 8'h48 == r_count_6_io_out ? io_r_72_b : _GEN_1571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1573 = 8'h49 == r_count_6_io_out ? io_r_73_b : _GEN_1572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1574 = 8'h4a == r_count_6_io_out ? io_r_74_b : _GEN_1573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1575 = 8'h4b == r_count_6_io_out ? io_r_75_b : _GEN_1574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1576 = 8'h4c == r_count_6_io_out ? io_r_76_b : _GEN_1575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1577 = 8'h4d == r_count_6_io_out ? io_r_77_b : _GEN_1576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1578 = 8'h4e == r_count_6_io_out ? io_r_78_b : _GEN_1577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1579 = 8'h4f == r_count_6_io_out ? io_r_79_b : _GEN_1578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1580 = 8'h50 == r_count_6_io_out ? io_r_80_b : _GEN_1579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1581 = 8'h51 == r_count_6_io_out ? io_r_81_b : _GEN_1580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1582 = 8'h52 == r_count_6_io_out ? io_r_82_b : _GEN_1581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1583 = 8'h53 == r_count_6_io_out ? io_r_83_b : _GEN_1582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1584 = 8'h54 == r_count_6_io_out ? io_r_84_b : _GEN_1583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1585 = 8'h55 == r_count_6_io_out ? io_r_85_b : _GEN_1584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1586 = 8'h56 == r_count_6_io_out ? io_r_86_b : _GEN_1585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1587 = 8'h57 == r_count_6_io_out ? io_r_87_b : _GEN_1586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1588 = 8'h58 == r_count_6_io_out ? io_r_88_b : _GEN_1587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1589 = 8'h59 == r_count_6_io_out ? io_r_89_b : _GEN_1588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1590 = 8'h5a == r_count_6_io_out ? io_r_90_b : _GEN_1589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1591 = 8'h5b == r_count_6_io_out ? io_r_91_b : _GEN_1590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1592 = 8'h5c == r_count_6_io_out ? io_r_92_b : _GEN_1591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1593 = 8'h5d == r_count_6_io_out ? io_r_93_b : _GEN_1592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1594 = 8'h5e == r_count_6_io_out ? io_r_94_b : _GEN_1593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1595 = 8'h5f == r_count_6_io_out ? io_r_95_b : _GEN_1594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1596 = 8'h60 == r_count_6_io_out ? io_r_96_b : _GEN_1595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1597 = 8'h61 == r_count_6_io_out ? io_r_97_b : _GEN_1596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1598 = 8'h62 == r_count_6_io_out ? io_r_98_b : _GEN_1597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1599 = 8'h63 == r_count_6_io_out ? io_r_99_b : _GEN_1598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1600 = 8'h64 == r_count_6_io_out ? io_r_100_b : _GEN_1599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1601 = 8'h65 == r_count_6_io_out ? io_r_101_b : _GEN_1600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1602 = 8'h66 == r_count_6_io_out ? io_r_102_b : _GEN_1601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1603 = 8'h67 == r_count_6_io_out ? io_r_103_b : _GEN_1602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1604 = 8'h68 == r_count_6_io_out ? io_r_104_b : _GEN_1603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1605 = 8'h69 == r_count_6_io_out ? io_r_105_b : _GEN_1604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1606 = 8'h6a == r_count_6_io_out ? io_r_106_b : _GEN_1605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1607 = 8'h6b == r_count_6_io_out ? io_r_107_b : _GEN_1606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1608 = 8'h6c == r_count_6_io_out ? io_r_108_b : _GEN_1607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1609 = 8'h6d == r_count_6_io_out ? io_r_109_b : _GEN_1608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1610 = 8'h6e == r_count_6_io_out ? io_r_110_b : _GEN_1609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1611 = 8'h6f == r_count_6_io_out ? io_r_111_b : _GEN_1610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1612 = 8'h70 == r_count_6_io_out ? io_r_112_b : _GEN_1611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1613 = 8'h71 == r_count_6_io_out ? io_r_113_b : _GEN_1612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1614 = 8'h72 == r_count_6_io_out ? io_r_114_b : _GEN_1613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1615 = 8'h73 == r_count_6_io_out ? io_r_115_b : _GEN_1614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1616 = 8'h74 == r_count_6_io_out ? io_r_116_b : _GEN_1615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1617 = 8'h75 == r_count_6_io_out ? io_r_117_b : _GEN_1616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1618 = 8'h76 == r_count_6_io_out ? io_r_118_b : _GEN_1617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1619 = 8'h77 == r_count_6_io_out ? io_r_119_b : _GEN_1618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1620 = 8'h78 == r_count_6_io_out ? io_r_120_b : _GEN_1619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1621 = 8'h79 == r_count_6_io_out ? io_r_121_b : _GEN_1620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1622 = 8'h7a == r_count_6_io_out ? io_r_122_b : _GEN_1621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1623 = 8'h7b == r_count_6_io_out ? io_r_123_b : _GEN_1622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1624 = 8'h7c == r_count_6_io_out ? io_r_124_b : _GEN_1623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1625 = 8'h7d == r_count_6_io_out ? io_r_125_b : _GEN_1624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1626 = 8'h7e == r_count_6_io_out ? io_r_126_b : _GEN_1625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1627 = 8'h7f == r_count_6_io_out ? io_r_127_b : _GEN_1626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1628 = 8'h80 == r_count_6_io_out ? io_r_128_b : _GEN_1627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1629 = 8'h81 == r_count_6_io_out ? io_r_129_b : _GEN_1628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1630 = 8'h82 == r_count_6_io_out ? io_r_130_b : _GEN_1629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1631 = 8'h83 == r_count_6_io_out ? io_r_131_b : _GEN_1630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1632 = 8'h84 == r_count_6_io_out ? io_r_132_b : _GEN_1631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1633 = 8'h85 == r_count_6_io_out ? io_r_133_b : _GEN_1632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1634 = 8'h86 == r_count_6_io_out ? io_r_134_b : _GEN_1633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1635 = 8'h87 == r_count_6_io_out ? io_r_135_b : _GEN_1634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1636 = 8'h88 == r_count_6_io_out ? io_r_136_b : _GEN_1635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1637 = 8'h89 == r_count_6_io_out ? io_r_137_b : _GEN_1636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1638 = 8'h8a == r_count_6_io_out ? io_r_138_b : _GEN_1637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1639 = 8'h8b == r_count_6_io_out ? io_r_139_b : _GEN_1638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1640 = 8'h8c == r_count_6_io_out ? io_r_140_b : _GEN_1639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1641 = 8'h8d == r_count_6_io_out ? io_r_141_b : _GEN_1640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1642 = 8'h8e == r_count_6_io_out ? io_r_142_b : _GEN_1641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1643 = 8'h8f == r_count_6_io_out ? io_r_143_b : _GEN_1642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1644 = 8'h90 == r_count_6_io_out ? io_r_144_b : _GEN_1643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1645 = 8'h91 == r_count_6_io_out ? io_r_145_b : _GEN_1644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1646 = 8'h92 == r_count_6_io_out ? io_r_146_b : _GEN_1645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1647 = 8'h93 == r_count_6_io_out ? io_r_147_b : _GEN_1646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1648 = 8'h94 == r_count_6_io_out ? io_r_148_b : _GEN_1647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1649 = 8'h95 == r_count_6_io_out ? io_r_149_b : _GEN_1648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1650 = 8'h96 == r_count_6_io_out ? io_r_150_b : _GEN_1649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1651 = 8'h97 == r_count_6_io_out ? io_r_151_b : _GEN_1650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1652 = 8'h98 == r_count_6_io_out ? io_r_152_b : _GEN_1651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1653 = 8'h99 == r_count_6_io_out ? io_r_153_b : _GEN_1652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1654 = 8'h9a == r_count_6_io_out ? io_r_154_b : _GEN_1653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1655 = 8'h9b == r_count_6_io_out ? io_r_155_b : _GEN_1654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1656 = 8'h9c == r_count_6_io_out ? io_r_156_b : _GEN_1655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1657 = 8'h9d == r_count_6_io_out ? io_r_157_b : _GEN_1656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1658 = 8'h9e == r_count_6_io_out ? io_r_158_b : _GEN_1657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1659 = 8'h9f == r_count_6_io_out ? io_r_159_b : _GEN_1658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1660 = 8'ha0 == r_count_6_io_out ? io_r_160_b : _GEN_1659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1661 = 8'ha1 == r_count_6_io_out ? io_r_161_b : _GEN_1660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1662 = 8'ha2 == r_count_6_io_out ? io_r_162_b : _GEN_1661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1663 = 8'ha3 == r_count_6_io_out ? io_r_163_b : _GEN_1662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1664 = 8'ha4 == r_count_6_io_out ? io_r_164_b : _GEN_1663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1665 = 8'ha5 == r_count_6_io_out ? io_r_165_b : _GEN_1664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1666 = 8'ha6 == r_count_6_io_out ? io_r_166_b : _GEN_1665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1667 = 8'ha7 == r_count_6_io_out ? io_r_167_b : _GEN_1666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1668 = 8'ha8 == r_count_6_io_out ? io_r_168_b : _GEN_1667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1669 = 8'ha9 == r_count_6_io_out ? io_r_169_b : _GEN_1668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1670 = 8'haa == r_count_6_io_out ? io_r_170_b : _GEN_1669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1671 = 8'hab == r_count_6_io_out ? io_r_171_b : _GEN_1670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1672 = 8'hac == r_count_6_io_out ? io_r_172_b : _GEN_1671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1673 = 8'had == r_count_6_io_out ? io_r_173_b : _GEN_1672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1674 = 8'hae == r_count_6_io_out ? io_r_174_b : _GEN_1673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1675 = 8'haf == r_count_6_io_out ? io_r_175_b : _GEN_1674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1676 = 8'hb0 == r_count_6_io_out ? io_r_176_b : _GEN_1675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1677 = 8'hb1 == r_count_6_io_out ? io_r_177_b : _GEN_1676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1678 = 8'hb2 == r_count_6_io_out ? io_r_178_b : _GEN_1677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1679 = 8'hb3 == r_count_6_io_out ? io_r_179_b : _GEN_1678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1680 = 8'hb4 == r_count_6_io_out ? io_r_180_b : _GEN_1679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1681 = 8'hb5 == r_count_6_io_out ? io_r_181_b : _GEN_1680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1682 = 8'hb6 == r_count_6_io_out ? io_r_182_b : _GEN_1681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1683 = 8'hb7 == r_count_6_io_out ? io_r_183_b : _GEN_1682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1684 = 8'hb8 == r_count_6_io_out ? io_r_184_b : _GEN_1683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1685 = 8'hb9 == r_count_6_io_out ? io_r_185_b : _GEN_1684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1686 = 8'hba == r_count_6_io_out ? io_r_186_b : _GEN_1685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1687 = 8'hbb == r_count_6_io_out ? io_r_187_b : _GEN_1686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1688 = 8'hbc == r_count_6_io_out ? io_r_188_b : _GEN_1687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1689 = 8'hbd == r_count_6_io_out ? io_r_189_b : _GEN_1688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1690 = 8'hbe == r_count_6_io_out ? io_r_190_b : _GEN_1689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1691 = 8'hbf == r_count_6_io_out ? io_r_191_b : _GEN_1690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1692 = 8'hc0 == r_count_6_io_out ? io_r_192_b : _GEN_1691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1693 = 8'hc1 == r_count_6_io_out ? io_r_193_b : _GEN_1692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1694 = 8'hc2 == r_count_6_io_out ? io_r_194_b : _GEN_1693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1695 = 8'hc3 == r_count_6_io_out ? io_r_195_b : _GEN_1694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1696 = 8'hc4 == r_count_6_io_out ? io_r_196_b : _GEN_1695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1697 = 8'hc5 == r_count_6_io_out ? io_r_197_b : _GEN_1696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1698 = 8'hc6 == r_count_6_io_out ? io_r_198_b : _GEN_1697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1701 = 8'h1 == r_count_7_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1702 = 8'h2 == r_count_7_io_out ? io_r_2_b : _GEN_1701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1703 = 8'h3 == r_count_7_io_out ? io_r_3_b : _GEN_1702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1704 = 8'h4 == r_count_7_io_out ? io_r_4_b : _GEN_1703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1705 = 8'h5 == r_count_7_io_out ? io_r_5_b : _GEN_1704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1706 = 8'h6 == r_count_7_io_out ? io_r_6_b : _GEN_1705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1707 = 8'h7 == r_count_7_io_out ? io_r_7_b : _GEN_1706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1708 = 8'h8 == r_count_7_io_out ? io_r_8_b : _GEN_1707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1709 = 8'h9 == r_count_7_io_out ? io_r_9_b : _GEN_1708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1710 = 8'ha == r_count_7_io_out ? io_r_10_b : _GEN_1709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1711 = 8'hb == r_count_7_io_out ? io_r_11_b : _GEN_1710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1712 = 8'hc == r_count_7_io_out ? io_r_12_b : _GEN_1711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1713 = 8'hd == r_count_7_io_out ? io_r_13_b : _GEN_1712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1714 = 8'he == r_count_7_io_out ? io_r_14_b : _GEN_1713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1715 = 8'hf == r_count_7_io_out ? io_r_15_b : _GEN_1714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1716 = 8'h10 == r_count_7_io_out ? io_r_16_b : _GEN_1715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1717 = 8'h11 == r_count_7_io_out ? io_r_17_b : _GEN_1716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1718 = 8'h12 == r_count_7_io_out ? io_r_18_b : _GEN_1717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1719 = 8'h13 == r_count_7_io_out ? io_r_19_b : _GEN_1718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1720 = 8'h14 == r_count_7_io_out ? io_r_20_b : _GEN_1719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1721 = 8'h15 == r_count_7_io_out ? io_r_21_b : _GEN_1720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1722 = 8'h16 == r_count_7_io_out ? io_r_22_b : _GEN_1721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1723 = 8'h17 == r_count_7_io_out ? io_r_23_b : _GEN_1722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1724 = 8'h18 == r_count_7_io_out ? io_r_24_b : _GEN_1723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1725 = 8'h19 == r_count_7_io_out ? io_r_25_b : _GEN_1724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1726 = 8'h1a == r_count_7_io_out ? io_r_26_b : _GEN_1725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1727 = 8'h1b == r_count_7_io_out ? io_r_27_b : _GEN_1726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1728 = 8'h1c == r_count_7_io_out ? io_r_28_b : _GEN_1727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1729 = 8'h1d == r_count_7_io_out ? io_r_29_b : _GEN_1728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1730 = 8'h1e == r_count_7_io_out ? io_r_30_b : _GEN_1729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1731 = 8'h1f == r_count_7_io_out ? io_r_31_b : _GEN_1730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1732 = 8'h20 == r_count_7_io_out ? io_r_32_b : _GEN_1731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1733 = 8'h21 == r_count_7_io_out ? io_r_33_b : _GEN_1732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1734 = 8'h22 == r_count_7_io_out ? io_r_34_b : _GEN_1733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1735 = 8'h23 == r_count_7_io_out ? io_r_35_b : _GEN_1734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1736 = 8'h24 == r_count_7_io_out ? io_r_36_b : _GEN_1735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1737 = 8'h25 == r_count_7_io_out ? io_r_37_b : _GEN_1736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1738 = 8'h26 == r_count_7_io_out ? io_r_38_b : _GEN_1737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1739 = 8'h27 == r_count_7_io_out ? io_r_39_b : _GEN_1738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1740 = 8'h28 == r_count_7_io_out ? io_r_40_b : _GEN_1739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1741 = 8'h29 == r_count_7_io_out ? io_r_41_b : _GEN_1740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1742 = 8'h2a == r_count_7_io_out ? io_r_42_b : _GEN_1741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1743 = 8'h2b == r_count_7_io_out ? io_r_43_b : _GEN_1742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1744 = 8'h2c == r_count_7_io_out ? io_r_44_b : _GEN_1743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1745 = 8'h2d == r_count_7_io_out ? io_r_45_b : _GEN_1744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1746 = 8'h2e == r_count_7_io_out ? io_r_46_b : _GEN_1745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1747 = 8'h2f == r_count_7_io_out ? io_r_47_b : _GEN_1746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1748 = 8'h30 == r_count_7_io_out ? io_r_48_b : _GEN_1747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1749 = 8'h31 == r_count_7_io_out ? io_r_49_b : _GEN_1748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1750 = 8'h32 == r_count_7_io_out ? io_r_50_b : _GEN_1749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1751 = 8'h33 == r_count_7_io_out ? io_r_51_b : _GEN_1750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1752 = 8'h34 == r_count_7_io_out ? io_r_52_b : _GEN_1751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1753 = 8'h35 == r_count_7_io_out ? io_r_53_b : _GEN_1752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1754 = 8'h36 == r_count_7_io_out ? io_r_54_b : _GEN_1753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1755 = 8'h37 == r_count_7_io_out ? io_r_55_b : _GEN_1754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1756 = 8'h38 == r_count_7_io_out ? io_r_56_b : _GEN_1755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1757 = 8'h39 == r_count_7_io_out ? io_r_57_b : _GEN_1756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1758 = 8'h3a == r_count_7_io_out ? io_r_58_b : _GEN_1757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1759 = 8'h3b == r_count_7_io_out ? io_r_59_b : _GEN_1758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1760 = 8'h3c == r_count_7_io_out ? io_r_60_b : _GEN_1759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1761 = 8'h3d == r_count_7_io_out ? io_r_61_b : _GEN_1760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1762 = 8'h3e == r_count_7_io_out ? io_r_62_b : _GEN_1761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1763 = 8'h3f == r_count_7_io_out ? io_r_63_b : _GEN_1762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1764 = 8'h40 == r_count_7_io_out ? io_r_64_b : _GEN_1763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1765 = 8'h41 == r_count_7_io_out ? io_r_65_b : _GEN_1764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1766 = 8'h42 == r_count_7_io_out ? io_r_66_b : _GEN_1765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1767 = 8'h43 == r_count_7_io_out ? io_r_67_b : _GEN_1766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1768 = 8'h44 == r_count_7_io_out ? io_r_68_b : _GEN_1767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1769 = 8'h45 == r_count_7_io_out ? io_r_69_b : _GEN_1768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1770 = 8'h46 == r_count_7_io_out ? io_r_70_b : _GEN_1769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1771 = 8'h47 == r_count_7_io_out ? io_r_71_b : _GEN_1770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1772 = 8'h48 == r_count_7_io_out ? io_r_72_b : _GEN_1771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1773 = 8'h49 == r_count_7_io_out ? io_r_73_b : _GEN_1772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1774 = 8'h4a == r_count_7_io_out ? io_r_74_b : _GEN_1773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1775 = 8'h4b == r_count_7_io_out ? io_r_75_b : _GEN_1774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1776 = 8'h4c == r_count_7_io_out ? io_r_76_b : _GEN_1775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1777 = 8'h4d == r_count_7_io_out ? io_r_77_b : _GEN_1776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1778 = 8'h4e == r_count_7_io_out ? io_r_78_b : _GEN_1777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1779 = 8'h4f == r_count_7_io_out ? io_r_79_b : _GEN_1778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1780 = 8'h50 == r_count_7_io_out ? io_r_80_b : _GEN_1779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1781 = 8'h51 == r_count_7_io_out ? io_r_81_b : _GEN_1780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1782 = 8'h52 == r_count_7_io_out ? io_r_82_b : _GEN_1781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1783 = 8'h53 == r_count_7_io_out ? io_r_83_b : _GEN_1782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1784 = 8'h54 == r_count_7_io_out ? io_r_84_b : _GEN_1783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1785 = 8'h55 == r_count_7_io_out ? io_r_85_b : _GEN_1784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1786 = 8'h56 == r_count_7_io_out ? io_r_86_b : _GEN_1785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1787 = 8'h57 == r_count_7_io_out ? io_r_87_b : _GEN_1786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1788 = 8'h58 == r_count_7_io_out ? io_r_88_b : _GEN_1787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1789 = 8'h59 == r_count_7_io_out ? io_r_89_b : _GEN_1788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1790 = 8'h5a == r_count_7_io_out ? io_r_90_b : _GEN_1789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1791 = 8'h5b == r_count_7_io_out ? io_r_91_b : _GEN_1790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1792 = 8'h5c == r_count_7_io_out ? io_r_92_b : _GEN_1791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1793 = 8'h5d == r_count_7_io_out ? io_r_93_b : _GEN_1792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1794 = 8'h5e == r_count_7_io_out ? io_r_94_b : _GEN_1793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1795 = 8'h5f == r_count_7_io_out ? io_r_95_b : _GEN_1794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1796 = 8'h60 == r_count_7_io_out ? io_r_96_b : _GEN_1795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1797 = 8'h61 == r_count_7_io_out ? io_r_97_b : _GEN_1796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1798 = 8'h62 == r_count_7_io_out ? io_r_98_b : _GEN_1797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1799 = 8'h63 == r_count_7_io_out ? io_r_99_b : _GEN_1798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1800 = 8'h64 == r_count_7_io_out ? io_r_100_b : _GEN_1799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1801 = 8'h65 == r_count_7_io_out ? io_r_101_b : _GEN_1800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1802 = 8'h66 == r_count_7_io_out ? io_r_102_b : _GEN_1801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1803 = 8'h67 == r_count_7_io_out ? io_r_103_b : _GEN_1802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1804 = 8'h68 == r_count_7_io_out ? io_r_104_b : _GEN_1803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1805 = 8'h69 == r_count_7_io_out ? io_r_105_b : _GEN_1804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1806 = 8'h6a == r_count_7_io_out ? io_r_106_b : _GEN_1805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1807 = 8'h6b == r_count_7_io_out ? io_r_107_b : _GEN_1806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1808 = 8'h6c == r_count_7_io_out ? io_r_108_b : _GEN_1807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1809 = 8'h6d == r_count_7_io_out ? io_r_109_b : _GEN_1808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1810 = 8'h6e == r_count_7_io_out ? io_r_110_b : _GEN_1809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1811 = 8'h6f == r_count_7_io_out ? io_r_111_b : _GEN_1810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1812 = 8'h70 == r_count_7_io_out ? io_r_112_b : _GEN_1811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1813 = 8'h71 == r_count_7_io_out ? io_r_113_b : _GEN_1812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1814 = 8'h72 == r_count_7_io_out ? io_r_114_b : _GEN_1813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1815 = 8'h73 == r_count_7_io_out ? io_r_115_b : _GEN_1814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1816 = 8'h74 == r_count_7_io_out ? io_r_116_b : _GEN_1815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1817 = 8'h75 == r_count_7_io_out ? io_r_117_b : _GEN_1816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1818 = 8'h76 == r_count_7_io_out ? io_r_118_b : _GEN_1817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1819 = 8'h77 == r_count_7_io_out ? io_r_119_b : _GEN_1818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1820 = 8'h78 == r_count_7_io_out ? io_r_120_b : _GEN_1819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1821 = 8'h79 == r_count_7_io_out ? io_r_121_b : _GEN_1820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1822 = 8'h7a == r_count_7_io_out ? io_r_122_b : _GEN_1821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1823 = 8'h7b == r_count_7_io_out ? io_r_123_b : _GEN_1822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1824 = 8'h7c == r_count_7_io_out ? io_r_124_b : _GEN_1823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1825 = 8'h7d == r_count_7_io_out ? io_r_125_b : _GEN_1824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1826 = 8'h7e == r_count_7_io_out ? io_r_126_b : _GEN_1825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1827 = 8'h7f == r_count_7_io_out ? io_r_127_b : _GEN_1826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1828 = 8'h80 == r_count_7_io_out ? io_r_128_b : _GEN_1827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1829 = 8'h81 == r_count_7_io_out ? io_r_129_b : _GEN_1828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1830 = 8'h82 == r_count_7_io_out ? io_r_130_b : _GEN_1829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1831 = 8'h83 == r_count_7_io_out ? io_r_131_b : _GEN_1830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1832 = 8'h84 == r_count_7_io_out ? io_r_132_b : _GEN_1831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1833 = 8'h85 == r_count_7_io_out ? io_r_133_b : _GEN_1832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1834 = 8'h86 == r_count_7_io_out ? io_r_134_b : _GEN_1833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1835 = 8'h87 == r_count_7_io_out ? io_r_135_b : _GEN_1834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1836 = 8'h88 == r_count_7_io_out ? io_r_136_b : _GEN_1835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1837 = 8'h89 == r_count_7_io_out ? io_r_137_b : _GEN_1836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1838 = 8'h8a == r_count_7_io_out ? io_r_138_b : _GEN_1837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1839 = 8'h8b == r_count_7_io_out ? io_r_139_b : _GEN_1838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1840 = 8'h8c == r_count_7_io_out ? io_r_140_b : _GEN_1839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1841 = 8'h8d == r_count_7_io_out ? io_r_141_b : _GEN_1840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1842 = 8'h8e == r_count_7_io_out ? io_r_142_b : _GEN_1841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1843 = 8'h8f == r_count_7_io_out ? io_r_143_b : _GEN_1842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1844 = 8'h90 == r_count_7_io_out ? io_r_144_b : _GEN_1843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1845 = 8'h91 == r_count_7_io_out ? io_r_145_b : _GEN_1844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1846 = 8'h92 == r_count_7_io_out ? io_r_146_b : _GEN_1845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1847 = 8'h93 == r_count_7_io_out ? io_r_147_b : _GEN_1846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1848 = 8'h94 == r_count_7_io_out ? io_r_148_b : _GEN_1847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1849 = 8'h95 == r_count_7_io_out ? io_r_149_b : _GEN_1848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1850 = 8'h96 == r_count_7_io_out ? io_r_150_b : _GEN_1849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1851 = 8'h97 == r_count_7_io_out ? io_r_151_b : _GEN_1850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1852 = 8'h98 == r_count_7_io_out ? io_r_152_b : _GEN_1851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1853 = 8'h99 == r_count_7_io_out ? io_r_153_b : _GEN_1852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1854 = 8'h9a == r_count_7_io_out ? io_r_154_b : _GEN_1853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1855 = 8'h9b == r_count_7_io_out ? io_r_155_b : _GEN_1854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1856 = 8'h9c == r_count_7_io_out ? io_r_156_b : _GEN_1855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1857 = 8'h9d == r_count_7_io_out ? io_r_157_b : _GEN_1856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1858 = 8'h9e == r_count_7_io_out ? io_r_158_b : _GEN_1857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1859 = 8'h9f == r_count_7_io_out ? io_r_159_b : _GEN_1858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1860 = 8'ha0 == r_count_7_io_out ? io_r_160_b : _GEN_1859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1861 = 8'ha1 == r_count_7_io_out ? io_r_161_b : _GEN_1860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1862 = 8'ha2 == r_count_7_io_out ? io_r_162_b : _GEN_1861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1863 = 8'ha3 == r_count_7_io_out ? io_r_163_b : _GEN_1862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1864 = 8'ha4 == r_count_7_io_out ? io_r_164_b : _GEN_1863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1865 = 8'ha5 == r_count_7_io_out ? io_r_165_b : _GEN_1864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1866 = 8'ha6 == r_count_7_io_out ? io_r_166_b : _GEN_1865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1867 = 8'ha7 == r_count_7_io_out ? io_r_167_b : _GEN_1866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1868 = 8'ha8 == r_count_7_io_out ? io_r_168_b : _GEN_1867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1869 = 8'ha9 == r_count_7_io_out ? io_r_169_b : _GEN_1868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1870 = 8'haa == r_count_7_io_out ? io_r_170_b : _GEN_1869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1871 = 8'hab == r_count_7_io_out ? io_r_171_b : _GEN_1870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1872 = 8'hac == r_count_7_io_out ? io_r_172_b : _GEN_1871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1873 = 8'had == r_count_7_io_out ? io_r_173_b : _GEN_1872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1874 = 8'hae == r_count_7_io_out ? io_r_174_b : _GEN_1873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1875 = 8'haf == r_count_7_io_out ? io_r_175_b : _GEN_1874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1876 = 8'hb0 == r_count_7_io_out ? io_r_176_b : _GEN_1875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1877 = 8'hb1 == r_count_7_io_out ? io_r_177_b : _GEN_1876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1878 = 8'hb2 == r_count_7_io_out ? io_r_178_b : _GEN_1877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1879 = 8'hb3 == r_count_7_io_out ? io_r_179_b : _GEN_1878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1880 = 8'hb4 == r_count_7_io_out ? io_r_180_b : _GEN_1879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1881 = 8'hb5 == r_count_7_io_out ? io_r_181_b : _GEN_1880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1882 = 8'hb6 == r_count_7_io_out ? io_r_182_b : _GEN_1881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1883 = 8'hb7 == r_count_7_io_out ? io_r_183_b : _GEN_1882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1884 = 8'hb8 == r_count_7_io_out ? io_r_184_b : _GEN_1883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1885 = 8'hb9 == r_count_7_io_out ? io_r_185_b : _GEN_1884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1886 = 8'hba == r_count_7_io_out ? io_r_186_b : _GEN_1885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1887 = 8'hbb == r_count_7_io_out ? io_r_187_b : _GEN_1886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1888 = 8'hbc == r_count_7_io_out ? io_r_188_b : _GEN_1887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1889 = 8'hbd == r_count_7_io_out ? io_r_189_b : _GEN_1888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1890 = 8'hbe == r_count_7_io_out ? io_r_190_b : _GEN_1889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1891 = 8'hbf == r_count_7_io_out ? io_r_191_b : _GEN_1890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1892 = 8'hc0 == r_count_7_io_out ? io_r_192_b : _GEN_1891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1893 = 8'hc1 == r_count_7_io_out ? io_r_193_b : _GEN_1892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1894 = 8'hc2 == r_count_7_io_out ? io_r_194_b : _GEN_1893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1895 = 8'hc3 == r_count_7_io_out ? io_r_195_b : _GEN_1894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1896 = 8'hc4 == r_count_7_io_out ? io_r_196_b : _GEN_1895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1897 = 8'hc5 == r_count_7_io_out ? io_r_197_b : _GEN_1896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1898 = 8'hc6 == r_count_7_io_out ? io_r_198_b : _GEN_1897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1901 = 8'h1 == r_count_8_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1902 = 8'h2 == r_count_8_io_out ? io_r_2_b : _GEN_1901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1903 = 8'h3 == r_count_8_io_out ? io_r_3_b : _GEN_1902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1904 = 8'h4 == r_count_8_io_out ? io_r_4_b : _GEN_1903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1905 = 8'h5 == r_count_8_io_out ? io_r_5_b : _GEN_1904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1906 = 8'h6 == r_count_8_io_out ? io_r_6_b : _GEN_1905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1907 = 8'h7 == r_count_8_io_out ? io_r_7_b : _GEN_1906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1908 = 8'h8 == r_count_8_io_out ? io_r_8_b : _GEN_1907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1909 = 8'h9 == r_count_8_io_out ? io_r_9_b : _GEN_1908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1910 = 8'ha == r_count_8_io_out ? io_r_10_b : _GEN_1909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1911 = 8'hb == r_count_8_io_out ? io_r_11_b : _GEN_1910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1912 = 8'hc == r_count_8_io_out ? io_r_12_b : _GEN_1911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1913 = 8'hd == r_count_8_io_out ? io_r_13_b : _GEN_1912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1914 = 8'he == r_count_8_io_out ? io_r_14_b : _GEN_1913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1915 = 8'hf == r_count_8_io_out ? io_r_15_b : _GEN_1914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1916 = 8'h10 == r_count_8_io_out ? io_r_16_b : _GEN_1915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1917 = 8'h11 == r_count_8_io_out ? io_r_17_b : _GEN_1916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1918 = 8'h12 == r_count_8_io_out ? io_r_18_b : _GEN_1917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1919 = 8'h13 == r_count_8_io_out ? io_r_19_b : _GEN_1918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1920 = 8'h14 == r_count_8_io_out ? io_r_20_b : _GEN_1919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1921 = 8'h15 == r_count_8_io_out ? io_r_21_b : _GEN_1920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1922 = 8'h16 == r_count_8_io_out ? io_r_22_b : _GEN_1921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1923 = 8'h17 == r_count_8_io_out ? io_r_23_b : _GEN_1922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1924 = 8'h18 == r_count_8_io_out ? io_r_24_b : _GEN_1923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1925 = 8'h19 == r_count_8_io_out ? io_r_25_b : _GEN_1924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1926 = 8'h1a == r_count_8_io_out ? io_r_26_b : _GEN_1925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1927 = 8'h1b == r_count_8_io_out ? io_r_27_b : _GEN_1926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1928 = 8'h1c == r_count_8_io_out ? io_r_28_b : _GEN_1927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1929 = 8'h1d == r_count_8_io_out ? io_r_29_b : _GEN_1928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1930 = 8'h1e == r_count_8_io_out ? io_r_30_b : _GEN_1929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1931 = 8'h1f == r_count_8_io_out ? io_r_31_b : _GEN_1930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1932 = 8'h20 == r_count_8_io_out ? io_r_32_b : _GEN_1931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1933 = 8'h21 == r_count_8_io_out ? io_r_33_b : _GEN_1932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1934 = 8'h22 == r_count_8_io_out ? io_r_34_b : _GEN_1933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1935 = 8'h23 == r_count_8_io_out ? io_r_35_b : _GEN_1934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1936 = 8'h24 == r_count_8_io_out ? io_r_36_b : _GEN_1935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1937 = 8'h25 == r_count_8_io_out ? io_r_37_b : _GEN_1936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1938 = 8'h26 == r_count_8_io_out ? io_r_38_b : _GEN_1937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1939 = 8'h27 == r_count_8_io_out ? io_r_39_b : _GEN_1938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1940 = 8'h28 == r_count_8_io_out ? io_r_40_b : _GEN_1939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1941 = 8'h29 == r_count_8_io_out ? io_r_41_b : _GEN_1940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1942 = 8'h2a == r_count_8_io_out ? io_r_42_b : _GEN_1941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1943 = 8'h2b == r_count_8_io_out ? io_r_43_b : _GEN_1942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1944 = 8'h2c == r_count_8_io_out ? io_r_44_b : _GEN_1943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1945 = 8'h2d == r_count_8_io_out ? io_r_45_b : _GEN_1944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1946 = 8'h2e == r_count_8_io_out ? io_r_46_b : _GEN_1945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1947 = 8'h2f == r_count_8_io_out ? io_r_47_b : _GEN_1946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1948 = 8'h30 == r_count_8_io_out ? io_r_48_b : _GEN_1947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1949 = 8'h31 == r_count_8_io_out ? io_r_49_b : _GEN_1948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1950 = 8'h32 == r_count_8_io_out ? io_r_50_b : _GEN_1949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1951 = 8'h33 == r_count_8_io_out ? io_r_51_b : _GEN_1950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1952 = 8'h34 == r_count_8_io_out ? io_r_52_b : _GEN_1951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1953 = 8'h35 == r_count_8_io_out ? io_r_53_b : _GEN_1952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1954 = 8'h36 == r_count_8_io_out ? io_r_54_b : _GEN_1953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1955 = 8'h37 == r_count_8_io_out ? io_r_55_b : _GEN_1954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1956 = 8'h38 == r_count_8_io_out ? io_r_56_b : _GEN_1955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1957 = 8'h39 == r_count_8_io_out ? io_r_57_b : _GEN_1956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1958 = 8'h3a == r_count_8_io_out ? io_r_58_b : _GEN_1957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1959 = 8'h3b == r_count_8_io_out ? io_r_59_b : _GEN_1958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1960 = 8'h3c == r_count_8_io_out ? io_r_60_b : _GEN_1959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1961 = 8'h3d == r_count_8_io_out ? io_r_61_b : _GEN_1960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1962 = 8'h3e == r_count_8_io_out ? io_r_62_b : _GEN_1961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1963 = 8'h3f == r_count_8_io_out ? io_r_63_b : _GEN_1962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1964 = 8'h40 == r_count_8_io_out ? io_r_64_b : _GEN_1963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1965 = 8'h41 == r_count_8_io_out ? io_r_65_b : _GEN_1964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1966 = 8'h42 == r_count_8_io_out ? io_r_66_b : _GEN_1965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1967 = 8'h43 == r_count_8_io_out ? io_r_67_b : _GEN_1966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1968 = 8'h44 == r_count_8_io_out ? io_r_68_b : _GEN_1967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1969 = 8'h45 == r_count_8_io_out ? io_r_69_b : _GEN_1968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1970 = 8'h46 == r_count_8_io_out ? io_r_70_b : _GEN_1969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1971 = 8'h47 == r_count_8_io_out ? io_r_71_b : _GEN_1970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1972 = 8'h48 == r_count_8_io_out ? io_r_72_b : _GEN_1971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1973 = 8'h49 == r_count_8_io_out ? io_r_73_b : _GEN_1972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1974 = 8'h4a == r_count_8_io_out ? io_r_74_b : _GEN_1973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1975 = 8'h4b == r_count_8_io_out ? io_r_75_b : _GEN_1974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1976 = 8'h4c == r_count_8_io_out ? io_r_76_b : _GEN_1975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1977 = 8'h4d == r_count_8_io_out ? io_r_77_b : _GEN_1976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1978 = 8'h4e == r_count_8_io_out ? io_r_78_b : _GEN_1977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1979 = 8'h4f == r_count_8_io_out ? io_r_79_b : _GEN_1978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1980 = 8'h50 == r_count_8_io_out ? io_r_80_b : _GEN_1979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1981 = 8'h51 == r_count_8_io_out ? io_r_81_b : _GEN_1980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1982 = 8'h52 == r_count_8_io_out ? io_r_82_b : _GEN_1981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1983 = 8'h53 == r_count_8_io_out ? io_r_83_b : _GEN_1982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1984 = 8'h54 == r_count_8_io_out ? io_r_84_b : _GEN_1983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1985 = 8'h55 == r_count_8_io_out ? io_r_85_b : _GEN_1984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1986 = 8'h56 == r_count_8_io_out ? io_r_86_b : _GEN_1985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1987 = 8'h57 == r_count_8_io_out ? io_r_87_b : _GEN_1986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1988 = 8'h58 == r_count_8_io_out ? io_r_88_b : _GEN_1987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1989 = 8'h59 == r_count_8_io_out ? io_r_89_b : _GEN_1988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1990 = 8'h5a == r_count_8_io_out ? io_r_90_b : _GEN_1989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1991 = 8'h5b == r_count_8_io_out ? io_r_91_b : _GEN_1990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1992 = 8'h5c == r_count_8_io_out ? io_r_92_b : _GEN_1991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1993 = 8'h5d == r_count_8_io_out ? io_r_93_b : _GEN_1992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1994 = 8'h5e == r_count_8_io_out ? io_r_94_b : _GEN_1993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1995 = 8'h5f == r_count_8_io_out ? io_r_95_b : _GEN_1994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1996 = 8'h60 == r_count_8_io_out ? io_r_96_b : _GEN_1995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1997 = 8'h61 == r_count_8_io_out ? io_r_97_b : _GEN_1996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1998 = 8'h62 == r_count_8_io_out ? io_r_98_b : _GEN_1997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1999 = 8'h63 == r_count_8_io_out ? io_r_99_b : _GEN_1998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2000 = 8'h64 == r_count_8_io_out ? io_r_100_b : _GEN_1999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2001 = 8'h65 == r_count_8_io_out ? io_r_101_b : _GEN_2000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2002 = 8'h66 == r_count_8_io_out ? io_r_102_b : _GEN_2001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2003 = 8'h67 == r_count_8_io_out ? io_r_103_b : _GEN_2002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2004 = 8'h68 == r_count_8_io_out ? io_r_104_b : _GEN_2003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2005 = 8'h69 == r_count_8_io_out ? io_r_105_b : _GEN_2004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2006 = 8'h6a == r_count_8_io_out ? io_r_106_b : _GEN_2005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2007 = 8'h6b == r_count_8_io_out ? io_r_107_b : _GEN_2006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2008 = 8'h6c == r_count_8_io_out ? io_r_108_b : _GEN_2007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2009 = 8'h6d == r_count_8_io_out ? io_r_109_b : _GEN_2008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2010 = 8'h6e == r_count_8_io_out ? io_r_110_b : _GEN_2009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2011 = 8'h6f == r_count_8_io_out ? io_r_111_b : _GEN_2010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2012 = 8'h70 == r_count_8_io_out ? io_r_112_b : _GEN_2011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2013 = 8'h71 == r_count_8_io_out ? io_r_113_b : _GEN_2012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2014 = 8'h72 == r_count_8_io_out ? io_r_114_b : _GEN_2013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2015 = 8'h73 == r_count_8_io_out ? io_r_115_b : _GEN_2014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2016 = 8'h74 == r_count_8_io_out ? io_r_116_b : _GEN_2015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2017 = 8'h75 == r_count_8_io_out ? io_r_117_b : _GEN_2016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2018 = 8'h76 == r_count_8_io_out ? io_r_118_b : _GEN_2017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2019 = 8'h77 == r_count_8_io_out ? io_r_119_b : _GEN_2018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2020 = 8'h78 == r_count_8_io_out ? io_r_120_b : _GEN_2019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2021 = 8'h79 == r_count_8_io_out ? io_r_121_b : _GEN_2020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2022 = 8'h7a == r_count_8_io_out ? io_r_122_b : _GEN_2021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2023 = 8'h7b == r_count_8_io_out ? io_r_123_b : _GEN_2022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2024 = 8'h7c == r_count_8_io_out ? io_r_124_b : _GEN_2023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2025 = 8'h7d == r_count_8_io_out ? io_r_125_b : _GEN_2024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2026 = 8'h7e == r_count_8_io_out ? io_r_126_b : _GEN_2025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2027 = 8'h7f == r_count_8_io_out ? io_r_127_b : _GEN_2026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2028 = 8'h80 == r_count_8_io_out ? io_r_128_b : _GEN_2027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2029 = 8'h81 == r_count_8_io_out ? io_r_129_b : _GEN_2028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2030 = 8'h82 == r_count_8_io_out ? io_r_130_b : _GEN_2029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2031 = 8'h83 == r_count_8_io_out ? io_r_131_b : _GEN_2030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2032 = 8'h84 == r_count_8_io_out ? io_r_132_b : _GEN_2031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2033 = 8'h85 == r_count_8_io_out ? io_r_133_b : _GEN_2032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2034 = 8'h86 == r_count_8_io_out ? io_r_134_b : _GEN_2033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2035 = 8'h87 == r_count_8_io_out ? io_r_135_b : _GEN_2034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2036 = 8'h88 == r_count_8_io_out ? io_r_136_b : _GEN_2035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2037 = 8'h89 == r_count_8_io_out ? io_r_137_b : _GEN_2036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2038 = 8'h8a == r_count_8_io_out ? io_r_138_b : _GEN_2037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2039 = 8'h8b == r_count_8_io_out ? io_r_139_b : _GEN_2038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2040 = 8'h8c == r_count_8_io_out ? io_r_140_b : _GEN_2039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2041 = 8'h8d == r_count_8_io_out ? io_r_141_b : _GEN_2040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2042 = 8'h8e == r_count_8_io_out ? io_r_142_b : _GEN_2041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2043 = 8'h8f == r_count_8_io_out ? io_r_143_b : _GEN_2042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2044 = 8'h90 == r_count_8_io_out ? io_r_144_b : _GEN_2043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2045 = 8'h91 == r_count_8_io_out ? io_r_145_b : _GEN_2044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2046 = 8'h92 == r_count_8_io_out ? io_r_146_b : _GEN_2045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2047 = 8'h93 == r_count_8_io_out ? io_r_147_b : _GEN_2046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2048 = 8'h94 == r_count_8_io_out ? io_r_148_b : _GEN_2047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2049 = 8'h95 == r_count_8_io_out ? io_r_149_b : _GEN_2048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2050 = 8'h96 == r_count_8_io_out ? io_r_150_b : _GEN_2049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2051 = 8'h97 == r_count_8_io_out ? io_r_151_b : _GEN_2050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2052 = 8'h98 == r_count_8_io_out ? io_r_152_b : _GEN_2051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2053 = 8'h99 == r_count_8_io_out ? io_r_153_b : _GEN_2052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2054 = 8'h9a == r_count_8_io_out ? io_r_154_b : _GEN_2053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2055 = 8'h9b == r_count_8_io_out ? io_r_155_b : _GEN_2054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2056 = 8'h9c == r_count_8_io_out ? io_r_156_b : _GEN_2055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2057 = 8'h9d == r_count_8_io_out ? io_r_157_b : _GEN_2056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2058 = 8'h9e == r_count_8_io_out ? io_r_158_b : _GEN_2057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2059 = 8'h9f == r_count_8_io_out ? io_r_159_b : _GEN_2058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2060 = 8'ha0 == r_count_8_io_out ? io_r_160_b : _GEN_2059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2061 = 8'ha1 == r_count_8_io_out ? io_r_161_b : _GEN_2060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2062 = 8'ha2 == r_count_8_io_out ? io_r_162_b : _GEN_2061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2063 = 8'ha3 == r_count_8_io_out ? io_r_163_b : _GEN_2062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2064 = 8'ha4 == r_count_8_io_out ? io_r_164_b : _GEN_2063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2065 = 8'ha5 == r_count_8_io_out ? io_r_165_b : _GEN_2064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2066 = 8'ha6 == r_count_8_io_out ? io_r_166_b : _GEN_2065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2067 = 8'ha7 == r_count_8_io_out ? io_r_167_b : _GEN_2066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2068 = 8'ha8 == r_count_8_io_out ? io_r_168_b : _GEN_2067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2069 = 8'ha9 == r_count_8_io_out ? io_r_169_b : _GEN_2068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2070 = 8'haa == r_count_8_io_out ? io_r_170_b : _GEN_2069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2071 = 8'hab == r_count_8_io_out ? io_r_171_b : _GEN_2070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2072 = 8'hac == r_count_8_io_out ? io_r_172_b : _GEN_2071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2073 = 8'had == r_count_8_io_out ? io_r_173_b : _GEN_2072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2074 = 8'hae == r_count_8_io_out ? io_r_174_b : _GEN_2073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2075 = 8'haf == r_count_8_io_out ? io_r_175_b : _GEN_2074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2076 = 8'hb0 == r_count_8_io_out ? io_r_176_b : _GEN_2075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2077 = 8'hb1 == r_count_8_io_out ? io_r_177_b : _GEN_2076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2078 = 8'hb2 == r_count_8_io_out ? io_r_178_b : _GEN_2077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2079 = 8'hb3 == r_count_8_io_out ? io_r_179_b : _GEN_2078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2080 = 8'hb4 == r_count_8_io_out ? io_r_180_b : _GEN_2079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2081 = 8'hb5 == r_count_8_io_out ? io_r_181_b : _GEN_2080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2082 = 8'hb6 == r_count_8_io_out ? io_r_182_b : _GEN_2081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2083 = 8'hb7 == r_count_8_io_out ? io_r_183_b : _GEN_2082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2084 = 8'hb8 == r_count_8_io_out ? io_r_184_b : _GEN_2083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2085 = 8'hb9 == r_count_8_io_out ? io_r_185_b : _GEN_2084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2086 = 8'hba == r_count_8_io_out ? io_r_186_b : _GEN_2085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2087 = 8'hbb == r_count_8_io_out ? io_r_187_b : _GEN_2086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2088 = 8'hbc == r_count_8_io_out ? io_r_188_b : _GEN_2087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2089 = 8'hbd == r_count_8_io_out ? io_r_189_b : _GEN_2088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2090 = 8'hbe == r_count_8_io_out ? io_r_190_b : _GEN_2089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2091 = 8'hbf == r_count_8_io_out ? io_r_191_b : _GEN_2090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2092 = 8'hc0 == r_count_8_io_out ? io_r_192_b : _GEN_2091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2093 = 8'hc1 == r_count_8_io_out ? io_r_193_b : _GEN_2092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2094 = 8'hc2 == r_count_8_io_out ? io_r_194_b : _GEN_2093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2095 = 8'hc3 == r_count_8_io_out ? io_r_195_b : _GEN_2094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2096 = 8'hc4 == r_count_8_io_out ? io_r_196_b : _GEN_2095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2097 = 8'hc5 == r_count_8_io_out ? io_r_197_b : _GEN_2096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2098 = 8'hc6 == r_count_8_io_out ? io_r_198_b : _GEN_2097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2101 = 8'h1 == r_count_9_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2102 = 8'h2 == r_count_9_io_out ? io_r_2_b : _GEN_2101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2103 = 8'h3 == r_count_9_io_out ? io_r_3_b : _GEN_2102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2104 = 8'h4 == r_count_9_io_out ? io_r_4_b : _GEN_2103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2105 = 8'h5 == r_count_9_io_out ? io_r_5_b : _GEN_2104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2106 = 8'h6 == r_count_9_io_out ? io_r_6_b : _GEN_2105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2107 = 8'h7 == r_count_9_io_out ? io_r_7_b : _GEN_2106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2108 = 8'h8 == r_count_9_io_out ? io_r_8_b : _GEN_2107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2109 = 8'h9 == r_count_9_io_out ? io_r_9_b : _GEN_2108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2110 = 8'ha == r_count_9_io_out ? io_r_10_b : _GEN_2109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2111 = 8'hb == r_count_9_io_out ? io_r_11_b : _GEN_2110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2112 = 8'hc == r_count_9_io_out ? io_r_12_b : _GEN_2111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2113 = 8'hd == r_count_9_io_out ? io_r_13_b : _GEN_2112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2114 = 8'he == r_count_9_io_out ? io_r_14_b : _GEN_2113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2115 = 8'hf == r_count_9_io_out ? io_r_15_b : _GEN_2114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2116 = 8'h10 == r_count_9_io_out ? io_r_16_b : _GEN_2115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2117 = 8'h11 == r_count_9_io_out ? io_r_17_b : _GEN_2116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2118 = 8'h12 == r_count_9_io_out ? io_r_18_b : _GEN_2117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2119 = 8'h13 == r_count_9_io_out ? io_r_19_b : _GEN_2118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2120 = 8'h14 == r_count_9_io_out ? io_r_20_b : _GEN_2119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2121 = 8'h15 == r_count_9_io_out ? io_r_21_b : _GEN_2120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2122 = 8'h16 == r_count_9_io_out ? io_r_22_b : _GEN_2121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2123 = 8'h17 == r_count_9_io_out ? io_r_23_b : _GEN_2122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2124 = 8'h18 == r_count_9_io_out ? io_r_24_b : _GEN_2123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2125 = 8'h19 == r_count_9_io_out ? io_r_25_b : _GEN_2124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2126 = 8'h1a == r_count_9_io_out ? io_r_26_b : _GEN_2125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2127 = 8'h1b == r_count_9_io_out ? io_r_27_b : _GEN_2126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2128 = 8'h1c == r_count_9_io_out ? io_r_28_b : _GEN_2127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2129 = 8'h1d == r_count_9_io_out ? io_r_29_b : _GEN_2128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2130 = 8'h1e == r_count_9_io_out ? io_r_30_b : _GEN_2129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2131 = 8'h1f == r_count_9_io_out ? io_r_31_b : _GEN_2130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2132 = 8'h20 == r_count_9_io_out ? io_r_32_b : _GEN_2131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2133 = 8'h21 == r_count_9_io_out ? io_r_33_b : _GEN_2132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2134 = 8'h22 == r_count_9_io_out ? io_r_34_b : _GEN_2133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2135 = 8'h23 == r_count_9_io_out ? io_r_35_b : _GEN_2134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2136 = 8'h24 == r_count_9_io_out ? io_r_36_b : _GEN_2135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2137 = 8'h25 == r_count_9_io_out ? io_r_37_b : _GEN_2136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2138 = 8'h26 == r_count_9_io_out ? io_r_38_b : _GEN_2137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2139 = 8'h27 == r_count_9_io_out ? io_r_39_b : _GEN_2138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2140 = 8'h28 == r_count_9_io_out ? io_r_40_b : _GEN_2139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2141 = 8'h29 == r_count_9_io_out ? io_r_41_b : _GEN_2140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2142 = 8'h2a == r_count_9_io_out ? io_r_42_b : _GEN_2141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2143 = 8'h2b == r_count_9_io_out ? io_r_43_b : _GEN_2142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2144 = 8'h2c == r_count_9_io_out ? io_r_44_b : _GEN_2143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2145 = 8'h2d == r_count_9_io_out ? io_r_45_b : _GEN_2144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2146 = 8'h2e == r_count_9_io_out ? io_r_46_b : _GEN_2145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2147 = 8'h2f == r_count_9_io_out ? io_r_47_b : _GEN_2146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2148 = 8'h30 == r_count_9_io_out ? io_r_48_b : _GEN_2147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2149 = 8'h31 == r_count_9_io_out ? io_r_49_b : _GEN_2148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2150 = 8'h32 == r_count_9_io_out ? io_r_50_b : _GEN_2149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2151 = 8'h33 == r_count_9_io_out ? io_r_51_b : _GEN_2150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2152 = 8'h34 == r_count_9_io_out ? io_r_52_b : _GEN_2151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2153 = 8'h35 == r_count_9_io_out ? io_r_53_b : _GEN_2152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2154 = 8'h36 == r_count_9_io_out ? io_r_54_b : _GEN_2153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2155 = 8'h37 == r_count_9_io_out ? io_r_55_b : _GEN_2154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2156 = 8'h38 == r_count_9_io_out ? io_r_56_b : _GEN_2155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2157 = 8'h39 == r_count_9_io_out ? io_r_57_b : _GEN_2156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2158 = 8'h3a == r_count_9_io_out ? io_r_58_b : _GEN_2157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2159 = 8'h3b == r_count_9_io_out ? io_r_59_b : _GEN_2158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2160 = 8'h3c == r_count_9_io_out ? io_r_60_b : _GEN_2159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2161 = 8'h3d == r_count_9_io_out ? io_r_61_b : _GEN_2160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2162 = 8'h3e == r_count_9_io_out ? io_r_62_b : _GEN_2161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2163 = 8'h3f == r_count_9_io_out ? io_r_63_b : _GEN_2162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2164 = 8'h40 == r_count_9_io_out ? io_r_64_b : _GEN_2163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2165 = 8'h41 == r_count_9_io_out ? io_r_65_b : _GEN_2164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2166 = 8'h42 == r_count_9_io_out ? io_r_66_b : _GEN_2165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2167 = 8'h43 == r_count_9_io_out ? io_r_67_b : _GEN_2166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2168 = 8'h44 == r_count_9_io_out ? io_r_68_b : _GEN_2167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2169 = 8'h45 == r_count_9_io_out ? io_r_69_b : _GEN_2168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2170 = 8'h46 == r_count_9_io_out ? io_r_70_b : _GEN_2169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2171 = 8'h47 == r_count_9_io_out ? io_r_71_b : _GEN_2170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2172 = 8'h48 == r_count_9_io_out ? io_r_72_b : _GEN_2171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2173 = 8'h49 == r_count_9_io_out ? io_r_73_b : _GEN_2172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2174 = 8'h4a == r_count_9_io_out ? io_r_74_b : _GEN_2173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2175 = 8'h4b == r_count_9_io_out ? io_r_75_b : _GEN_2174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2176 = 8'h4c == r_count_9_io_out ? io_r_76_b : _GEN_2175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2177 = 8'h4d == r_count_9_io_out ? io_r_77_b : _GEN_2176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2178 = 8'h4e == r_count_9_io_out ? io_r_78_b : _GEN_2177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2179 = 8'h4f == r_count_9_io_out ? io_r_79_b : _GEN_2178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2180 = 8'h50 == r_count_9_io_out ? io_r_80_b : _GEN_2179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2181 = 8'h51 == r_count_9_io_out ? io_r_81_b : _GEN_2180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2182 = 8'h52 == r_count_9_io_out ? io_r_82_b : _GEN_2181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2183 = 8'h53 == r_count_9_io_out ? io_r_83_b : _GEN_2182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2184 = 8'h54 == r_count_9_io_out ? io_r_84_b : _GEN_2183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2185 = 8'h55 == r_count_9_io_out ? io_r_85_b : _GEN_2184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2186 = 8'h56 == r_count_9_io_out ? io_r_86_b : _GEN_2185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2187 = 8'h57 == r_count_9_io_out ? io_r_87_b : _GEN_2186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2188 = 8'h58 == r_count_9_io_out ? io_r_88_b : _GEN_2187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2189 = 8'h59 == r_count_9_io_out ? io_r_89_b : _GEN_2188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2190 = 8'h5a == r_count_9_io_out ? io_r_90_b : _GEN_2189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2191 = 8'h5b == r_count_9_io_out ? io_r_91_b : _GEN_2190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2192 = 8'h5c == r_count_9_io_out ? io_r_92_b : _GEN_2191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2193 = 8'h5d == r_count_9_io_out ? io_r_93_b : _GEN_2192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2194 = 8'h5e == r_count_9_io_out ? io_r_94_b : _GEN_2193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2195 = 8'h5f == r_count_9_io_out ? io_r_95_b : _GEN_2194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2196 = 8'h60 == r_count_9_io_out ? io_r_96_b : _GEN_2195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2197 = 8'h61 == r_count_9_io_out ? io_r_97_b : _GEN_2196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2198 = 8'h62 == r_count_9_io_out ? io_r_98_b : _GEN_2197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2199 = 8'h63 == r_count_9_io_out ? io_r_99_b : _GEN_2198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2200 = 8'h64 == r_count_9_io_out ? io_r_100_b : _GEN_2199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2201 = 8'h65 == r_count_9_io_out ? io_r_101_b : _GEN_2200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2202 = 8'h66 == r_count_9_io_out ? io_r_102_b : _GEN_2201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2203 = 8'h67 == r_count_9_io_out ? io_r_103_b : _GEN_2202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2204 = 8'h68 == r_count_9_io_out ? io_r_104_b : _GEN_2203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2205 = 8'h69 == r_count_9_io_out ? io_r_105_b : _GEN_2204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2206 = 8'h6a == r_count_9_io_out ? io_r_106_b : _GEN_2205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2207 = 8'h6b == r_count_9_io_out ? io_r_107_b : _GEN_2206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2208 = 8'h6c == r_count_9_io_out ? io_r_108_b : _GEN_2207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2209 = 8'h6d == r_count_9_io_out ? io_r_109_b : _GEN_2208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2210 = 8'h6e == r_count_9_io_out ? io_r_110_b : _GEN_2209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2211 = 8'h6f == r_count_9_io_out ? io_r_111_b : _GEN_2210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2212 = 8'h70 == r_count_9_io_out ? io_r_112_b : _GEN_2211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2213 = 8'h71 == r_count_9_io_out ? io_r_113_b : _GEN_2212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2214 = 8'h72 == r_count_9_io_out ? io_r_114_b : _GEN_2213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2215 = 8'h73 == r_count_9_io_out ? io_r_115_b : _GEN_2214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2216 = 8'h74 == r_count_9_io_out ? io_r_116_b : _GEN_2215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2217 = 8'h75 == r_count_9_io_out ? io_r_117_b : _GEN_2216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2218 = 8'h76 == r_count_9_io_out ? io_r_118_b : _GEN_2217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2219 = 8'h77 == r_count_9_io_out ? io_r_119_b : _GEN_2218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2220 = 8'h78 == r_count_9_io_out ? io_r_120_b : _GEN_2219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2221 = 8'h79 == r_count_9_io_out ? io_r_121_b : _GEN_2220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2222 = 8'h7a == r_count_9_io_out ? io_r_122_b : _GEN_2221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2223 = 8'h7b == r_count_9_io_out ? io_r_123_b : _GEN_2222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2224 = 8'h7c == r_count_9_io_out ? io_r_124_b : _GEN_2223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2225 = 8'h7d == r_count_9_io_out ? io_r_125_b : _GEN_2224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2226 = 8'h7e == r_count_9_io_out ? io_r_126_b : _GEN_2225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2227 = 8'h7f == r_count_9_io_out ? io_r_127_b : _GEN_2226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2228 = 8'h80 == r_count_9_io_out ? io_r_128_b : _GEN_2227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2229 = 8'h81 == r_count_9_io_out ? io_r_129_b : _GEN_2228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2230 = 8'h82 == r_count_9_io_out ? io_r_130_b : _GEN_2229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2231 = 8'h83 == r_count_9_io_out ? io_r_131_b : _GEN_2230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2232 = 8'h84 == r_count_9_io_out ? io_r_132_b : _GEN_2231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2233 = 8'h85 == r_count_9_io_out ? io_r_133_b : _GEN_2232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2234 = 8'h86 == r_count_9_io_out ? io_r_134_b : _GEN_2233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2235 = 8'h87 == r_count_9_io_out ? io_r_135_b : _GEN_2234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2236 = 8'h88 == r_count_9_io_out ? io_r_136_b : _GEN_2235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2237 = 8'h89 == r_count_9_io_out ? io_r_137_b : _GEN_2236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2238 = 8'h8a == r_count_9_io_out ? io_r_138_b : _GEN_2237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2239 = 8'h8b == r_count_9_io_out ? io_r_139_b : _GEN_2238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2240 = 8'h8c == r_count_9_io_out ? io_r_140_b : _GEN_2239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2241 = 8'h8d == r_count_9_io_out ? io_r_141_b : _GEN_2240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2242 = 8'h8e == r_count_9_io_out ? io_r_142_b : _GEN_2241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2243 = 8'h8f == r_count_9_io_out ? io_r_143_b : _GEN_2242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2244 = 8'h90 == r_count_9_io_out ? io_r_144_b : _GEN_2243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2245 = 8'h91 == r_count_9_io_out ? io_r_145_b : _GEN_2244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2246 = 8'h92 == r_count_9_io_out ? io_r_146_b : _GEN_2245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2247 = 8'h93 == r_count_9_io_out ? io_r_147_b : _GEN_2246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2248 = 8'h94 == r_count_9_io_out ? io_r_148_b : _GEN_2247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2249 = 8'h95 == r_count_9_io_out ? io_r_149_b : _GEN_2248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2250 = 8'h96 == r_count_9_io_out ? io_r_150_b : _GEN_2249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2251 = 8'h97 == r_count_9_io_out ? io_r_151_b : _GEN_2250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2252 = 8'h98 == r_count_9_io_out ? io_r_152_b : _GEN_2251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2253 = 8'h99 == r_count_9_io_out ? io_r_153_b : _GEN_2252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2254 = 8'h9a == r_count_9_io_out ? io_r_154_b : _GEN_2253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2255 = 8'h9b == r_count_9_io_out ? io_r_155_b : _GEN_2254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2256 = 8'h9c == r_count_9_io_out ? io_r_156_b : _GEN_2255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2257 = 8'h9d == r_count_9_io_out ? io_r_157_b : _GEN_2256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2258 = 8'h9e == r_count_9_io_out ? io_r_158_b : _GEN_2257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2259 = 8'h9f == r_count_9_io_out ? io_r_159_b : _GEN_2258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2260 = 8'ha0 == r_count_9_io_out ? io_r_160_b : _GEN_2259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2261 = 8'ha1 == r_count_9_io_out ? io_r_161_b : _GEN_2260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2262 = 8'ha2 == r_count_9_io_out ? io_r_162_b : _GEN_2261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2263 = 8'ha3 == r_count_9_io_out ? io_r_163_b : _GEN_2262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2264 = 8'ha4 == r_count_9_io_out ? io_r_164_b : _GEN_2263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2265 = 8'ha5 == r_count_9_io_out ? io_r_165_b : _GEN_2264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2266 = 8'ha6 == r_count_9_io_out ? io_r_166_b : _GEN_2265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2267 = 8'ha7 == r_count_9_io_out ? io_r_167_b : _GEN_2266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2268 = 8'ha8 == r_count_9_io_out ? io_r_168_b : _GEN_2267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2269 = 8'ha9 == r_count_9_io_out ? io_r_169_b : _GEN_2268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2270 = 8'haa == r_count_9_io_out ? io_r_170_b : _GEN_2269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2271 = 8'hab == r_count_9_io_out ? io_r_171_b : _GEN_2270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2272 = 8'hac == r_count_9_io_out ? io_r_172_b : _GEN_2271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2273 = 8'had == r_count_9_io_out ? io_r_173_b : _GEN_2272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2274 = 8'hae == r_count_9_io_out ? io_r_174_b : _GEN_2273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2275 = 8'haf == r_count_9_io_out ? io_r_175_b : _GEN_2274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2276 = 8'hb0 == r_count_9_io_out ? io_r_176_b : _GEN_2275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2277 = 8'hb1 == r_count_9_io_out ? io_r_177_b : _GEN_2276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2278 = 8'hb2 == r_count_9_io_out ? io_r_178_b : _GEN_2277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2279 = 8'hb3 == r_count_9_io_out ? io_r_179_b : _GEN_2278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2280 = 8'hb4 == r_count_9_io_out ? io_r_180_b : _GEN_2279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2281 = 8'hb5 == r_count_9_io_out ? io_r_181_b : _GEN_2280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2282 = 8'hb6 == r_count_9_io_out ? io_r_182_b : _GEN_2281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2283 = 8'hb7 == r_count_9_io_out ? io_r_183_b : _GEN_2282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2284 = 8'hb8 == r_count_9_io_out ? io_r_184_b : _GEN_2283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2285 = 8'hb9 == r_count_9_io_out ? io_r_185_b : _GEN_2284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2286 = 8'hba == r_count_9_io_out ? io_r_186_b : _GEN_2285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2287 = 8'hbb == r_count_9_io_out ? io_r_187_b : _GEN_2286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2288 = 8'hbc == r_count_9_io_out ? io_r_188_b : _GEN_2287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2289 = 8'hbd == r_count_9_io_out ? io_r_189_b : _GEN_2288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2290 = 8'hbe == r_count_9_io_out ? io_r_190_b : _GEN_2289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2291 = 8'hbf == r_count_9_io_out ? io_r_191_b : _GEN_2290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2292 = 8'hc0 == r_count_9_io_out ? io_r_192_b : _GEN_2291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2293 = 8'hc1 == r_count_9_io_out ? io_r_193_b : _GEN_2292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2294 = 8'hc2 == r_count_9_io_out ? io_r_194_b : _GEN_2293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2295 = 8'hc3 == r_count_9_io_out ? io_r_195_b : _GEN_2294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2296 = 8'hc4 == r_count_9_io_out ? io_r_196_b : _GEN_2295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2297 = 8'hc5 == r_count_9_io_out ? io_r_197_b : _GEN_2296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2298 = 8'hc6 == r_count_9_io_out ? io_r_198_b : _GEN_2297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2301 = 8'h1 == r_count_10_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2302 = 8'h2 == r_count_10_io_out ? io_r_2_b : _GEN_2301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2303 = 8'h3 == r_count_10_io_out ? io_r_3_b : _GEN_2302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2304 = 8'h4 == r_count_10_io_out ? io_r_4_b : _GEN_2303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2305 = 8'h5 == r_count_10_io_out ? io_r_5_b : _GEN_2304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2306 = 8'h6 == r_count_10_io_out ? io_r_6_b : _GEN_2305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2307 = 8'h7 == r_count_10_io_out ? io_r_7_b : _GEN_2306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2308 = 8'h8 == r_count_10_io_out ? io_r_8_b : _GEN_2307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2309 = 8'h9 == r_count_10_io_out ? io_r_9_b : _GEN_2308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2310 = 8'ha == r_count_10_io_out ? io_r_10_b : _GEN_2309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2311 = 8'hb == r_count_10_io_out ? io_r_11_b : _GEN_2310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2312 = 8'hc == r_count_10_io_out ? io_r_12_b : _GEN_2311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2313 = 8'hd == r_count_10_io_out ? io_r_13_b : _GEN_2312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2314 = 8'he == r_count_10_io_out ? io_r_14_b : _GEN_2313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2315 = 8'hf == r_count_10_io_out ? io_r_15_b : _GEN_2314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2316 = 8'h10 == r_count_10_io_out ? io_r_16_b : _GEN_2315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2317 = 8'h11 == r_count_10_io_out ? io_r_17_b : _GEN_2316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2318 = 8'h12 == r_count_10_io_out ? io_r_18_b : _GEN_2317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2319 = 8'h13 == r_count_10_io_out ? io_r_19_b : _GEN_2318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2320 = 8'h14 == r_count_10_io_out ? io_r_20_b : _GEN_2319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2321 = 8'h15 == r_count_10_io_out ? io_r_21_b : _GEN_2320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2322 = 8'h16 == r_count_10_io_out ? io_r_22_b : _GEN_2321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2323 = 8'h17 == r_count_10_io_out ? io_r_23_b : _GEN_2322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2324 = 8'h18 == r_count_10_io_out ? io_r_24_b : _GEN_2323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2325 = 8'h19 == r_count_10_io_out ? io_r_25_b : _GEN_2324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2326 = 8'h1a == r_count_10_io_out ? io_r_26_b : _GEN_2325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2327 = 8'h1b == r_count_10_io_out ? io_r_27_b : _GEN_2326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2328 = 8'h1c == r_count_10_io_out ? io_r_28_b : _GEN_2327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2329 = 8'h1d == r_count_10_io_out ? io_r_29_b : _GEN_2328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2330 = 8'h1e == r_count_10_io_out ? io_r_30_b : _GEN_2329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2331 = 8'h1f == r_count_10_io_out ? io_r_31_b : _GEN_2330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2332 = 8'h20 == r_count_10_io_out ? io_r_32_b : _GEN_2331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2333 = 8'h21 == r_count_10_io_out ? io_r_33_b : _GEN_2332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2334 = 8'h22 == r_count_10_io_out ? io_r_34_b : _GEN_2333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2335 = 8'h23 == r_count_10_io_out ? io_r_35_b : _GEN_2334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2336 = 8'h24 == r_count_10_io_out ? io_r_36_b : _GEN_2335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2337 = 8'h25 == r_count_10_io_out ? io_r_37_b : _GEN_2336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2338 = 8'h26 == r_count_10_io_out ? io_r_38_b : _GEN_2337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2339 = 8'h27 == r_count_10_io_out ? io_r_39_b : _GEN_2338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2340 = 8'h28 == r_count_10_io_out ? io_r_40_b : _GEN_2339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2341 = 8'h29 == r_count_10_io_out ? io_r_41_b : _GEN_2340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2342 = 8'h2a == r_count_10_io_out ? io_r_42_b : _GEN_2341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2343 = 8'h2b == r_count_10_io_out ? io_r_43_b : _GEN_2342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2344 = 8'h2c == r_count_10_io_out ? io_r_44_b : _GEN_2343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2345 = 8'h2d == r_count_10_io_out ? io_r_45_b : _GEN_2344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2346 = 8'h2e == r_count_10_io_out ? io_r_46_b : _GEN_2345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2347 = 8'h2f == r_count_10_io_out ? io_r_47_b : _GEN_2346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2348 = 8'h30 == r_count_10_io_out ? io_r_48_b : _GEN_2347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2349 = 8'h31 == r_count_10_io_out ? io_r_49_b : _GEN_2348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2350 = 8'h32 == r_count_10_io_out ? io_r_50_b : _GEN_2349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2351 = 8'h33 == r_count_10_io_out ? io_r_51_b : _GEN_2350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2352 = 8'h34 == r_count_10_io_out ? io_r_52_b : _GEN_2351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2353 = 8'h35 == r_count_10_io_out ? io_r_53_b : _GEN_2352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2354 = 8'h36 == r_count_10_io_out ? io_r_54_b : _GEN_2353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2355 = 8'h37 == r_count_10_io_out ? io_r_55_b : _GEN_2354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2356 = 8'h38 == r_count_10_io_out ? io_r_56_b : _GEN_2355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2357 = 8'h39 == r_count_10_io_out ? io_r_57_b : _GEN_2356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2358 = 8'h3a == r_count_10_io_out ? io_r_58_b : _GEN_2357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2359 = 8'h3b == r_count_10_io_out ? io_r_59_b : _GEN_2358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2360 = 8'h3c == r_count_10_io_out ? io_r_60_b : _GEN_2359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2361 = 8'h3d == r_count_10_io_out ? io_r_61_b : _GEN_2360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2362 = 8'h3e == r_count_10_io_out ? io_r_62_b : _GEN_2361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2363 = 8'h3f == r_count_10_io_out ? io_r_63_b : _GEN_2362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2364 = 8'h40 == r_count_10_io_out ? io_r_64_b : _GEN_2363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2365 = 8'h41 == r_count_10_io_out ? io_r_65_b : _GEN_2364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2366 = 8'h42 == r_count_10_io_out ? io_r_66_b : _GEN_2365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2367 = 8'h43 == r_count_10_io_out ? io_r_67_b : _GEN_2366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2368 = 8'h44 == r_count_10_io_out ? io_r_68_b : _GEN_2367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2369 = 8'h45 == r_count_10_io_out ? io_r_69_b : _GEN_2368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2370 = 8'h46 == r_count_10_io_out ? io_r_70_b : _GEN_2369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2371 = 8'h47 == r_count_10_io_out ? io_r_71_b : _GEN_2370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2372 = 8'h48 == r_count_10_io_out ? io_r_72_b : _GEN_2371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2373 = 8'h49 == r_count_10_io_out ? io_r_73_b : _GEN_2372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2374 = 8'h4a == r_count_10_io_out ? io_r_74_b : _GEN_2373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2375 = 8'h4b == r_count_10_io_out ? io_r_75_b : _GEN_2374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2376 = 8'h4c == r_count_10_io_out ? io_r_76_b : _GEN_2375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2377 = 8'h4d == r_count_10_io_out ? io_r_77_b : _GEN_2376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2378 = 8'h4e == r_count_10_io_out ? io_r_78_b : _GEN_2377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2379 = 8'h4f == r_count_10_io_out ? io_r_79_b : _GEN_2378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2380 = 8'h50 == r_count_10_io_out ? io_r_80_b : _GEN_2379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2381 = 8'h51 == r_count_10_io_out ? io_r_81_b : _GEN_2380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2382 = 8'h52 == r_count_10_io_out ? io_r_82_b : _GEN_2381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2383 = 8'h53 == r_count_10_io_out ? io_r_83_b : _GEN_2382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2384 = 8'h54 == r_count_10_io_out ? io_r_84_b : _GEN_2383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2385 = 8'h55 == r_count_10_io_out ? io_r_85_b : _GEN_2384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2386 = 8'h56 == r_count_10_io_out ? io_r_86_b : _GEN_2385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2387 = 8'h57 == r_count_10_io_out ? io_r_87_b : _GEN_2386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2388 = 8'h58 == r_count_10_io_out ? io_r_88_b : _GEN_2387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2389 = 8'h59 == r_count_10_io_out ? io_r_89_b : _GEN_2388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2390 = 8'h5a == r_count_10_io_out ? io_r_90_b : _GEN_2389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2391 = 8'h5b == r_count_10_io_out ? io_r_91_b : _GEN_2390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2392 = 8'h5c == r_count_10_io_out ? io_r_92_b : _GEN_2391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2393 = 8'h5d == r_count_10_io_out ? io_r_93_b : _GEN_2392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2394 = 8'h5e == r_count_10_io_out ? io_r_94_b : _GEN_2393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2395 = 8'h5f == r_count_10_io_out ? io_r_95_b : _GEN_2394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2396 = 8'h60 == r_count_10_io_out ? io_r_96_b : _GEN_2395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2397 = 8'h61 == r_count_10_io_out ? io_r_97_b : _GEN_2396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2398 = 8'h62 == r_count_10_io_out ? io_r_98_b : _GEN_2397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2399 = 8'h63 == r_count_10_io_out ? io_r_99_b : _GEN_2398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2400 = 8'h64 == r_count_10_io_out ? io_r_100_b : _GEN_2399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2401 = 8'h65 == r_count_10_io_out ? io_r_101_b : _GEN_2400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2402 = 8'h66 == r_count_10_io_out ? io_r_102_b : _GEN_2401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2403 = 8'h67 == r_count_10_io_out ? io_r_103_b : _GEN_2402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2404 = 8'h68 == r_count_10_io_out ? io_r_104_b : _GEN_2403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2405 = 8'h69 == r_count_10_io_out ? io_r_105_b : _GEN_2404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2406 = 8'h6a == r_count_10_io_out ? io_r_106_b : _GEN_2405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2407 = 8'h6b == r_count_10_io_out ? io_r_107_b : _GEN_2406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2408 = 8'h6c == r_count_10_io_out ? io_r_108_b : _GEN_2407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2409 = 8'h6d == r_count_10_io_out ? io_r_109_b : _GEN_2408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2410 = 8'h6e == r_count_10_io_out ? io_r_110_b : _GEN_2409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2411 = 8'h6f == r_count_10_io_out ? io_r_111_b : _GEN_2410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2412 = 8'h70 == r_count_10_io_out ? io_r_112_b : _GEN_2411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2413 = 8'h71 == r_count_10_io_out ? io_r_113_b : _GEN_2412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2414 = 8'h72 == r_count_10_io_out ? io_r_114_b : _GEN_2413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2415 = 8'h73 == r_count_10_io_out ? io_r_115_b : _GEN_2414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2416 = 8'h74 == r_count_10_io_out ? io_r_116_b : _GEN_2415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2417 = 8'h75 == r_count_10_io_out ? io_r_117_b : _GEN_2416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2418 = 8'h76 == r_count_10_io_out ? io_r_118_b : _GEN_2417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2419 = 8'h77 == r_count_10_io_out ? io_r_119_b : _GEN_2418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2420 = 8'h78 == r_count_10_io_out ? io_r_120_b : _GEN_2419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2421 = 8'h79 == r_count_10_io_out ? io_r_121_b : _GEN_2420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2422 = 8'h7a == r_count_10_io_out ? io_r_122_b : _GEN_2421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2423 = 8'h7b == r_count_10_io_out ? io_r_123_b : _GEN_2422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2424 = 8'h7c == r_count_10_io_out ? io_r_124_b : _GEN_2423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2425 = 8'h7d == r_count_10_io_out ? io_r_125_b : _GEN_2424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2426 = 8'h7e == r_count_10_io_out ? io_r_126_b : _GEN_2425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2427 = 8'h7f == r_count_10_io_out ? io_r_127_b : _GEN_2426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2428 = 8'h80 == r_count_10_io_out ? io_r_128_b : _GEN_2427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2429 = 8'h81 == r_count_10_io_out ? io_r_129_b : _GEN_2428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2430 = 8'h82 == r_count_10_io_out ? io_r_130_b : _GEN_2429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2431 = 8'h83 == r_count_10_io_out ? io_r_131_b : _GEN_2430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2432 = 8'h84 == r_count_10_io_out ? io_r_132_b : _GEN_2431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2433 = 8'h85 == r_count_10_io_out ? io_r_133_b : _GEN_2432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2434 = 8'h86 == r_count_10_io_out ? io_r_134_b : _GEN_2433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2435 = 8'h87 == r_count_10_io_out ? io_r_135_b : _GEN_2434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2436 = 8'h88 == r_count_10_io_out ? io_r_136_b : _GEN_2435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2437 = 8'h89 == r_count_10_io_out ? io_r_137_b : _GEN_2436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2438 = 8'h8a == r_count_10_io_out ? io_r_138_b : _GEN_2437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2439 = 8'h8b == r_count_10_io_out ? io_r_139_b : _GEN_2438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2440 = 8'h8c == r_count_10_io_out ? io_r_140_b : _GEN_2439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2441 = 8'h8d == r_count_10_io_out ? io_r_141_b : _GEN_2440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2442 = 8'h8e == r_count_10_io_out ? io_r_142_b : _GEN_2441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2443 = 8'h8f == r_count_10_io_out ? io_r_143_b : _GEN_2442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2444 = 8'h90 == r_count_10_io_out ? io_r_144_b : _GEN_2443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2445 = 8'h91 == r_count_10_io_out ? io_r_145_b : _GEN_2444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2446 = 8'h92 == r_count_10_io_out ? io_r_146_b : _GEN_2445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2447 = 8'h93 == r_count_10_io_out ? io_r_147_b : _GEN_2446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2448 = 8'h94 == r_count_10_io_out ? io_r_148_b : _GEN_2447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2449 = 8'h95 == r_count_10_io_out ? io_r_149_b : _GEN_2448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2450 = 8'h96 == r_count_10_io_out ? io_r_150_b : _GEN_2449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2451 = 8'h97 == r_count_10_io_out ? io_r_151_b : _GEN_2450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2452 = 8'h98 == r_count_10_io_out ? io_r_152_b : _GEN_2451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2453 = 8'h99 == r_count_10_io_out ? io_r_153_b : _GEN_2452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2454 = 8'h9a == r_count_10_io_out ? io_r_154_b : _GEN_2453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2455 = 8'h9b == r_count_10_io_out ? io_r_155_b : _GEN_2454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2456 = 8'h9c == r_count_10_io_out ? io_r_156_b : _GEN_2455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2457 = 8'h9d == r_count_10_io_out ? io_r_157_b : _GEN_2456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2458 = 8'h9e == r_count_10_io_out ? io_r_158_b : _GEN_2457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2459 = 8'h9f == r_count_10_io_out ? io_r_159_b : _GEN_2458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2460 = 8'ha0 == r_count_10_io_out ? io_r_160_b : _GEN_2459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2461 = 8'ha1 == r_count_10_io_out ? io_r_161_b : _GEN_2460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2462 = 8'ha2 == r_count_10_io_out ? io_r_162_b : _GEN_2461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2463 = 8'ha3 == r_count_10_io_out ? io_r_163_b : _GEN_2462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2464 = 8'ha4 == r_count_10_io_out ? io_r_164_b : _GEN_2463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2465 = 8'ha5 == r_count_10_io_out ? io_r_165_b : _GEN_2464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2466 = 8'ha6 == r_count_10_io_out ? io_r_166_b : _GEN_2465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2467 = 8'ha7 == r_count_10_io_out ? io_r_167_b : _GEN_2466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2468 = 8'ha8 == r_count_10_io_out ? io_r_168_b : _GEN_2467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2469 = 8'ha9 == r_count_10_io_out ? io_r_169_b : _GEN_2468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2470 = 8'haa == r_count_10_io_out ? io_r_170_b : _GEN_2469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2471 = 8'hab == r_count_10_io_out ? io_r_171_b : _GEN_2470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2472 = 8'hac == r_count_10_io_out ? io_r_172_b : _GEN_2471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2473 = 8'had == r_count_10_io_out ? io_r_173_b : _GEN_2472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2474 = 8'hae == r_count_10_io_out ? io_r_174_b : _GEN_2473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2475 = 8'haf == r_count_10_io_out ? io_r_175_b : _GEN_2474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2476 = 8'hb0 == r_count_10_io_out ? io_r_176_b : _GEN_2475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2477 = 8'hb1 == r_count_10_io_out ? io_r_177_b : _GEN_2476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2478 = 8'hb2 == r_count_10_io_out ? io_r_178_b : _GEN_2477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2479 = 8'hb3 == r_count_10_io_out ? io_r_179_b : _GEN_2478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2480 = 8'hb4 == r_count_10_io_out ? io_r_180_b : _GEN_2479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2481 = 8'hb5 == r_count_10_io_out ? io_r_181_b : _GEN_2480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2482 = 8'hb6 == r_count_10_io_out ? io_r_182_b : _GEN_2481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2483 = 8'hb7 == r_count_10_io_out ? io_r_183_b : _GEN_2482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2484 = 8'hb8 == r_count_10_io_out ? io_r_184_b : _GEN_2483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2485 = 8'hb9 == r_count_10_io_out ? io_r_185_b : _GEN_2484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2486 = 8'hba == r_count_10_io_out ? io_r_186_b : _GEN_2485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2487 = 8'hbb == r_count_10_io_out ? io_r_187_b : _GEN_2486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2488 = 8'hbc == r_count_10_io_out ? io_r_188_b : _GEN_2487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2489 = 8'hbd == r_count_10_io_out ? io_r_189_b : _GEN_2488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2490 = 8'hbe == r_count_10_io_out ? io_r_190_b : _GEN_2489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2491 = 8'hbf == r_count_10_io_out ? io_r_191_b : _GEN_2490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2492 = 8'hc0 == r_count_10_io_out ? io_r_192_b : _GEN_2491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2493 = 8'hc1 == r_count_10_io_out ? io_r_193_b : _GEN_2492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2494 = 8'hc2 == r_count_10_io_out ? io_r_194_b : _GEN_2493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2495 = 8'hc3 == r_count_10_io_out ? io_r_195_b : _GEN_2494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2496 = 8'hc4 == r_count_10_io_out ? io_r_196_b : _GEN_2495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2497 = 8'hc5 == r_count_10_io_out ? io_r_197_b : _GEN_2496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2498 = 8'hc6 == r_count_10_io_out ? io_r_198_b : _GEN_2497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2501 = 8'h1 == r_count_11_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2502 = 8'h2 == r_count_11_io_out ? io_r_2_b : _GEN_2501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2503 = 8'h3 == r_count_11_io_out ? io_r_3_b : _GEN_2502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2504 = 8'h4 == r_count_11_io_out ? io_r_4_b : _GEN_2503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2505 = 8'h5 == r_count_11_io_out ? io_r_5_b : _GEN_2504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2506 = 8'h6 == r_count_11_io_out ? io_r_6_b : _GEN_2505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2507 = 8'h7 == r_count_11_io_out ? io_r_7_b : _GEN_2506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2508 = 8'h8 == r_count_11_io_out ? io_r_8_b : _GEN_2507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2509 = 8'h9 == r_count_11_io_out ? io_r_9_b : _GEN_2508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2510 = 8'ha == r_count_11_io_out ? io_r_10_b : _GEN_2509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2511 = 8'hb == r_count_11_io_out ? io_r_11_b : _GEN_2510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2512 = 8'hc == r_count_11_io_out ? io_r_12_b : _GEN_2511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2513 = 8'hd == r_count_11_io_out ? io_r_13_b : _GEN_2512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2514 = 8'he == r_count_11_io_out ? io_r_14_b : _GEN_2513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2515 = 8'hf == r_count_11_io_out ? io_r_15_b : _GEN_2514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2516 = 8'h10 == r_count_11_io_out ? io_r_16_b : _GEN_2515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2517 = 8'h11 == r_count_11_io_out ? io_r_17_b : _GEN_2516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2518 = 8'h12 == r_count_11_io_out ? io_r_18_b : _GEN_2517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2519 = 8'h13 == r_count_11_io_out ? io_r_19_b : _GEN_2518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2520 = 8'h14 == r_count_11_io_out ? io_r_20_b : _GEN_2519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2521 = 8'h15 == r_count_11_io_out ? io_r_21_b : _GEN_2520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2522 = 8'h16 == r_count_11_io_out ? io_r_22_b : _GEN_2521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2523 = 8'h17 == r_count_11_io_out ? io_r_23_b : _GEN_2522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2524 = 8'h18 == r_count_11_io_out ? io_r_24_b : _GEN_2523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2525 = 8'h19 == r_count_11_io_out ? io_r_25_b : _GEN_2524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2526 = 8'h1a == r_count_11_io_out ? io_r_26_b : _GEN_2525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2527 = 8'h1b == r_count_11_io_out ? io_r_27_b : _GEN_2526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2528 = 8'h1c == r_count_11_io_out ? io_r_28_b : _GEN_2527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2529 = 8'h1d == r_count_11_io_out ? io_r_29_b : _GEN_2528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2530 = 8'h1e == r_count_11_io_out ? io_r_30_b : _GEN_2529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2531 = 8'h1f == r_count_11_io_out ? io_r_31_b : _GEN_2530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2532 = 8'h20 == r_count_11_io_out ? io_r_32_b : _GEN_2531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2533 = 8'h21 == r_count_11_io_out ? io_r_33_b : _GEN_2532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2534 = 8'h22 == r_count_11_io_out ? io_r_34_b : _GEN_2533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2535 = 8'h23 == r_count_11_io_out ? io_r_35_b : _GEN_2534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2536 = 8'h24 == r_count_11_io_out ? io_r_36_b : _GEN_2535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2537 = 8'h25 == r_count_11_io_out ? io_r_37_b : _GEN_2536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2538 = 8'h26 == r_count_11_io_out ? io_r_38_b : _GEN_2537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2539 = 8'h27 == r_count_11_io_out ? io_r_39_b : _GEN_2538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2540 = 8'h28 == r_count_11_io_out ? io_r_40_b : _GEN_2539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2541 = 8'h29 == r_count_11_io_out ? io_r_41_b : _GEN_2540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2542 = 8'h2a == r_count_11_io_out ? io_r_42_b : _GEN_2541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2543 = 8'h2b == r_count_11_io_out ? io_r_43_b : _GEN_2542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2544 = 8'h2c == r_count_11_io_out ? io_r_44_b : _GEN_2543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2545 = 8'h2d == r_count_11_io_out ? io_r_45_b : _GEN_2544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2546 = 8'h2e == r_count_11_io_out ? io_r_46_b : _GEN_2545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2547 = 8'h2f == r_count_11_io_out ? io_r_47_b : _GEN_2546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2548 = 8'h30 == r_count_11_io_out ? io_r_48_b : _GEN_2547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2549 = 8'h31 == r_count_11_io_out ? io_r_49_b : _GEN_2548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2550 = 8'h32 == r_count_11_io_out ? io_r_50_b : _GEN_2549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2551 = 8'h33 == r_count_11_io_out ? io_r_51_b : _GEN_2550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2552 = 8'h34 == r_count_11_io_out ? io_r_52_b : _GEN_2551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2553 = 8'h35 == r_count_11_io_out ? io_r_53_b : _GEN_2552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2554 = 8'h36 == r_count_11_io_out ? io_r_54_b : _GEN_2553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2555 = 8'h37 == r_count_11_io_out ? io_r_55_b : _GEN_2554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2556 = 8'h38 == r_count_11_io_out ? io_r_56_b : _GEN_2555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2557 = 8'h39 == r_count_11_io_out ? io_r_57_b : _GEN_2556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2558 = 8'h3a == r_count_11_io_out ? io_r_58_b : _GEN_2557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2559 = 8'h3b == r_count_11_io_out ? io_r_59_b : _GEN_2558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2560 = 8'h3c == r_count_11_io_out ? io_r_60_b : _GEN_2559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2561 = 8'h3d == r_count_11_io_out ? io_r_61_b : _GEN_2560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2562 = 8'h3e == r_count_11_io_out ? io_r_62_b : _GEN_2561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2563 = 8'h3f == r_count_11_io_out ? io_r_63_b : _GEN_2562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2564 = 8'h40 == r_count_11_io_out ? io_r_64_b : _GEN_2563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2565 = 8'h41 == r_count_11_io_out ? io_r_65_b : _GEN_2564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2566 = 8'h42 == r_count_11_io_out ? io_r_66_b : _GEN_2565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2567 = 8'h43 == r_count_11_io_out ? io_r_67_b : _GEN_2566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2568 = 8'h44 == r_count_11_io_out ? io_r_68_b : _GEN_2567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2569 = 8'h45 == r_count_11_io_out ? io_r_69_b : _GEN_2568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2570 = 8'h46 == r_count_11_io_out ? io_r_70_b : _GEN_2569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2571 = 8'h47 == r_count_11_io_out ? io_r_71_b : _GEN_2570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2572 = 8'h48 == r_count_11_io_out ? io_r_72_b : _GEN_2571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2573 = 8'h49 == r_count_11_io_out ? io_r_73_b : _GEN_2572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2574 = 8'h4a == r_count_11_io_out ? io_r_74_b : _GEN_2573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2575 = 8'h4b == r_count_11_io_out ? io_r_75_b : _GEN_2574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2576 = 8'h4c == r_count_11_io_out ? io_r_76_b : _GEN_2575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2577 = 8'h4d == r_count_11_io_out ? io_r_77_b : _GEN_2576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2578 = 8'h4e == r_count_11_io_out ? io_r_78_b : _GEN_2577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2579 = 8'h4f == r_count_11_io_out ? io_r_79_b : _GEN_2578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2580 = 8'h50 == r_count_11_io_out ? io_r_80_b : _GEN_2579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2581 = 8'h51 == r_count_11_io_out ? io_r_81_b : _GEN_2580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2582 = 8'h52 == r_count_11_io_out ? io_r_82_b : _GEN_2581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2583 = 8'h53 == r_count_11_io_out ? io_r_83_b : _GEN_2582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2584 = 8'h54 == r_count_11_io_out ? io_r_84_b : _GEN_2583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2585 = 8'h55 == r_count_11_io_out ? io_r_85_b : _GEN_2584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2586 = 8'h56 == r_count_11_io_out ? io_r_86_b : _GEN_2585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2587 = 8'h57 == r_count_11_io_out ? io_r_87_b : _GEN_2586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2588 = 8'h58 == r_count_11_io_out ? io_r_88_b : _GEN_2587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2589 = 8'h59 == r_count_11_io_out ? io_r_89_b : _GEN_2588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2590 = 8'h5a == r_count_11_io_out ? io_r_90_b : _GEN_2589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2591 = 8'h5b == r_count_11_io_out ? io_r_91_b : _GEN_2590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2592 = 8'h5c == r_count_11_io_out ? io_r_92_b : _GEN_2591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2593 = 8'h5d == r_count_11_io_out ? io_r_93_b : _GEN_2592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2594 = 8'h5e == r_count_11_io_out ? io_r_94_b : _GEN_2593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2595 = 8'h5f == r_count_11_io_out ? io_r_95_b : _GEN_2594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2596 = 8'h60 == r_count_11_io_out ? io_r_96_b : _GEN_2595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2597 = 8'h61 == r_count_11_io_out ? io_r_97_b : _GEN_2596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2598 = 8'h62 == r_count_11_io_out ? io_r_98_b : _GEN_2597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2599 = 8'h63 == r_count_11_io_out ? io_r_99_b : _GEN_2598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2600 = 8'h64 == r_count_11_io_out ? io_r_100_b : _GEN_2599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2601 = 8'h65 == r_count_11_io_out ? io_r_101_b : _GEN_2600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2602 = 8'h66 == r_count_11_io_out ? io_r_102_b : _GEN_2601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2603 = 8'h67 == r_count_11_io_out ? io_r_103_b : _GEN_2602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2604 = 8'h68 == r_count_11_io_out ? io_r_104_b : _GEN_2603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2605 = 8'h69 == r_count_11_io_out ? io_r_105_b : _GEN_2604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2606 = 8'h6a == r_count_11_io_out ? io_r_106_b : _GEN_2605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2607 = 8'h6b == r_count_11_io_out ? io_r_107_b : _GEN_2606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2608 = 8'h6c == r_count_11_io_out ? io_r_108_b : _GEN_2607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2609 = 8'h6d == r_count_11_io_out ? io_r_109_b : _GEN_2608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2610 = 8'h6e == r_count_11_io_out ? io_r_110_b : _GEN_2609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2611 = 8'h6f == r_count_11_io_out ? io_r_111_b : _GEN_2610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2612 = 8'h70 == r_count_11_io_out ? io_r_112_b : _GEN_2611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2613 = 8'h71 == r_count_11_io_out ? io_r_113_b : _GEN_2612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2614 = 8'h72 == r_count_11_io_out ? io_r_114_b : _GEN_2613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2615 = 8'h73 == r_count_11_io_out ? io_r_115_b : _GEN_2614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2616 = 8'h74 == r_count_11_io_out ? io_r_116_b : _GEN_2615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2617 = 8'h75 == r_count_11_io_out ? io_r_117_b : _GEN_2616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2618 = 8'h76 == r_count_11_io_out ? io_r_118_b : _GEN_2617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2619 = 8'h77 == r_count_11_io_out ? io_r_119_b : _GEN_2618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2620 = 8'h78 == r_count_11_io_out ? io_r_120_b : _GEN_2619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2621 = 8'h79 == r_count_11_io_out ? io_r_121_b : _GEN_2620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2622 = 8'h7a == r_count_11_io_out ? io_r_122_b : _GEN_2621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2623 = 8'h7b == r_count_11_io_out ? io_r_123_b : _GEN_2622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2624 = 8'h7c == r_count_11_io_out ? io_r_124_b : _GEN_2623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2625 = 8'h7d == r_count_11_io_out ? io_r_125_b : _GEN_2624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2626 = 8'h7e == r_count_11_io_out ? io_r_126_b : _GEN_2625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2627 = 8'h7f == r_count_11_io_out ? io_r_127_b : _GEN_2626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2628 = 8'h80 == r_count_11_io_out ? io_r_128_b : _GEN_2627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2629 = 8'h81 == r_count_11_io_out ? io_r_129_b : _GEN_2628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2630 = 8'h82 == r_count_11_io_out ? io_r_130_b : _GEN_2629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2631 = 8'h83 == r_count_11_io_out ? io_r_131_b : _GEN_2630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2632 = 8'h84 == r_count_11_io_out ? io_r_132_b : _GEN_2631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2633 = 8'h85 == r_count_11_io_out ? io_r_133_b : _GEN_2632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2634 = 8'h86 == r_count_11_io_out ? io_r_134_b : _GEN_2633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2635 = 8'h87 == r_count_11_io_out ? io_r_135_b : _GEN_2634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2636 = 8'h88 == r_count_11_io_out ? io_r_136_b : _GEN_2635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2637 = 8'h89 == r_count_11_io_out ? io_r_137_b : _GEN_2636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2638 = 8'h8a == r_count_11_io_out ? io_r_138_b : _GEN_2637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2639 = 8'h8b == r_count_11_io_out ? io_r_139_b : _GEN_2638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2640 = 8'h8c == r_count_11_io_out ? io_r_140_b : _GEN_2639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2641 = 8'h8d == r_count_11_io_out ? io_r_141_b : _GEN_2640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2642 = 8'h8e == r_count_11_io_out ? io_r_142_b : _GEN_2641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2643 = 8'h8f == r_count_11_io_out ? io_r_143_b : _GEN_2642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2644 = 8'h90 == r_count_11_io_out ? io_r_144_b : _GEN_2643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2645 = 8'h91 == r_count_11_io_out ? io_r_145_b : _GEN_2644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2646 = 8'h92 == r_count_11_io_out ? io_r_146_b : _GEN_2645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2647 = 8'h93 == r_count_11_io_out ? io_r_147_b : _GEN_2646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2648 = 8'h94 == r_count_11_io_out ? io_r_148_b : _GEN_2647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2649 = 8'h95 == r_count_11_io_out ? io_r_149_b : _GEN_2648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2650 = 8'h96 == r_count_11_io_out ? io_r_150_b : _GEN_2649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2651 = 8'h97 == r_count_11_io_out ? io_r_151_b : _GEN_2650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2652 = 8'h98 == r_count_11_io_out ? io_r_152_b : _GEN_2651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2653 = 8'h99 == r_count_11_io_out ? io_r_153_b : _GEN_2652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2654 = 8'h9a == r_count_11_io_out ? io_r_154_b : _GEN_2653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2655 = 8'h9b == r_count_11_io_out ? io_r_155_b : _GEN_2654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2656 = 8'h9c == r_count_11_io_out ? io_r_156_b : _GEN_2655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2657 = 8'h9d == r_count_11_io_out ? io_r_157_b : _GEN_2656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2658 = 8'h9e == r_count_11_io_out ? io_r_158_b : _GEN_2657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2659 = 8'h9f == r_count_11_io_out ? io_r_159_b : _GEN_2658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2660 = 8'ha0 == r_count_11_io_out ? io_r_160_b : _GEN_2659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2661 = 8'ha1 == r_count_11_io_out ? io_r_161_b : _GEN_2660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2662 = 8'ha2 == r_count_11_io_out ? io_r_162_b : _GEN_2661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2663 = 8'ha3 == r_count_11_io_out ? io_r_163_b : _GEN_2662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2664 = 8'ha4 == r_count_11_io_out ? io_r_164_b : _GEN_2663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2665 = 8'ha5 == r_count_11_io_out ? io_r_165_b : _GEN_2664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2666 = 8'ha6 == r_count_11_io_out ? io_r_166_b : _GEN_2665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2667 = 8'ha7 == r_count_11_io_out ? io_r_167_b : _GEN_2666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2668 = 8'ha8 == r_count_11_io_out ? io_r_168_b : _GEN_2667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2669 = 8'ha9 == r_count_11_io_out ? io_r_169_b : _GEN_2668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2670 = 8'haa == r_count_11_io_out ? io_r_170_b : _GEN_2669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2671 = 8'hab == r_count_11_io_out ? io_r_171_b : _GEN_2670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2672 = 8'hac == r_count_11_io_out ? io_r_172_b : _GEN_2671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2673 = 8'had == r_count_11_io_out ? io_r_173_b : _GEN_2672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2674 = 8'hae == r_count_11_io_out ? io_r_174_b : _GEN_2673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2675 = 8'haf == r_count_11_io_out ? io_r_175_b : _GEN_2674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2676 = 8'hb0 == r_count_11_io_out ? io_r_176_b : _GEN_2675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2677 = 8'hb1 == r_count_11_io_out ? io_r_177_b : _GEN_2676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2678 = 8'hb2 == r_count_11_io_out ? io_r_178_b : _GEN_2677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2679 = 8'hb3 == r_count_11_io_out ? io_r_179_b : _GEN_2678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2680 = 8'hb4 == r_count_11_io_out ? io_r_180_b : _GEN_2679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2681 = 8'hb5 == r_count_11_io_out ? io_r_181_b : _GEN_2680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2682 = 8'hb6 == r_count_11_io_out ? io_r_182_b : _GEN_2681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2683 = 8'hb7 == r_count_11_io_out ? io_r_183_b : _GEN_2682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2684 = 8'hb8 == r_count_11_io_out ? io_r_184_b : _GEN_2683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2685 = 8'hb9 == r_count_11_io_out ? io_r_185_b : _GEN_2684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2686 = 8'hba == r_count_11_io_out ? io_r_186_b : _GEN_2685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2687 = 8'hbb == r_count_11_io_out ? io_r_187_b : _GEN_2686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2688 = 8'hbc == r_count_11_io_out ? io_r_188_b : _GEN_2687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2689 = 8'hbd == r_count_11_io_out ? io_r_189_b : _GEN_2688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2690 = 8'hbe == r_count_11_io_out ? io_r_190_b : _GEN_2689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2691 = 8'hbf == r_count_11_io_out ? io_r_191_b : _GEN_2690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2692 = 8'hc0 == r_count_11_io_out ? io_r_192_b : _GEN_2691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2693 = 8'hc1 == r_count_11_io_out ? io_r_193_b : _GEN_2692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2694 = 8'hc2 == r_count_11_io_out ? io_r_194_b : _GEN_2693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2695 = 8'hc3 == r_count_11_io_out ? io_r_195_b : _GEN_2694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2696 = 8'hc4 == r_count_11_io_out ? io_r_196_b : _GEN_2695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2697 = 8'hc5 == r_count_11_io_out ? io_r_197_b : _GEN_2696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2698 = 8'hc6 == r_count_11_io_out ? io_r_198_b : _GEN_2697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2701 = 8'h1 == r_count_12_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2702 = 8'h2 == r_count_12_io_out ? io_r_2_b : _GEN_2701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2703 = 8'h3 == r_count_12_io_out ? io_r_3_b : _GEN_2702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2704 = 8'h4 == r_count_12_io_out ? io_r_4_b : _GEN_2703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2705 = 8'h5 == r_count_12_io_out ? io_r_5_b : _GEN_2704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2706 = 8'h6 == r_count_12_io_out ? io_r_6_b : _GEN_2705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2707 = 8'h7 == r_count_12_io_out ? io_r_7_b : _GEN_2706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2708 = 8'h8 == r_count_12_io_out ? io_r_8_b : _GEN_2707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2709 = 8'h9 == r_count_12_io_out ? io_r_9_b : _GEN_2708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2710 = 8'ha == r_count_12_io_out ? io_r_10_b : _GEN_2709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2711 = 8'hb == r_count_12_io_out ? io_r_11_b : _GEN_2710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2712 = 8'hc == r_count_12_io_out ? io_r_12_b : _GEN_2711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2713 = 8'hd == r_count_12_io_out ? io_r_13_b : _GEN_2712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2714 = 8'he == r_count_12_io_out ? io_r_14_b : _GEN_2713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2715 = 8'hf == r_count_12_io_out ? io_r_15_b : _GEN_2714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2716 = 8'h10 == r_count_12_io_out ? io_r_16_b : _GEN_2715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2717 = 8'h11 == r_count_12_io_out ? io_r_17_b : _GEN_2716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2718 = 8'h12 == r_count_12_io_out ? io_r_18_b : _GEN_2717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2719 = 8'h13 == r_count_12_io_out ? io_r_19_b : _GEN_2718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2720 = 8'h14 == r_count_12_io_out ? io_r_20_b : _GEN_2719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2721 = 8'h15 == r_count_12_io_out ? io_r_21_b : _GEN_2720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2722 = 8'h16 == r_count_12_io_out ? io_r_22_b : _GEN_2721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2723 = 8'h17 == r_count_12_io_out ? io_r_23_b : _GEN_2722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2724 = 8'h18 == r_count_12_io_out ? io_r_24_b : _GEN_2723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2725 = 8'h19 == r_count_12_io_out ? io_r_25_b : _GEN_2724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2726 = 8'h1a == r_count_12_io_out ? io_r_26_b : _GEN_2725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2727 = 8'h1b == r_count_12_io_out ? io_r_27_b : _GEN_2726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2728 = 8'h1c == r_count_12_io_out ? io_r_28_b : _GEN_2727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2729 = 8'h1d == r_count_12_io_out ? io_r_29_b : _GEN_2728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2730 = 8'h1e == r_count_12_io_out ? io_r_30_b : _GEN_2729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2731 = 8'h1f == r_count_12_io_out ? io_r_31_b : _GEN_2730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2732 = 8'h20 == r_count_12_io_out ? io_r_32_b : _GEN_2731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2733 = 8'h21 == r_count_12_io_out ? io_r_33_b : _GEN_2732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2734 = 8'h22 == r_count_12_io_out ? io_r_34_b : _GEN_2733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2735 = 8'h23 == r_count_12_io_out ? io_r_35_b : _GEN_2734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2736 = 8'h24 == r_count_12_io_out ? io_r_36_b : _GEN_2735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2737 = 8'h25 == r_count_12_io_out ? io_r_37_b : _GEN_2736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2738 = 8'h26 == r_count_12_io_out ? io_r_38_b : _GEN_2737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2739 = 8'h27 == r_count_12_io_out ? io_r_39_b : _GEN_2738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2740 = 8'h28 == r_count_12_io_out ? io_r_40_b : _GEN_2739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2741 = 8'h29 == r_count_12_io_out ? io_r_41_b : _GEN_2740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2742 = 8'h2a == r_count_12_io_out ? io_r_42_b : _GEN_2741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2743 = 8'h2b == r_count_12_io_out ? io_r_43_b : _GEN_2742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2744 = 8'h2c == r_count_12_io_out ? io_r_44_b : _GEN_2743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2745 = 8'h2d == r_count_12_io_out ? io_r_45_b : _GEN_2744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2746 = 8'h2e == r_count_12_io_out ? io_r_46_b : _GEN_2745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2747 = 8'h2f == r_count_12_io_out ? io_r_47_b : _GEN_2746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2748 = 8'h30 == r_count_12_io_out ? io_r_48_b : _GEN_2747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2749 = 8'h31 == r_count_12_io_out ? io_r_49_b : _GEN_2748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2750 = 8'h32 == r_count_12_io_out ? io_r_50_b : _GEN_2749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2751 = 8'h33 == r_count_12_io_out ? io_r_51_b : _GEN_2750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2752 = 8'h34 == r_count_12_io_out ? io_r_52_b : _GEN_2751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2753 = 8'h35 == r_count_12_io_out ? io_r_53_b : _GEN_2752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2754 = 8'h36 == r_count_12_io_out ? io_r_54_b : _GEN_2753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2755 = 8'h37 == r_count_12_io_out ? io_r_55_b : _GEN_2754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2756 = 8'h38 == r_count_12_io_out ? io_r_56_b : _GEN_2755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2757 = 8'h39 == r_count_12_io_out ? io_r_57_b : _GEN_2756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2758 = 8'h3a == r_count_12_io_out ? io_r_58_b : _GEN_2757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2759 = 8'h3b == r_count_12_io_out ? io_r_59_b : _GEN_2758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2760 = 8'h3c == r_count_12_io_out ? io_r_60_b : _GEN_2759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2761 = 8'h3d == r_count_12_io_out ? io_r_61_b : _GEN_2760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2762 = 8'h3e == r_count_12_io_out ? io_r_62_b : _GEN_2761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2763 = 8'h3f == r_count_12_io_out ? io_r_63_b : _GEN_2762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2764 = 8'h40 == r_count_12_io_out ? io_r_64_b : _GEN_2763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2765 = 8'h41 == r_count_12_io_out ? io_r_65_b : _GEN_2764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2766 = 8'h42 == r_count_12_io_out ? io_r_66_b : _GEN_2765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2767 = 8'h43 == r_count_12_io_out ? io_r_67_b : _GEN_2766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2768 = 8'h44 == r_count_12_io_out ? io_r_68_b : _GEN_2767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2769 = 8'h45 == r_count_12_io_out ? io_r_69_b : _GEN_2768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2770 = 8'h46 == r_count_12_io_out ? io_r_70_b : _GEN_2769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2771 = 8'h47 == r_count_12_io_out ? io_r_71_b : _GEN_2770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2772 = 8'h48 == r_count_12_io_out ? io_r_72_b : _GEN_2771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2773 = 8'h49 == r_count_12_io_out ? io_r_73_b : _GEN_2772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2774 = 8'h4a == r_count_12_io_out ? io_r_74_b : _GEN_2773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2775 = 8'h4b == r_count_12_io_out ? io_r_75_b : _GEN_2774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2776 = 8'h4c == r_count_12_io_out ? io_r_76_b : _GEN_2775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2777 = 8'h4d == r_count_12_io_out ? io_r_77_b : _GEN_2776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2778 = 8'h4e == r_count_12_io_out ? io_r_78_b : _GEN_2777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2779 = 8'h4f == r_count_12_io_out ? io_r_79_b : _GEN_2778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2780 = 8'h50 == r_count_12_io_out ? io_r_80_b : _GEN_2779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2781 = 8'h51 == r_count_12_io_out ? io_r_81_b : _GEN_2780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2782 = 8'h52 == r_count_12_io_out ? io_r_82_b : _GEN_2781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2783 = 8'h53 == r_count_12_io_out ? io_r_83_b : _GEN_2782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2784 = 8'h54 == r_count_12_io_out ? io_r_84_b : _GEN_2783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2785 = 8'h55 == r_count_12_io_out ? io_r_85_b : _GEN_2784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2786 = 8'h56 == r_count_12_io_out ? io_r_86_b : _GEN_2785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2787 = 8'h57 == r_count_12_io_out ? io_r_87_b : _GEN_2786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2788 = 8'h58 == r_count_12_io_out ? io_r_88_b : _GEN_2787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2789 = 8'h59 == r_count_12_io_out ? io_r_89_b : _GEN_2788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2790 = 8'h5a == r_count_12_io_out ? io_r_90_b : _GEN_2789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2791 = 8'h5b == r_count_12_io_out ? io_r_91_b : _GEN_2790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2792 = 8'h5c == r_count_12_io_out ? io_r_92_b : _GEN_2791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2793 = 8'h5d == r_count_12_io_out ? io_r_93_b : _GEN_2792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2794 = 8'h5e == r_count_12_io_out ? io_r_94_b : _GEN_2793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2795 = 8'h5f == r_count_12_io_out ? io_r_95_b : _GEN_2794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2796 = 8'h60 == r_count_12_io_out ? io_r_96_b : _GEN_2795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2797 = 8'h61 == r_count_12_io_out ? io_r_97_b : _GEN_2796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2798 = 8'h62 == r_count_12_io_out ? io_r_98_b : _GEN_2797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2799 = 8'h63 == r_count_12_io_out ? io_r_99_b : _GEN_2798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2800 = 8'h64 == r_count_12_io_out ? io_r_100_b : _GEN_2799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2801 = 8'h65 == r_count_12_io_out ? io_r_101_b : _GEN_2800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2802 = 8'h66 == r_count_12_io_out ? io_r_102_b : _GEN_2801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2803 = 8'h67 == r_count_12_io_out ? io_r_103_b : _GEN_2802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2804 = 8'h68 == r_count_12_io_out ? io_r_104_b : _GEN_2803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2805 = 8'h69 == r_count_12_io_out ? io_r_105_b : _GEN_2804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2806 = 8'h6a == r_count_12_io_out ? io_r_106_b : _GEN_2805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2807 = 8'h6b == r_count_12_io_out ? io_r_107_b : _GEN_2806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2808 = 8'h6c == r_count_12_io_out ? io_r_108_b : _GEN_2807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2809 = 8'h6d == r_count_12_io_out ? io_r_109_b : _GEN_2808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2810 = 8'h6e == r_count_12_io_out ? io_r_110_b : _GEN_2809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2811 = 8'h6f == r_count_12_io_out ? io_r_111_b : _GEN_2810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2812 = 8'h70 == r_count_12_io_out ? io_r_112_b : _GEN_2811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2813 = 8'h71 == r_count_12_io_out ? io_r_113_b : _GEN_2812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2814 = 8'h72 == r_count_12_io_out ? io_r_114_b : _GEN_2813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2815 = 8'h73 == r_count_12_io_out ? io_r_115_b : _GEN_2814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2816 = 8'h74 == r_count_12_io_out ? io_r_116_b : _GEN_2815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2817 = 8'h75 == r_count_12_io_out ? io_r_117_b : _GEN_2816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2818 = 8'h76 == r_count_12_io_out ? io_r_118_b : _GEN_2817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2819 = 8'h77 == r_count_12_io_out ? io_r_119_b : _GEN_2818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2820 = 8'h78 == r_count_12_io_out ? io_r_120_b : _GEN_2819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2821 = 8'h79 == r_count_12_io_out ? io_r_121_b : _GEN_2820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2822 = 8'h7a == r_count_12_io_out ? io_r_122_b : _GEN_2821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2823 = 8'h7b == r_count_12_io_out ? io_r_123_b : _GEN_2822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2824 = 8'h7c == r_count_12_io_out ? io_r_124_b : _GEN_2823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2825 = 8'h7d == r_count_12_io_out ? io_r_125_b : _GEN_2824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2826 = 8'h7e == r_count_12_io_out ? io_r_126_b : _GEN_2825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2827 = 8'h7f == r_count_12_io_out ? io_r_127_b : _GEN_2826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2828 = 8'h80 == r_count_12_io_out ? io_r_128_b : _GEN_2827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2829 = 8'h81 == r_count_12_io_out ? io_r_129_b : _GEN_2828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2830 = 8'h82 == r_count_12_io_out ? io_r_130_b : _GEN_2829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2831 = 8'h83 == r_count_12_io_out ? io_r_131_b : _GEN_2830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2832 = 8'h84 == r_count_12_io_out ? io_r_132_b : _GEN_2831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2833 = 8'h85 == r_count_12_io_out ? io_r_133_b : _GEN_2832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2834 = 8'h86 == r_count_12_io_out ? io_r_134_b : _GEN_2833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2835 = 8'h87 == r_count_12_io_out ? io_r_135_b : _GEN_2834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2836 = 8'h88 == r_count_12_io_out ? io_r_136_b : _GEN_2835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2837 = 8'h89 == r_count_12_io_out ? io_r_137_b : _GEN_2836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2838 = 8'h8a == r_count_12_io_out ? io_r_138_b : _GEN_2837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2839 = 8'h8b == r_count_12_io_out ? io_r_139_b : _GEN_2838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2840 = 8'h8c == r_count_12_io_out ? io_r_140_b : _GEN_2839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2841 = 8'h8d == r_count_12_io_out ? io_r_141_b : _GEN_2840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2842 = 8'h8e == r_count_12_io_out ? io_r_142_b : _GEN_2841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2843 = 8'h8f == r_count_12_io_out ? io_r_143_b : _GEN_2842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2844 = 8'h90 == r_count_12_io_out ? io_r_144_b : _GEN_2843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2845 = 8'h91 == r_count_12_io_out ? io_r_145_b : _GEN_2844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2846 = 8'h92 == r_count_12_io_out ? io_r_146_b : _GEN_2845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2847 = 8'h93 == r_count_12_io_out ? io_r_147_b : _GEN_2846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2848 = 8'h94 == r_count_12_io_out ? io_r_148_b : _GEN_2847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2849 = 8'h95 == r_count_12_io_out ? io_r_149_b : _GEN_2848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2850 = 8'h96 == r_count_12_io_out ? io_r_150_b : _GEN_2849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2851 = 8'h97 == r_count_12_io_out ? io_r_151_b : _GEN_2850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2852 = 8'h98 == r_count_12_io_out ? io_r_152_b : _GEN_2851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2853 = 8'h99 == r_count_12_io_out ? io_r_153_b : _GEN_2852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2854 = 8'h9a == r_count_12_io_out ? io_r_154_b : _GEN_2853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2855 = 8'h9b == r_count_12_io_out ? io_r_155_b : _GEN_2854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2856 = 8'h9c == r_count_12_io_out ? io_r_156_b : _GEN_2855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2857 = 8'h9d == r_count_12_io_out ? io_r_157_b : _GEN_2856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2858 = 8'h9e == r_count_12_io_out ? io_r_158_b : _GEN_2857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2859 = 8'h9f == r_count_12_io_out ? io_r_159_b : _GEN_2858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2860 = 8'ha0 == r_count_12_io_out ? io_r_160_b : _GEN_2859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2861 = 8'ha1 == r_count_12_io_out ? io_r_161_b : _GEN_2860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2862 = 8'ha2 == r_count_12_io_out ? io_r_162_b : _GEN_2861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2863 = 8'ha3 == r_count_12_io_out ? io_r_163_b : _GEN_2862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2864 = 8'ha4 == r_count_12_io_out ? io_r_164_b : _GEN_2863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2865 = 8'ha5 == r_count_12_io_out ? io_r_165_b : _GEN_2864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2866 = 8'ha6 == r_count_12_io_out ? io_r_166_b : _GEN_2865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2867 = 8'ha7 == r_count_12_io_out ? io_r_167_b : _GEN_2866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2868 = 8'ha8 == r_count_12_io_out ? io_r_168_b : _GEN_2867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2869 = 8'ha9 == r_count_12_io_out ? io_r_169_b : _GEN_2868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2870 = 8'haa == r_count_12_io_out ? io_r_170_b : _GEN_2869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2871 = 8'hab == r_count_12_io_out ? io_r_171_b : _GEN_2870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2872 = 8'hac == r_count_12_io_out ? io_r_172_b : _GEN_2871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2873 = 8'had == r_count_12_io_out ? io_r_173_b : _GEN_2872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2874 = 8'hae == r_count_12_io_out ? io_r_174_b : _GEN_2873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2875 = 8'haf == r_count_12_io_out ? io_r_175_b : _GEN_2874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2876 = 8'hb0 == r_count_12_io_out ? io_r_176_b : _GEN_2875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2877 = 8'hb1 == r_count_12_io_out ? io_r_177_b : _GEN_2876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2878 = 8'hb2 == r_count_12_io_out ? io_r_178_b : _GEN_2877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2879 = 8'hb3 == r_count_12_io_out ? io_r_179_b : _GEN_2878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2880 = 8'hb4 == r_count_12_io_out ? io_r_180_b : _GEN_2879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2881 = 8'hb5 == r_count_12_io_out ? io_r_181_b : _GEN_2880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2882 = 8'hb6 == r_count_12_io_out ? io_r_182_b : _GEN_2881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2883 = 8'hb7 == r_count_12_io_out ? io_r_183_b : _GEN_2882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2884 = 8'hb8 == r_count_12_io_out ? io_r_184_b : _GEN_2883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2885 = 8'hb9 == r_count_12_io_out ? io_r_185_b : _GEN_2884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2886 = 8'hba == r_count_12_io_out ? io_r_186_b : _GEN_2885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2887 = 8'hbb == r_count_12_io_out ? io_r_187_b : _GEN_2886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2888 = 8'hbc == r_count_12_io_out ? io_r_188_b : _GEN_2887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2889 = 8'hbd == r_count_12_io_out ? io_r_189_b : _GEN_2888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2890 = 8'hbe == r_count_12_io_out ? io_r_190_b : _GEN_2889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2891 = 8'hbf == r_count_12_io_out ? io_r_191_b : _GEN_2890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2892 = 8'hc0 == r_count_12_io_out ? io_r_192_b : _GEN_2891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2893 = 8'hc1 == r_count_12_io_out ? io_r_193_b : _GEN_2892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2894 = 8'hc2 == r_count_12_io_out ? io_r_194_b : _GEN_2893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2895 = 8'hc3 == r_count_12_io_out ? io_r_195_b : _GEN_2894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2896 = 8'hc4 == r_count_12_io_out ? io_r_196_b : _GEN_2895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2897 = 8'hc5 == r_count_12_io_out ? io_r_197_b : _GEN_2896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2898 = 8'hc6 == r_count_12_io_out ? io_r_198_b : _GEN_2897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2901 = 8'h1 == r_count_13_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2902 = 8'h2 == r_count_13_io_out ? io_r_2_b : _GEN_2901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2903 = 8'h3 == r_count_13_io_out ? io_r_3_b : _GEN_2902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2904 = 8'h4 == r_count_13_io_out ? io_r_4_b : _GEN_2903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2905 = 8'h5 == r_count_13_io_out ? io_r_5_b : _GEN_2904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2906 = 8'h6 == r_count_13_io_out ? io_r_6_b : _GEN_2905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2907 = 8'h7 == r_count_13_io_out ? io_r_7_b : _GEN_2906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2908 = 8'h8 == r_count_13_io_out ? io_r_8_b : _GEN_2907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2909 = 8'h9 == r_count_13_io_out ? io_r_9_b : _GEN_2908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2910 = 8'ha == r_count_13_io_out ? io_r_10_b : _GEN_2909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2911 = 8'hb == r_count_13_io_out ? io_r_11_b : _GEN_2910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2912 = 8'hc == r_count_13_io_out ? io_r_12_b : _GEN_2911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2913 = 8'hd == r_count_13_io_out ? io_r_13_b : _GEN_2912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2914 = 8'he == r_count_13_io_out ? io_r_14_b : _GEN_2913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2915 = 8'hf == r_count_13_io_out ? io_r_15_b : _GEN_2914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2916 = 8'h10 == r_count_13_io_out ? io_r_16_b : _GEN_2915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2917 = 8'h11 == r_count_13_io_out ? io_r_17_b : _GEN_2916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2918 = 8'h12 == r_count_13_io_out ? io_r_18_b : _GEN_2917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2919 = 8'h13 == r_count_13_io_out ? io_r_19_b : _GEN_2918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2920 = 8'h14 == r_count_13_io_out ? io_r_20_b : _GEN_2919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2921 = 8'h15 == r_count_13_io_out ? io_r_21_b : _GEN_2920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2922 = 8'h16 == r_count_13_io_out ? io_r_22_b : _GEN_2921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2923 = 8'h17 == r_count_13_io_out ? io_r_23_b : _GEN_2922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2924 = 8'h18 == r_count_13_io_out ? io_r_24_b : _GEN_2923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2925 = 8'h19 == r_count_13_io_out ? io_r_25_b : _GEN_2924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2926 = 8'h1a == r_count_13_io_out ? io_r_26_b : _GEN_2925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2927 = 8'h1b == r_count_13_io_out ? io_r_27_b : _GEN_2926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2928 = 8'h1c == r_count_13_io_out ? io_r_28_b : _GEN_2927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2929 = 8'h1d == r_count_13_io_out ? io_r_29_b : _GEN_2928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2930 = 8'h1e == r_count_13_io_out ? io_r_30_b : _GEN_2929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2931 = 8'h1f == r_count_13_io_out ? io_r_31_b : _GEN_2930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2932 = 8'h20 == r_count_13_io_out ? io_r_32_b : _GEN_2931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2933 = 8'h21 == r_count_13_io_out ? io_r_33_b : _GEN_2932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2934 = 8'h22 == r_count_13_io_out ? io_r_34_b : _GEN_2933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2935 = 8'h23 == r_count_13_io_out ? io_r_35_b : _GEN_2934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2936 = 8'h24 == r_count_13_io_out ? io_r_36_b : _GEN_2935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2937 = 8'h25 == r_count_13_io_out ? io_r_37_b : _GEN_2936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2938 = 8'h26 == r_count_13_io_out ? io_r_38_b : _GEN_2937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2939 = 8'h27 == r_count_13_io_out ? io_r_39_b : _GEN_2938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2940 = 8'h28 == r_count_13_io_out ? io_r_40_b : _GEN_2939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2941 = 8'h29 == r_count_13_io_out ? io_r_41_b : _GEN_2940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2942 = 8'h2a == r_count_13_io_out ? io_r_42_b : _GEN_2941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2943 = 8'h2b == r_count_13_io_out ? io_r_43_b : _GEN_2942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2944 = 8'h2c == r_count_13_io_out ? io_r_44_b : _GEN_2943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2945 = 8'h2d == r_count_13_io_out ? io_r_45_b : _GEN_2944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2946 = 8'h2e == r_count_13_io_out ? io_r_46_b : _GEN_2945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2947 = 8'h2f == r_count_13_io_out ? io_r_47_b : _GEN_2946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2948 = 8'h30 == r_count_13_io_out ? io_r_48_b : _GEN_2947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2949 = 8'h31 == r_count_13_io_out ? io_r_49_b : _GEN_2948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2950 = 8'h32 == r_count_13_io_out ? io_r_50_b : _GEN_2949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2951 = 8'h33 == r_count_13_io_out ? io_r_51_b : _GEN_2950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2952 = 8'h34 == r_count_13_io_out ? io_r_52_b : _GEN_2951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2953 = 8'h35 == r_count_13_io_out ? io_r_53_b : _GEN_2952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2954 = 8'h36 == r_count_13_io_out ? io_r_54_b : _GEN_2953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2955 = 8'h37 == r_count_13_io_out ? io_r_55_b : _GEN_2954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2956 = 8'h38 == r_count_13_io_out ? io_r_56_b : _GEN_2955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2957 = 8'h39 == r_count_13_io_out ? io_r_57_b : _GEN_2956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2958 = 8'h3a == r_count_13_io_out ? io_r_58_b : _GEN_2957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2959 = 8'h3b == r_count_13_io_out ? io_r_59_b : _GEN_2958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2960 = 8'h3c == r_count_13_io_out ? io_r_60_b : _GEN_2959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2961 = 8'h3d == r_count_13_io_out ? io_r_61_b : _GEN_2960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2962 = 8'h3e == r_count_13_io_out ? io_r_62_b : _GEN_2961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2963 = 8'h3f == r_count_13_io_out ? io_r_63_b : _GEN_2962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2964 = 8'h40 == r_count_13_io_out ? io_r_64_b : _GEN_2963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2965 = 8'h41 == r_count_13_io_out ? io_r_65_b : _GEN_2964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2966 = 8'h42 == r_count_13_io_out ? io_r_66_b : _GEN_2965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2967 = 8'h43 == r_count_13_io_out ? io_r_67_b : _GEN_2966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2968 = 8'h44 == r_count_13_io_out ? io_r_68_b : _GEN_2967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2969 = 8'h45 == r_count_13_io_out ? io_r_69_b : _GEN_2968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2970 = 8'h46 == r_count_13_io_out ? io_r_70_b : _GEN_2969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2971 = 8'h47 == r_count_13_io_out ? io_r_71_b : _GEN_2970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2972 = 8'h48 == r_count_13_io_out ? io_r_72_b : _GEN_2971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2973 = 8'h49 == r_count_13_io_out ? io_r_73_b : _GEN_2972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2974 = 8'h4a == r_count_13_io_out ? io_r_74_b : _GEN_2973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2975 = 8'h4b == r_count_13_io_out ? io_r_75_b : _GEN_2974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2976 = 8'h4c == r_count_13_io_out ? io_r_76_b : _GEN_2975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2977 = 8'h4d == r_count_13_io_out ? io_r_77_b : _GEN_2976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2978 = 8'h4e == r_count_13_io_out ? io_r_78_b : _GEN_2977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2979 = 8'h4f == r_count_13_io_out ? io_r_79_b : _GEN_2978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2980 = 8'h50 == r_count_13_io_out ? io_r_80_b : _GEN_2979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2981 = 8'h51 == r_count_13_io_out ? io_r_81_b : _GEN_2980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2982 = 8'h52 == r_count_13_io_out ? io_r_82_b : _GEN_2981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2983 = 8'h53 == r_count_13_io_out ? io_r_83_b : _GEN_2982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2984 = 8'h54 == r_count_13_io_out ? io_r_84_b : _GEN_2983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2985 = 8'h55 == r_count_13_io_out ? io_r_85_b : _GEN_2984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2986 = 8'h56 == r_count_13_io_out ? io_r_86_b : _GEN_2985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2987 = 8'h57 == r_count_13_io_out ? io_r_87_b : _GEN_2986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2988 = 8'h58 == r_count_13_io_out ? io_r_88_b : _GEN_2987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2989 = 8'h59 == r_count_13_io_out ? io_r_89_b : _GEN_2988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2990 = 8'h5a == r_count_13_io_out ? io_r_90_b : _GEN_2989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2991 = 8'h5b == r_count_13_io_out ? io_r_91_b : _GEN_2990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2992 = 8'h5c == r_count_13_io_out ? io_r_92_b : _GEN_2991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2993 = 8'h5d == r_count_13_io_out ? io_r_93_b : _GEN_2992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2994 = 8'h5e == r_count_13_io_out ? io_r_94_b : _GEN_2993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2995 = 8'h5f == r_count_13_io_out ? io_r_95_b : _GEN_2994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2996 = 8'h60 == r_count_13_io_out ? io_r_96_b : _GEN_2995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2997 = 8'h61 == r_count_13_io_out ? io_r_97_b : _GEN_2996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2998 = 8'h62 == r_count_13_io_out ? io_r_98_b : _GEN_2997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2999 = 8'h63 == r_count_13_io_out ? io_r_99_b : _GEN_2998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3000 = 8'h64 == r_count_13_io_out ? io_r_100_b : _GEN_2999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3001 = 8'h65 == r_count_13_io_out ? io_r_101_b : _GEN_3000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3002 = 8'h66 == r_count_13_io_out ? io_r_102_b : _GEN_3001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3003 = 8'h67 == r_count_13_io_out ? io_r_103_b : _GEN_3002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3004 = 8'h68 == r_count_13_io_out ? io_r_104_b : _GEN_3003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3005 = 8'h69 == r_count_13_io_out ? io_r_105_b : _GEN_3004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3006 = 8'h6a == r_count_13_io_out ? io_r_106_b : _GEN_3005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3007 = 8'h6b == r_count_13_io_out ? io_r_107_b : _GEN_3006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3008 = 8'h6c == r_count_13_io_out ? io_r_108_b : _GEN_3007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3009 = 8'h6d == r_count_13_io_out ? io_r_109_b : _GEN_3008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3010 = 8'h6e == r_count_13_io_out ? io_r_110_b : _GEN_3009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3011 = 8'h6f == r_count_13_io_out ? io_r_111_b : _GEN_3010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3012 = 8'h70 == r_count_13_io_out ? io_r_112_b : _GEN_3011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3013 = 8'h71 == r_count_13_io_out ? io_r_113_b : _GEN_3012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3014 = 8'h72 == r_count_13_io_out ? io_r_114_b : _GEN_3013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3015 = 8'h73 == r_count_13_io_out ? io_r_115_b : _GEN_3014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3016 = 8'h74 == r_count_13_io_out ? io_r_116_b : _GEN_3015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3017 = 8'h75 == r_count_13_io_out ? io_r_117_b : _GEN_3016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3018 = 8'h76 == r_count_13_io_out ? io_r_118_b : _GEN_3017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3019 = 8'h77 == r_count_13_io_out ? io_r_119_b : _GEN_3018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3020 = 8'h78 == r_count_13_io_out ? io_r_120_b : _GEN_3019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3021 = 8'h79 == r_count_13_io_out ? io_r_121_b : _GEN_3020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3022 = 8'h7a == r_count_13_io_out ? io_r_122_b : _GEN_3021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3023 = 8'h7b == r_count_13_io_out ? io_r_123_b : _GEN_3022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3024 = 8'h7c == r_count_13_io_out ? io_r_124_b : _GEN_3023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3025 = 8'h7d == r_count_13_io_out ? io_r_125_b : _GEN_3024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3026 = 8'h7e == r_count_13_io_out ? io_r_126_b : _GEN_3025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3027 = 8'h7f == r_count_13_io_out ? io_r_127_b : _GEN_3026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3028 = 8'h80 == r_count_13_io_out ? io_r_128_b : _GEN_3027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3029 = 8'h81 == r_count_13_io_out ? io_r_129_b : _GEN_3028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3030 = 8'h82 == r_count_13_io_out ? io_r_130_b : _GEN_3029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3031 = 8'h83 == r_count_13_io_out ? io_r_131_b : _GEN_3030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3032 = 8'h84 == r_count_13_io_out ? io_r_132_b : _GEN_3031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3033 = 8'h85 == r_count_13_io_out ? io_r_133_b : _GEN_3032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3034 = 8'h86 == r_count_13_io_out ? io_r_134_b : _GEN_3033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3035 = 8'h87 == r_count_13_io_out ? io_r_135_b : _GEN_3034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3036 = 8'h88 == r_count_13_io_out ? io_r_136_b : _GEN_3035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3037 = 8'h89 == r_count_13_io_out ? io_r_137_b : _GEN_3036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3038 = 8'h8a == r_count_13_io_out ? io_r_138_b : _GEN_3037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3039 = 8'h8b == r_count_13_io_out ? io_r_139_b : _GEN_3038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3040 = 8'h8c == r_count_13_io_out ? io_r_140_b : _GEN_3039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3041 = 8'h8d == r_count_13_io_out ? io_r_141_b : _GEN_3040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3042 = 8'h8e == r_count_13_io_out ? io_r_142_b : _GEN_3041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3043 = 8'h8f == r_count_13_io_out ? io_r_143_b : _GEN_3042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3044 = 8'h90 == r_count_13_io_out ? io_r_144_b : _GEN_3043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3045 = 8'h91 == r_count_13_io_out ? io_r_145_b : _GEN_3044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3046 = 8'h92 == r_count_13_io_out ? io_r_146_b : _GEN_3045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3047 = 8'h93 == r_count_13_io_out ? io_r_147_b : _GEN_3046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3048 = 8'h94 == r_count_13_io_out ? io_r_148_b : _GEN_3047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3049 = 8'h95 == r_count_13_io_out ? io_r_149_b : _GEN_3048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3050 = 8'h96 == r_count_13_io_out ? io_r_150_b : _GEN_3049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3051 = 8'h97 == r_count_13_io_out ? io_r_151_b : _GEN_3050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3052 = 8'h98 == r_count_13_io_out ? io_r_152_b : _GEN_3051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3053 = 8'h99 == r_count_13_io_out ? io_r_153_b : _GEN_3052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3054 = 8'h9a == r_count_13_io_out ? io_r_154_b : _GEN_3053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3055 = 8'h9b == r_count_13_io_out ? io_r_155_b : _GEN_3054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3056 = 8'h9c == r_count_13_io_out ? io_r_156_b : _GEN_3055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3057 = 8'h9d == r_count_13_io_out ? io_r_157_b : _GEN_3056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3058 = 8'h9e == r_count_13_io_out ? io_r_158_b : _GEN_3057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3059 = 8'h9f == r_count_13_io_out ? io_r_159_b : _GEN_3058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3060 = 8'ha0 == r_count_13_io_out ? io_r_160_b : _GEN_3059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3061 = 8'ha1 == r_count_13_io_out ? io_r_161_b : _GEN_3060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3062 = 8'ha2 == r_count_13_io_out ? io_r_162_b : _GEN_3061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3063 = 8'ha3 == r_count_13_io_out ? io_r_163_b : _GEN_3062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3064 = 8'ha4 == r_count_13_io_out ? io_r_164_b : _GEN_3063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3065 = 8'ha5 == r_count_13_io_out ? io_r_165_b : _GEN_3064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3066 = 8'ha6 == r_count_13_io_out ? io_r_166_b : _GEN_3065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3067 = 8'ha7 == r_count_13_io_out ? io_r_167_b : _GEN_3066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3068 = 8'ha8 == r_count_13_io_out ? io_r_168_b : _GEN_3067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3069 = 8'ha9 == r_count_13_io_out ? io_r_169_b : _GEN_3068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3070 = 8'haa == r_count_13_io_out ? io_r_170_b : _GEN_3069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3071 = 8'hab == r_count_13_io_out ? io_r_171_b : _GEN_3070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3072 = 8'hac == r_count_13_io_out ? io_r_172_b : _GEN_3071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3073 = 8'had == r_count_13_io_out ? io_r_173_b : _GEN_3072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3074 = 8'hae == r_count_13_io_out ? io_r_174_b : _GEN_3073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3075 = 8'haf == r_count_13_io_out ? io_r_175_b : _GEN_3074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3076 = 8'hb0 == r_count_13_io_out ? io_r_176_b : _GEN_3075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3077 = 8'hb1 == r_count_13_io_out ? io_r_177_b : _GEN_3076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3078 = 8'hb2 == r_count_13_io_out ? io_r_178_b : _GEN_3077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3079 = 8'hb3 == r_count_13_io_out ? io_r_179_b : _GEN_3078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3080 = 8'hb4 == r_count_13_io_out ? io_r_180_b : _GEN_3079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3081 = 8'hb5 == r_count_13_io_out ? io_r_181_b : _GEN_3080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3082 = 8'hb6 == r_count_13_io_out ? io_r_182_b : _GEN_3081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3083 = 8'hb7 == r_count_13_io_out ? io_r_183_b : _GEN_3082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3084 = 8'hb8 == r_count_13_io_out ? io_r_184_b : _GEN_3083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3085 = 8'hb9 == r_count_13_io_out ? io_r_185_b : _GEN_3084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3086 = 8'hba == r_count_13_io_out ? io_r_186_b : _GEN_3085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3087 = 8'hbb == r_count_13_io_out ? io_r_187_b : _GEN_3086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3088 = 8'hbc == r_count_13_io_out ? io_r_188_b : _GEN_3087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3089 = 8'hbd == r_count_13_io_out ? io_r_189_b : _GEN_3088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3090 = 8'hbe == r_count_13_io_out ? io_r_190_b : _GEN_3089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3091 = 8'hbf == r_count_13_io_out ? io_r_191_b : _GEN_3090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3092 = 8'hc0 == r_count_13_io_out ? io_r_192_b : _GEN_3091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3093 = 8'hc1 == r_count_13_io_out ? io_r_193_b : _GEN_3092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3094 = 8'hc2 == r_count_13_io_out ? io_r_194_b : _GEN_3093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3095 = 8'hc3 == r_count_13_io_out ? io_r_195_b : _GEN_3094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3096 = 8'hc4 == r_count_13_io_out ? io_r_196_b : _GEN_3095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3097 = 8'hc5 == r_count_13_io_out ? io_r_197_b : _GEN_3096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3098 = 8'hc6 == r_count_13_io_out ? io_r_198_b : _GEN_3097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3101 = 8'h1 == r_count_14_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3102 = 8'h2 == r_count_14_io_out ? io_r_2_b : _GEN_3101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3103 = 8'h3 == r_count_14_io_out ? io_r_3_b : _GEN_3102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3104 = 8'h4 == r_count_14_io_out ? io_r_4_b : _GEN_3103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3105 = 8'h5 == r_count_14_io_out ? io_r_5_b : _GEN_3104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3106 = 8'h6 == r_count_14_io_out ? io_r_6_b : _GEN_3105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3107 = 8'h7 == r_count_14_io_out ? io_r_7_b : _GEN_3106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3108 = 8'h8 == r_count_14_io_out ? io_r_8_b : _GEN_3107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3109 = 8'h9 == r_count_14_io_out ? io_r_9_b : _GEN_3108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3110 = 8'ha == r_count_14_io_out ? io_r_10_b : _GEN_3109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3111 = 8'hb == r_count_14_io_out ? io_r_11_b : _GEN_3110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3112 = 8'hc == r_count_14_io_out ? io_r_12_b : _GEN_3111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3113 = 8'hd == r_count_14_io_out ? io_r_13_b : _GEN_3112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3114 = 8'he == r_count_14_io_out ? io_r_14_b : _GEN_3113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3115 = 8'hf == r_count_14_io_out ? io_r_15_b : _GEN_3114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3116 = 8'h10 == r_count_14_io_out ? io_r_16_b : _GEN_3115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3117 = 8'h11 == r_count_14_io_out ? io_r_17_b : _GEN_3116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3118 = 8'h12 == r_count_14_io_out ? io_r_18_b : _GEN_3117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3119 = 8'h13 == r_count_14_io_out ? io_r_19_b : _GEN_3118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3120 = 8'h14 == r_count_14_io_out ? io_r_20_b : _GEN_3119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3121 = 8'h15 == r_count_14_io_out ? io_r_21_b : _GEN_3120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3122 = 8'h16 == r_count_14_io_out ? io_r_22_b : _GEN_3121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3123 = 8'h17 == r_count_14_io_out ? io_r_23_b : _GEN_3122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3124 = 8'h18 == r_count_14_io_out ? io_r_24_b : _GEN_3123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3125 = 8'h19 == r_count_14_io_out ? io_r_25_b : _GEN_3124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3126 = 8'h1a == r_count_14_io_out ? io_r_26_b : _GEN_3125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3127 = 8'h1b == r_count_14_io_out ? io_r_27_b : _GEN_3126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3128 = 8'h1c == r_count_14_io_out ? io_r_28_b : _GEN_3127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3129 = 8'h1d == r_count_14_io_out ? io_r_29_b : _GEN_3128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3130 = 8'h1e == r_count_14_io_out ? io_r_30_b : _GEN_3129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3131 = 8'h1f == r_count_14_io_out ? io_r_31_b : _GEN_3130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3132 = 8'h20 == r_count_14_io_out ? io_r_32_b : _GEN_3131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3133 = 8'h21 == r_count_14_io_out ? io_r_33_b : _GEN_3132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3134 = 8'h22 == r_count_14_io_out ? io_r_34_b : _GEN_3133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3135 = 8'h23 == r_count_14_io_out ? io_r_35_b : _GEN_3134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3136 = 8'h24 == r_count_14_io_out ? io_r_36_b : _GEN_3135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3137 = 8'h25 == r_count_14_io_out ? io_r_37_b : _GEN_3136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3138 = 8'h26 == r_count_14_io_out ? io_r_38_b : _GEN_3137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3139 = 8'h27 == r_count_14_io_out ? io_r_39_b : _GEN_3138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3140 = 8'h28 == r_count_14_io_out ? io_r_40_b : _GEN_3139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3141 = 8'h29 == r_count_14_io_out ? io_r_41_b : _GEN_3140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3142 = 8'h2a == r_count_14_io_out ? io_r_42_b : _GEN_3141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3143 = 8'h2b == r_count_14_io_out ? io_r_43_b : _GEN_3142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3144 = 8'h2c == r_count_14_io_out ? io_r_44_b : _GEN_3143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3145 = 8'h2d == r_count_14_io_out ? io_r_45_b : _GEN_3144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3146 = 8'h2e == r_count_14_io_out ? io_r_46_b : _GEN_3145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3147 = 8'h2f == r_count_14_io_out ? io_r_47_b : _GEN_3146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3148 = 8'h30 == r_count_14_io_out ? io_r_48_b : _GEN_3147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3149 = 8'h31 == r_count_14_io_out ? io_r_49_b : _GEN_3148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3150 = 8'h32 == r_count_14_io_out ? io_r_50_b : _GEN_3149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3151 = 8'h33 == r_count_14_io_out ? io_r_51_b : _GEN_3150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3152 = 8'h34 == r_count_14_io_out ? io_r_52_b : _GEN_3151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3153 = 8'h35 == r_count_14_io_out ? io_r_53_b : _GEN_3152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3154 = 8'h36 == r_count_14_io_out ? io_r_54_b : _GEN_3153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3155 = 8'h37 == r_count_14_io_out ? io_r_55_b : _GEN_3154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3156 = 8'h38 == r_count_14_io_out ? io_r_56_b : _GEN_3155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3157 = 8'h39 == r_count_14_io_out ? io_r_57_b : _GEN_3156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3158 = 8'h3a == r_count_14_io_out ? io_r_58_b : _GEN_3157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3159 = 8'h3b == r_count_14_io_out ? io_r_59_b : _GEN_3158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3160 = 8'h3c == r_count_14_io_out ? io_r_60_b : _GEN_3159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3161 = 8'h3d == r_count_14_io_out ? io_r_61_b : _GEN_3160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3162 = 8'h3e == r_count_14_io_out ? io_r_62_b : _GEN_3161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3163 = 8'h3f == r_count_14_io_out ? io_r_63_b : _GEN_3162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3164 = 8'h40 == r_count_14_io_out ? io_r_64_b : _GEN_3163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3165 = 8'h41 == r_count_14_io_out ? io_r_65_b : _GEN_3164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3166 = 8'h42 == r_count_14_io_out ? io_r_66_b : _GEN_3165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3167 = 8'h43 == r_count_14_io_out ? io_r_67_b : _GEN_3166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3168 = 8'h44 == r_count_14_io_out ? io_r_68_b : _GEN_3167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3169 = 8'h45 == r_count_14_io_out ? io_r_69_b : _GEN_3168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3170 = 8'h46 == r_count_14_io_out ? io_r_70_b : _GEN_3169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3171 = 8'h47 == r_count_14_io_out ? io_r_71_b : _GEN_3170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3172 = 8'h48 == r_count_14_io_out ? io_r_72_b : _GEN_3171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3173 = 8'h49 == r_count_14_io_out ? io_r_73_b : _GEN_3172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3174 = 8'h4a == r_count_14_io_out ? io_r_74_b : _GEN_3173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3175 = 8'h4b == r_count_14_io_out ? io_r_75_b : _GEN_3174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3176 = 8'h4c == r_count_14_io_out ? io_r_76_b : _GEN_3175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3177 = 8'h4d == r_count_14_io_out ? io_r_77_b : _GEN_3176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3178 = 8'h4e == r_count_14_io_out ? io_r_78_b : _GEN_3177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3179 = 8'h4f == r_count_14_io_out ? io_r_79_b : _GEN_3178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3180 = 8'h50 == r_count_14_io_out ? io_r_80_b : _GEN_3179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3181 = 8'h51 == r_count_14_io_out ? io_r_81_b : _GEN_3180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3182 = 8'h52 == r_count_14_io_out ? io_r_82_b : _GEN_3181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3183 = 8'h53 == r_count_14_io_out ? io_r_83_b : _GEN_3182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3184 = 8'h54 == r_count_14_io_out ? io_r_84_b : _GEN_3183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3185 = 8'h55 == r_count_14_io_out ? io_r_85_b : _GEN_3184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3186 = 8'h56 == r_count_14_io_out ? io_r_86_b : _GEN_3185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3187 = 8'h57 == r_count_14_io_out ? io_r_87_b : _GEN_3186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3188 = 8'h58 == r_count_14_io_out ? io_r_88_b : _GEN_3187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3189 = 8'h59 == r_count_14_io_out ? io_r_89_b : _GEN_3188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3190 = 8'h5a == r_count_14_io_out ? io_r_90_b : _GEN_3189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3191 = 8'h5b == r_count_14_io_out ? io_r_91_b : _GEN_3190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3192 = 8'h5c == r_count_14_io_out ? io_r_92_b : _GEN_3191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3193 = 8'h5d == r_count_14_io_out ? io_r_93_b : _GEN_3192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3194 = 8'h5e == r_count_14_io_out ? io_r_94_b : _GEN_3193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3195 = 8'h5f == r_count_14_io_out ? io_r_95_b : _GEN_3194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3196 = 8'h60 == r_count_14_io_out ? io_r_96_b : _GEN_3195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3197 = 8'h61 == r_count_14_io_out ? io_r_97_b : _GEN_3196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3198 = 8'h62 == r_count_14_io_out ? io_r_98_b : _GEN_3197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3199 = 8'h63 == r_count_14_io_out ? io_r_99_b : _GEN_3198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3200 = 8'h64 == r_count_14_io_out ? io_r_100_b : _GEN_3199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3201 = 8'h65 == r_count_14_io_out ? io_r_101_b : _GEN_3200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3202 = 8'h66 == r_count_14_io_out ? io_r_102_b : _GEN_3201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3203 = 8'h67 == r_count_14_io_out ? io_r_103_b : _GEN_3202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3204 = 8'h68 == r_count_14_io_out ? io_r_104_b : _GEN_3203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3205 = 8'h69 == r_count_14_io_out ? io_r_105_b : _GEN_3204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3206 = 8'h6a == r_count_14_io_out ? io_r_106_b : _GEN_3205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3207 = 8'h6b == r_count_14_io_out ? io_r_107_b : _GEN_3206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3208 = 8'h6c == r_count_14_io_out ? io_r_108_b : _GEN_3207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3209 = 8'h6d == r_count_14_io_out ? io_r_109_b : _GEN_3208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3210 = 8'h6e == r_count_14_io_out ? io_r_110_b : _GEN_3209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3211 = 8'h6f == r_count_14_io_out ? io_r_111_b : _GEN_3210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3212 = 8'h70 == r_count_14_io_out ? io_r_112_b : _GEN_3211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3213 = 8'h71 == r_count_14_io_out ? io_r_113_b : _GEN_3212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3214 = 8'h72 == r_count_14_io_out ? io_r_114_b : _GEN_3213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3215 = 8'h73 == r_count_14_io_out ? io_r_115_b : _GEN_3214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3216 = 8'h74 == r_count_14_io_out ? io_r_116_b : _GEN_3215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3217 = 8'h75 == r_count_14_io_out ? io_r_117_b : _GEN_3216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3218 = 8'h76 == r_count_14_io_out ? io_r_118_b : _GEN_3217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3219 = 8'h77 == r_count_14_io_out ? io_r_119_b : _GEN_3218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3220 = 8'h78 == r_count_14_io_out ? io_r_120_b : _GEN_3219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3221 = 8'h79 == r_count_14_io_out ? io_r_121_b : _GEN_3220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3222 = 8'h7a == r_count_14_io_out ? io_r_122_b : _GEN_3221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3223 = 8'h7b == r_count_14_io_out ? io_r_123_b : _GEN_3222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3224 = 8'h7c == r_count_14_io_out ? io_r_124_b : _GEN_3223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3225 = 8'h7d == r_count_14_io_out ? io_r_125_b : _GEN_3224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3226 = 8'h7e == r_count_14_io_out ? io_r_126_b : _GEN_3225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3227 = 8'h7f == r_count_14_io_out ? io_r_127_b : _GEN_3226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3228 = 8'h80 == r_count_14_io_out ? io_r_128_b : _GEN_3227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3229 = 8'h81 == r_count_14_io_out ? io_r_129_b : _GEN_3228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3230 = 8'h82 == r_count_14_io_out ? io_r_130_b : _GEN_3229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3231 = 8'h83 == r_count_14_io_out ? io_r_131_b : _GEN_3230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3232 = 8'h84 == r_count_14_io_out ? io_r_132_b : _GEN_3231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3233 = 8'h85 == r_count_14_io_out ? io_r_133_b : _GEN_3232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3234 = 8'h86 == r_count_14_io_out ? io_r_134_b : _GEN_3233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3235 = 8'h87 == r_count_14_io_out ? io_r_135_b : _GEN_3234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3236 = 8'h88 == r_count_14_io_out ? io_r_136_b : _GEN_3235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3237 = 8'h89 == r_count_14_io_out ? io_r_137_b : _GEN_3236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3238 = 8'h8a == r_count_14_io_out ? io_r_138_b : _GEN_3237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3239 = 8'h8b == r_count_14_io_out ? io_r_139_b : _GEN_3238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3240 = 8'h8c == r_count_14_io_out ? io_r_140_b : _GEN_3239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3241 = 8'h8d == r_count_14_io_out ? io_r_141_b : _GEN_3240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3242 = 8'h8e == r_count_14_io_out ? io_r_142_b : _GEN_3241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3243 = 8'h8f == r_count_14_io_out ? io_r_143_b : _GEN_3242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3244 = 8'h90 == r_count_14_io_out ? io_r_144_b : _GEN_3243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3245 = 8'h91 == r_count_14_io_out ? io_r_145_b : _GEN_3244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3246 = 8'h92 == r_count_14_io_out ? io_r_146_b : _GEN_3245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3247 = 8'h93 == r_count_14_io_out ? io_r_147_b : _GEN_3246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3248 = 8'h94 == r_count_14_io_out ? io_r_148_b : _GEN_3247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3249 = 8'h95 == r_count_14_io_out ? io_r_149_b : _GEN_3248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3250 = 8'h96 == r_count_14_io_out ? io_r_150_b : _GEN_3249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3251 = 8'h97 == r_count_14_io_out ? io_r_151_b : _GEN_3250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3252 = 8'h98 == r_count_14_io_out ? io_r_152_b : _GEN_3251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3253 = 8'h99 == r_count_14_io_out ? io_r_153_b : _GEN_3252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3254 = 8'h9a == r_count_14_io_out ? io_r_154_b : _GEN_3253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3255 = 8'h9b == r_count_14_io_out ? io_r_155_b : _GEN_3254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3256 = 8'h9c == r_count_14_io_out ? io_r_156_b : _GEN_3255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3257 = 8'h9d == r_count_14_io_out ? io_r_157_b : _GEN_3256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3258 = 8'h9e == r_count_14_io_out ? io_r_158_b : _GEN_3257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3259 = 8'h9f == r_count_14_io_out ? io_r_159_b : _GEN_3258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3260 = 8'ha0 == r_count_14_io_out ? io_r_160_b : _GEN_3259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3261 = 8'ha1 == r_count_14_io_out ? io_r_161_b : _GEN_3260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3262 = 8'ha2 == r_count_14_io_out ? io_r_162_b : _GEN_3261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3263 = 8'ha3 == r_count_14_io_out ? io_r_163_b : _GEN_3262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3264 = 8'ha4 == r_count_14_io_out ? io_r_164_b : _GEN_3263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3265 = 8'ha5 == r_count_14_io_out ? io_r_165_b : _GEN_3264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3266 = 8'ha6 == r_count_14_io_out ? io_r_166_b : _GEN_3265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3267 = 8'ha7 == r_count_14_io_out ? io_r_167_b : _GEN_3266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3268 = 8'ha8 == r_count_14_io_out ? io_r_168_b : _GEN_3267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3269 = 8'ha9 == r_count_14_io_out ? io_r_169_b : _GEN_3268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3270 = 8'haa == r_count_14_io_out ? io_r_170_b : _GEN_3269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3271 = 8'hab == r_count_14_io_out ? io_r_171_b : _GEN_3270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3272 = 8'hac == r_count_14_io_out ? io_r_172_b : _GEN_3271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3273 = 8'had == r_count_14_io_out ? io_r_173_b : _GEN_3272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3274 = 8'hae == r_count_14_io_out ? io_r_174_b : _GEN_3273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3275 = 8'haf == r_count_14_io_out ? io_r_175_b : _GEN_3274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3276 = 8'hb0 == r_count_14_io_out ? io_r_176_b : _GEN_3275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3277 = 8'hb1 == r_count_14_io_out ? io_r_177_b : _GEN_3276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3278 = 8'hb2 == r_count_14_io_out ? io_r_178_b : _GEN_3277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3279 = 8'hb3 == r_count_14_io_out ? io_r_179_b : _GEN_3278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3280 = 8'hb4 == r_count_14_io_out ? io_r_180_b : _GEN_3279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3281 = 8'hb5 == r_count_14_io_out ? io_r_181_b : _GEN_3280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3282 = 8'hb6 == r_count_14_io_out ? io_r_182_b : _GEN_3281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3283 = 8'hb7 == r_count_14_io_out ? io_r_183_b : _GEN_3282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3284 = 8'hb8 == r_count_14_io_out ? io_r_184_b : _GEN_3283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3285 = 8'hb9 == r_count_14_io_out ? io_r_185_b : _GEN_3284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3286 = 8'hba == r_count_14_io_out ? io_r_186_b : _GEN_3285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3287 = 8'hbb == r_count_14_io_out ? io_r_187_b : _GEN_3286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3288 = 8'hbc == r_count_14_io_out ? io_r_188_b : _GEN_3287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3289 = 8'hbd == r_count_14_io_out ? io_r_189_b : _GEN_3288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3290 = 8'hbe == r_count_14_io_out ? io_r_190_b : _GEN_3289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3291 = 8'hbf == r_count_14_io_out ? io_r_191_b : _GEN_3290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3292 = 8'hc0 == r_count_14_io_out ? io_r_192_b : _GEN_3291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3293 = 8'hc1 == r_count_14_io_out ? io_r_193_b : _GEN_3292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3294 = 8'hc2 == r_count_14_io_out ? io_r_194_b : _GEN_3293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3295 = 8'hc3 == r_count_14_io_out ? io_r_195_b : _GEN_3294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3296 = 8'hc4 == r_count_14_io_out ? io_r_196_b : _GEN_3295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3297 = 8'hc5 == r_count_14_io_out ? io_r_197_b : _GEN_3296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3298 = 8'hc6 == r_count_14_io_out ? io_r_198_b : _GEN_3297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3301 = 8'h1 == r_count_15_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3302 = 8'h2 == r_count_15_io_out ? io_r_2_b : _GEN_3301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3303 = 8'h3 == r_count_15_io_out ? io_r_3_b : _GEN_3302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3304 = 8'h4 == r_count_15_io_out ? io_r_4_b : _GEN_3303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3305 = 8'h5 == r_count_15_io_out ? io_r_5_b : _GEN_3304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3306 = 8'h6 == r_count_15_io_out ? io_r_6_b : _GEN_3305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3307 = 8'h7 == r_count_15_io_out ? io_r_7_b : _GEN_3306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3308 = 8'h8 == r_count_15_io_out ? io_r_8_b : _GEN_3307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3309 = 8'h9 == r_count_15_io_out ? io_r_9_b : _GEN_3308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3310 = 8'ha == r_count_15_io_out ? io_r_10_b : _GEN_3309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3311 = 8'hb == r_count_15_io_out ? io_r_11_b : _GEN_3310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3312 = 8'hc == r_count_15_io_out ? io_r_12_b : _GEN_3311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3313 = 8'hd == r_count_15_io_out ? io_r_13_b : _GEN_3312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3314 = 8'he == r_count_15_io_out ? io_r_14_b : _GEN_3313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3315 = 8'hf == r_count_15_io_out ? io_r_15_b : _GEN_3314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3316 = 8'h10 == r_count_15_io_out ? io_r_16_b : _GEN_3315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3317 = 8'h11 == r_count_15_io_out ? io_r_17_b : _GEN_3316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3318 = 8'h12 == r_count_15_io_out ? io_r_18_b : _GEN_3317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3319 = 8'h13 == r_count_15_io_out ? io_r_19_b : _GEN_3318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3320 = 8'h14 == r_count_15_io_out ? io_r_20_b : _GEN_3319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3321 = 8'h15 == r_count_15_io_out ? io_r_21_b : _GEN_3320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3322 = 8'h16 == r_count_15_io_out ? io_r_22_b : _GEN_3321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3323 = 8'h17 == r_count_15_io_out ? io_r_23_b : _GEN_3322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3324 = 8'h18 == r_count_15_io_out ? io_r_24_b : _GEN_3323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3325 = 8'h19 == r_count_15_io_out ? io_r_25_b : _GEN_3324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3326 = 8'h1a == r_count_15_io_out ? io_r_26_b : _GEN_3325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3327 = 8'h1b == r_count_15_io_out ? io_r_27_b : _GEN_3326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3328 = 8'h1c == r_count_15_io_out ? io_r_28_b : _GEN_3327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3329 = 8'h1d == r_count_15_io_out ? io_r_29_b : _GEN_3328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3330 = 8'h1e == r_count_15_io_out ? io_r_30_b : _GEN_3329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3331 = 8'h1f == r_count_15_io_out ? io_r_31_b : _GEN_3330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3332 = 8'h20 == r_count_15_io_out ? io_r_32_b : _GEN_3331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3333 = 8'h21 == r_count_15_io_out ? io_r_33_b : _GEN_3332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3334 = 8'h22 == r_count_15_io_out ? io_r_34_b : _GEN_3333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3335 = 8'h23 == r_count_15_io_out ? io_r_35_b : _GEN_3334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3336 = 8'h24 == r_count_15_io_out ? io_r_36_b : _GEN_3335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3337 = 8'h25 == r_count_15_io_out ? io_r_37_b : _GEN_3336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3338 = 8'h26 == r_count_15_io_out ? io_r_38_b : _GEN_3337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3339 = 8'h27 == r_count_15_io_out ? io_r_39_b : _GEN_3338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3340 = 8'h28 == r_count_15_io_out ? io_r_40_b : _GEN_3339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3341 = 8'h29 == r_count_15_io_out ? io_r_41_b : _GEN_3340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3342 = 8'h2a == r_count_15_io_out ? io_r_42_b : _GEN_3341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3343 = 8'h2b == r_count_15_io_out ? io_r_43_b : _GEN_3342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3344 = 8'h2c == r_count_15_io_out ? io_r_44_b : _GEN_3343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3345 = 8'h2d == r_count_15_io_out ? io_r_45_b : _GEN_3344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3346 = 8'h2e == r_count_15_io_out ? io_r_46_b : _GEN_3345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3347 = 8'h2f == r_count_15_io_out ? io_r_47_b : _GEN_3346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3348 = 8'h30 == r_count_15_io_out ? io_r_48_b : _GEN_3347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3349 = 8'h31 == r_count_15_io_out ? io_r_49_b : _GEN_3348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3350 = 8'h32 == r_count_15_io_out ? io_r_50_b : _GEN_3349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3351 = 8'h33 == r_count_15_io_out ? io_r_51_b : _GEN_3350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3352 = 8'h34 == r_count_15_io_out ? io_r_52_b : _GEN_3351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3353 = 8'h35 == r_count_15_io_out ? io_r_53_b : _GEN_3352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3354 = 8'h36 == r_count_15_io_out ? io_r_54_b : _GEN_3353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3355 = 8'h37 == r_count_15_io_out ? io_r_55_b : _GEN_3354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3356 = 8'h38 == r_count_15_io_out ? io_r_56_b : _GEN_3355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3357 = 8'h39 == r_count_15_io_out ? io_r_57_b : _GEN_3356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3358 = 8'h3a == r_count_15_io_out ? io_r_58_b : _GEN_3357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3359 = 8'h3b == r_count_15_io_out ? io_r_59_b : _GEN_3358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3360 = 8'h3c == r_count_15_io_out ? io_r_60_b : _GEN_3359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3361 = 8'h3d == r_count_15_io_out ? io_r_61_b : _GEN_3360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3362 = 8'h3e == r_count_15_io_out ? io_r_62_b : _GEN_3361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3363 = 8'h3f == r_count_15_io_out ? io_r_63_b : _GEN_3362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3364 = 8'h40 == r_count_15_io_out ? io_r_64_b : _GEN_3363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3365 = 8'h41 == r_count_15_io_out ? io_r_65_b : _GEN_3364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3366 = 8'h42 == r_count_15_io_out ? io_r_66_b : _GEN_3365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3367 = 8'h43 == r_count_15_io_out ? io_r_67_b : _GEN_3366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3368 = 8'h44 == r_count_15_io_out ? io_r_68_b : _GEN_3367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3369 = 8'h45 == r_count_15_io_out ? io_r_69_b : _GEN_3368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3370 = 8'h46 == r_count_15_io_out ? io_r_70_b : _GEN_3369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3371 = 8'h47 == r_count_15_io_out ? io_r_71_b : _GEN_3370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3372 = 8'h48 == r_count_15_io_out ? io_r_72_b : _GEN_3371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3373 = 8'h49 == r_count_15_io_out ? io_r_73_b : _GEN_3372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3374 = 8'h4a == r_count_15_io_out ? io_r_74_b : _GEN_3373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3375 = 8'h4b == r_count_15_io_out ? io_r_75_b : _GEN_3374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3376 = 8'h4c == r_count_15_io_out ? io_r_76_b : _GEN_3375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3377 = 8'h4d == r_count_15_io_out ? io_r_77_b : _GEN_3376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3378 = 8'h4e == r_count_15_io_out ? io_r_78_b : _GEN_3377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3379 = 8'h4f == r_count_15_io_out ? io_r_79_b : _GEN_3378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3380 = 8'h50 == r_count_15_io_out ? io_r_80_b : _GEN_3379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3381 = 8'h51 == r_count_15_io_out ? io_r_81_b : _GEN_3380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3382 = 8'h52 == r_count_15_io_out ? io_r_82_b : _GEN_3381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3383 = 8'h53 == r_count_15_io_out ? io_r_83_b : _GEN_3382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3384 = 8'h54 == r_count_15_io_out ? io_r_84_b : _GEN_3383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3385 = 8'h55 == r_count_15_io_out ? io_r_85_b : _GEN_3384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3386 = 8'h56 == r_count_15_io_out ? io_r_86_b : _GEN_3385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3387 = 8'h57 == r_count_15_io_out ? io_r_87_b : _GEN_3386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3388 = 8'h58 == r_count_15_io_out ? io_r_88_b : _GEN_3387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3389 = 8'h59 == r_count_15_io_out ? io_r_89_b : _GEN_3388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3390 = 8'h5a == r_count_15_io_out ? io_r_90_b : _GEN_3389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3391 = 8'h5b == r_count_15_io_out ? io_r_91_b : _GEN_3390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3392 = 8'h5c == r_count_15_io_out ? io_r_92_b : _GEN_3391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3393 = 8'h5d == r_count_15_io_out ? io_r_93_b : _GEN_3392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3394 = 8'h5e == r_count_15_io_out ? io_r_94_b : _GEN_3393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3395 = 8'h5f == r_count_15_io_out ? io_r_95_b : _GEN_3394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3396 = 8'h60 == r_count_15_io_out ? io_r_96_b : _GEN_3395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3397 = 8'h61 == r_count_15_io_out ? io_r_97_b : _GEN_3396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3398 = 8'h62 == r_count_15_io_out ? io_r_98_b : _GEN_3397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3399 = 8'h63 == r_count_15_io_out ? io_r_99_b : _GEN_3398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3400 = 8'h64 == r_count_15_io_out ? io_r_100_b : _GEN_3399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3401 = 8'h65 == r_count_15_io_out ? io_r_101_b : _GEN_3400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3402 = 8'h66 == r_count_15_io_out ? io_r_102_b : _GEN_3401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3403 = 8'h67 == r_count_15_io_out ? io_r_103_b : _GEN_3402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3404 = 8'h68 == r_count_15_io_out ? io_r_104_b : _GEN_3403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3405 = 8'h69 == r_count_15_io_out ? io_r_105_b : _GEN_3404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3406 = 8'h6a == r_count_15_io_out ? io_r_106_b : _GEN_3405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3407 = 8'h6b == r_count_15_io_out ? io_r_107_b : _GEN_3406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3408 = 8'h6c == r_count_15_io_out ? io_r_108_b : _GEN_3407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3409 = 8'h6d == r_count_15_io_out ? io_r_109_b : _GEN_3408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3410 = 8'h6e == r_count_15_io_out ? io_r_110_b : _GEN_3409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3411 = 8'h6f == r_count_15_io_out ? io_r_111_b : _GEN_3410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3412 = 8'h70 == r_count_15_io_out ? io_r_112_b : _GEN_3411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3413 = 8'h71 == r_count_15_io_out ? io_r_113_b : _GEN_3412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3414 = 8'h72 == r_count_15_io_out ? io_r_114_b : _GEN_3413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3415 = 8'h73 == r_count_15_io_out ? io_r_115_b : _GEN_3414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3416 = 8'h74 == r_count_15_io_out ? io_r_116_b : _GEN_3415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3417 = 8'h75 == r_count_15_io_out ? io_r_117_b : _GEN_3416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3418 = 8'h76 == r_count_15_io_out ? io_r_118_b : _GEN_3417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3419 = 8'h77 == r_count_15_io_out ? io_r_119_b : _GEN_3418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3420 = 8'h78 == r_count_15_io_out ? io_r_120_b : _GEN_3419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3421 = 8'h79 == r_count_15_io_out ? io_r_121_b : _GEN_3420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3422 = 8'h7a == r_count_15_io_out ? io_r_122_b : _GEN_3421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3423 = 8'h7b == r_count_15_io_out ? io_r_123_b : _GEN_3422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3424 = 8'h7c == r_count_15_io_out ? io_r_124_b : _GEN_3423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3425 = 8'h7d == r_count_15_io_out ? io_r_125_b : _GEN_3424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3426 = 8'h7e == r_count_15_io_out ? io_r_126_b : _GEN_3425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3427 = 8'h7f == r_count_15_io_out ? io_r_127_b : _GEN_3426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3428 = 8'h80 == r_count_15_io_out ? io_r_128_b : _GEN_3427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3429 = 8'h81 == r_count_15_io_out ? io_r_129_b : _GEN_3428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3430 = 8'h82 == r_count_15_io_out ? io_r_130_b : _GEN_3429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3431 = 8'h83 == r_count_15_io_out ? io_r_131_b : _GEN_3430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3432 = 8'h84 == r_count_15_io_out ? io_r_132_b : _GEN_3431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3433 = 8'h85 == r_count_15_io_out ? io_r_133_b : _GEN_3432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3434 = 8'h86 == r_count_15_io_out ? io_r_134_b : _GEN_3433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3435 = 8'h87 == r_count_15_io_out ? io_r_135_b : _GEN_3434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3436 = 8'h88 == r_count_15_io_out ? io_r_136_b : _GEN_3435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3437 = 8'h89 == r_count_15_io_out ? io_r_137_b : _GEN_3436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3438 = 8'h8a == r_count_15_io_out ? io_r_138_b : _GEN_3437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3439 = 8'h8b == r_count_15_io_out ? io_r_139_b : _GEN_3438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3440 = 8'h8c == r_count_15_io_out ? io_r_140_b : _GEN_3439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3441 = 8'h8d == r_count_15_io_out ? io_r_141_b : _GEN_3440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3442 = 8'h8e == r_count_15_io_out ? io_r_142_b : _GEN_3441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3443 = 8'h8f == r_count_15_io_out ? io_r_143_b : _GEN_3442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3444 = 8'h90 == r_count_15_io_out ? io_r_144_b : _GEN_3443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3445 = 8'h91 == r_count_15_io_out ? io_r_145_b : _GEN_3444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3446 = 8'h92 == r_count_15_io_out ? io_r_146_b : _GEN_3445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3447 = 8'h93 == r_count_15_io_out ? io_r_147_b : _GEN_3446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3448 = 8'h94 == r_count_15_io_out ? io_r_148_b : _GEN_3447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3449 = 8'h95 == r_count_15_io_out ? io_r_149_b : _GEN_3448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3450 = 8'h96 == r_count_15_io_out ? io_r_150_b : _GEN_3449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3451 = 8'h97 == r_count_15_io_out ? io_r_151_b : _GEN_3450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3452 = 8'h98 == r_count_15_io_out ? io_r_152_b : _GEN_3451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3453 = 8'h99 == r_count_15_io_out ? io_r_153_b : _GEN_3452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3454 = 8'h9a == r_count_15_io_out ? io_r_154_b : _GEN_3453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3455 = 8'h9b == r_count_15_io_out ? io_r_155_b : _GEN_3454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3456 = 8'h9c == r_count_15_io_out ? io_r_156_b : _GEN_3455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3457 = 8'h9d == r_count_15_io_out ? io_r_157_b : _GEN_3456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3458 = 8'h9e == r_count_15_io_out ? io_r_158_b : _GEN_3457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3459 = 8'h9f == r_count_15_io_out ? io_r_159_b : _GEN_3458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3460 = 8'ha0 == r_count_15_io_out ? io_r_160_b : _GEN_3459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3461 = 8'ha1 == r_count_15_io_out ? io_r_161_b : _GEN_3460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3462 = 8'ha2 == r_count_15_io_out ? io_r_162_b : _GEN_3461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3463 = 8'ha3 == r_count_15_io_out ? io_r_163_b : _GEN_3462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3464 = 8'ha4 == r_count_15_io_out ? io_r_164_b : _GEN_3463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3465 = 8'ha5 == r_count_15_io_out ? io_r_165_b : _GEN_3464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3466 = 8'ha6 == r_count_15_io_out ? io_r_166_b : _GEN_3465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3467 = 8'ha7 == r_count_15_io_out ? io_r_167_b : _GEN_3466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3468 = 8'ha8 == r_count_15_io_out ? io_r_168_b : _GEN_3467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3469 = 8'ha9 == r_count_15_io_out ? io_r_169_b : _GEN_3468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3470 = 8'haa == r_count_15_io_out ? io_r_170_b : _GEN_3469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3471 = 8'hab == r_count_15_io_out ? io_r_171_b : _GEN_3470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3472 = 8'hac == r_count_15_io_out ? io_r_172_b : _GEN_3471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3473 = 8'had == r_count_15_io_out ? io_r_173_b : _GEN_3472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3474 = 8'hae == r_count_15_io_out ? io_r_174_b : _GEN_3473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3475 = 8'haf == r_count_15_io_out ? io_r_175_b : _GEN_3474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3476 = 8'hb0 == r_count_15_io_out ? io_r_176_b : _GEN_3475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3477 = 8'hb1 == r_count_15_io_out ? io_r_177_b : _GEN_3476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3478 = 8'hb2 == r_count_15_io_out ? io_r_178_b : _GEN_3477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3479 = 8'hb3 == r_count_15_io_out ? io_r_179_b : _GEN_3478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3480 = 8'hb4 == r_count_15_io_out ? io_r_180_b : _GEN_3479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3481 = 8'hb5 == r_count_15_io_out ? io_r_181_b : _GEN_3480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3482 = 8'hb6 == r_count_15_io_out ? io_r_182_b : _GEN_3481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3483 = 8'hb7 == r_count_15_io_out ? io_r_183_b : _GEN_3482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3484 = 8'hb8 == r_count_15_io_out ? io_r_184_b : _GEN_3483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3485 = 8'hb9 == r_count_15_io_out ? io_r_185_b : _GEN_3484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3486 = 8'hba == r_count_15_io_out ? io_r_186_b : _GEN_3485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3487 = 8'hbb == r_count_15_io_out ? io_r_187_b : _GEN_3486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3488 = 8'hbc == r_count_15_io_out ? io_r_188_b : _GEN_3487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3489 = 8'hbd == r_count_15_io_out ? io_r_189_b : _GEN_3488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3490 = 8'hbe == r_count_15_io_out ? io_r_190_b : _GEN_3489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3491 = 8'hbf == r_count_15_io_out ? io_r_191_b : _GEN_3490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3492 = 8'hc0 == r_count_15_io_out ? io_r_192_b : _GEN_3491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3493 = 8'hc1 == r_count_15_io_out ? io_r_193_b : _GEN_3492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3494 = 8'hc2 == r_count_15_io_out ? io_r_194_b : _GEN_3493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3495 = 8'hc3 == r_count_15_io_out ? io_r_195_b : _GEN_3494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3496 = 8'hc4 == r_count_15_io_out ? io_r_196_b : _GEN_3495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3497 = 8'hc5 == r_count_15_io_out ? io_r_197_b : _GEN_3496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3498 = 8'hc6 == r_count_15_io_out ? io_r_198_b : _GEN_3497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3501 = 8'h1 == r_count_16_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3502 = 8'h2 == r_count_16_io_out ? io_r_2_b : _GEN_3501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3503 = 8'h3 == r_count_16_io_out ? io_r_3_b : _GEN_3502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3504 = 8'h4 == r_count_16_io_out ? io_r_4_b : _GEN_3503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3505 = 8'h5 == r_count_16_io_out ? io_r_5_b : _GEN_3504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3506 = 8'h6 == r_count_16_io_out ? io_r_6_b : _GEN_3505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3507 = 8'h7 == r_count_16_io_out ? io_r_7_b : _GEN_3506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3508 = 8'h8 == r_count_16_io_out ? io_r_8_b : _GEN_3507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3509 = 8'h9 == r_count_16_io_out ? io_r_9_b : _GEN_3508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3510 = 8'ha == r_count_16_io_out ? io_r_10_b : _GEN_3509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3511 = 8'hb == r_count_16_io_out ? io_r_11_b : _GEN_3510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3512 = 8'hc == r_count_16_io_out ? io_r_12_b : _GEN_3511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3513 = 8'hd == r_count_16_io_out ? io_r_13_b : _GEN_3512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3514 = 8'he == r_count_16_io_out ? io_r_14_b : _GEN_3513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3515 = 8'hf == r_count_16_io_out ? io_r_15_b : _GEN_3514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3516 = 8'h10 == r_count_16_io_out ? io_r_16_b : _GEN_3515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3517 = 8'h11 == r_count_16_io_out ? io_r_17_b : _GEN_3516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3518 = 8'h12 == r_count_16_io_out ? io_r_18_b : _GEN_3517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3519 = 8'h13 == r_count_16_io_out ? io_r_19_b : _GEN_3518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3520 = 8'h14 == r_count_16_io_out ? io_r_20_b : _GEN_3519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3521 = 8'h15 == r_count_16_io_out ? io_r_21_b : _GEN_3520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3522 = 8'h16 == r_count_16_io_out ? io_r_22_b : _GEN_3521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3523 = 8'h17 == r_count_16_io_out ? io_r_23_b : _GEN_3522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3524 = 8'h18 == r_count_16_io_out ? io_r_24_b : _GEN_3523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3525 = 8'h19 == r_count_16_io_out ? io_r_25_b : _GEN_3524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3526 = 8'h1a == r_count_16_io_out ? io_r_26_b : _GEN_3525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3527 = 8'h1b == r_count_16_io_out ? io_r_27_b : _GEN_3526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3528 = 8'h1c == r_count_16_io_out ? io_r_28_b : _GEN_3527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3529 = 8'h1d == r_count_16_io_out ? io_r_29_b : _GEN_3528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3530 = 8'h1e == r_count_16_io_out ? io_r_30_b : _GEN_3529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3531 = 8'h1f == r_count_16_io_out ? io_r_31_b : _GEN_3530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3532 = 8'h20 == r_count_16_io_out ? io_r_32_b : _GEN_3531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3533 = 8'h21 == r_count_16_io_out ? io_r_33_b : _GEN_3532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3534 = 8'h22 == r_count_16_io_out ? io_r_34_b : _GEN_3533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3535 = 8'h23 == r_count_16_io_out ? io_r_35_b : _GEN_3534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3536 = 8'h24 == r_count_16_io_out ? io_r_36_b : _GEN_3535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3537 = 8'h25 == r_count_16_io_out ? io_r_37_b : _GEN_3536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3538 = 8'h26 == r_count_16_io_out ? io_r_38_b : _GEN_3537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3539 = 8'h27 == r_count_16_io_out ? io_r_39_b : _GEN_3538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3540 = 8'h28 == r_count_16_io_out ? io_r_40_b : _GEN_3539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3541 = 8'h29 == r_count_16_io_out ? io_r_41_b : _GEN_3540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3542 = 8'h2a == r_count_16_io_out ? io_r_42_b : _GEN_3541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3543 = 8'h2b == r_count_16_io_out ? io_r_43_b : _GEN_3542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3544 = 8'h2c == r_count_16_io_out ? io_r_44_b : _GEN_3543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3545 = 8'h2d == r_count_16_io_out ? io_r_45_b : _GEN_3544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3546 = 8'h2e == r_count_16_io_out ? io_r_46_b : _GEN_3545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3547 = 8'h2f == r_count_16_io_out ? io_r_47_b : _GEN_3546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3548 = 8'h30 == r_count_16_io_out ? io_r_48_b : _GEN_3547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3549 = 8'h31 == r_count_16_io_out ? io_r_49_b : _GEN_3548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3550 = 8'h32 == r_count_16_io_out ? io_r_50_b : _GEN_3549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3551 = 8'h33 == r_count_16_io_out ? io_r_51_b : _GEN_3550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3552 = 8'h34 == r_count_16_io_out ? io_r_52_b : _GEN_3551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3553 = 8'h35 == r_count_16_io_out ? io_r_53_b : _GEN_3552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3554 = 8'h36 == r_count_16_io_out ? io_r_54_b : _GEN_3553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3555 = 8'h37 == r_count_16_io_out ? io_r_55_b : _GEN_3554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3556 = 8'h38 == r_count_16_io_out ? io_r_56_b : _GEN_3555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3557 = 8'h39 == r_count_16_io_out ? io_r_57_b : _GEN_3556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3558 = 8'h3a == r_count_16_io_out ? io_r_58_b : _GEN_3557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3559 = 8'h3b == r_count_16_io_out ? io_r_59_b : _GEN_3558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3560 = 8'h3c == r_count_16_io_out ? io_r_60_b : _GEN_3559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3561 = 8'h3d == r_count_16_io_out ? io_r_61_b : _GEN_3560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3562 = 8'h3e == r_count_16_io_out ? io_r_62_b : _GEN_3561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3563 = 8'h3f == r_count_16_io_out ? io_r_63_b : _GEN_3562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3564 = 8'h40 == r_count_16_io_out ? io_r_64_b : _GEN_3563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3565 = 8'h41 == r_count_16_io_out ? io_r_65_b : _GEN_3564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3566 = 8'h42 == r_count_16_io_out ? io_r_66_b : _GEN_3565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3567 = 8'h43 == r_count_16_io_out ? io_r_67_b : _GEN_3566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3568 = 8'h44 == r_count_16_io_out ? io_r_68_b : _GEN_3567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3569 = 8'h45 == r_count_16_io_out ? io_r_69_b : _GEN_3568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3570 = 8'h46 == r_count_16_io_out ? io_r_70_b : _GEN_3569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3571 = 8'h47 == r_count_16_io_out ? io_r_71_b : _GEN_3570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3572 = 8'h48 == r_count_16_io_out ? io_r_72_b : _GEN_3571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3573 = 8'h49 == r_count_16_io_out ? io_r_73_b : _GEN_3572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3574 = 8'h4a == r_count_16_io_out ? io_r_74_b : _GEN_3573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3575 = 8'h4b == r_count_16_io_out ? io_r_75_b : _GEN_3574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3576 = 8'h4c == r_count_16_io_out ? io_r_76_b : _GEN_3575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3577 = 8'h4d == r_count_16_io_out ? io_r_77_b : _GEN_3576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3578 = 8'h4e == r_count_16_io_out ? io_r_78_b : _GEN_3577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3579 = 8'h4f == r_count_16_io_out ? io_r_79_b : _GEN_3578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3580 = 8'h50 == r_count_16_io_out ? io_r_80_b : _GEN_3579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3581 = 8'h51 == r_count_16_io_out ? io_r_81_b : _GEN_3580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3582 = 8'h52 == r_count_16_io_out ? io_r_82_b : _GEN_3581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3583 = 8'h53 == r_count_16_io_out ? io_r_83_b : _GEN_3582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3584 = 8'h54 == r_count_16_io_out ? io_r_84_b : _GEN_3583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3585 = 8'h55 == r_count_16_io_out ? io_r_85_b : _GEN_3584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3586 = 8'h56 == r_count_16_io_out ? io_r_86_b : _GEN_3585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3587 = 8'h57 == r_count_16_io_out ? io_r_87_b : _GEN_3586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3588 = 8'h58 == r_count_16_io_out ? io_r_88_b : _GEN_3587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3589 = 8'h59 == r_count_16_io_out ? io_r_89_b : _GEN_3588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3590 = 8'h5a == r_count_16_io_out ? io_r_90_b : _GEN_3589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3591 = 8'h5b == r_count_16_io_out ? io_r_91_b : _GEN_3590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3592 = 8'h5c == r_count_16_io_out ? io_r_92_b : _GEN_3591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3593 = 8'h5d == r_count_16_io_out ? io_r_93_b : _GEN_3592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3594 = 8'h5e == r_count_16_io_out ? io_r_94_b : _GEN_3593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3595 = 8'h5f == r_count_16_io_out ? io_r_95_b : _GEN_3594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3596 = 8'h60 == r_count_16_io_out ? io_r_96_b : _GEN_3595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3597 = 8'h61 == r_count_16_io_out ? io_r_97_b : _GEN_3596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3598 = 8'h62 == r_count_16_io_out ? io_r_98_b : _GEN_3597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3599 = 8'h63 == r_count_16_io_out ? io_r_99_b : _GEN_3598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3600 = 8'h64 == r_count_16_io_out ? io_r_100_b : _GEN_3599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3601 = 8'h65 == r_count_16_io_out ? io_r_101_b : _GEN_3600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3602 = 8'h66 == r_count_16_io_out ? io_r_102_b : _GEN_3601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3603 = 8'h67 == r_count_16_io_out ? io_r_103_b : _GEN_3602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3604 = 8'h68 == r_count_16_io_out ? io_r_104_b : _GEN_3603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3605 = 8'h69 == r_count_16_io_out ? io_r_105_b : _GEN_3604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3606 = 8'h6a == r_count_16_io_out ? io_r_106_b : _GEN_3605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3607 = 8'h6b == r_count_16_io_out ? io_r_107_b : _GEN_3606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3608 = 8'h6c == r_count_16_io_out ? io_r_108_b : _GEN_3607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3609 = 8'h6d == r_count_16_io_out ? io_r_109_b : _GEN_3608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3610 = 8'h6e == r_count_16_io_out ? io_r_110_b : _GEN_3609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3611 = 8'h6f == r_count_16_io_out ? io_r_111_b : _GEN_3610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3612 = 8'h70 == r_count_16_io_out ? io_r_112_b : _GEN_3611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3613 = 8'h71 == r_count_16_io_out ? io_r_113_b : _GEN_3612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3614 = 8'h72 == r_count_16_io_out ? io_r_114_b : _GEN_3613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3615 = 8'h73 == r_count_16_io_out ? io_r_115_b : _GEN_3614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3616 = 8'h74 == r_count_16_io_out ? io_r_116_b : _GEN_3615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3617 = 8'h75 == r_count_16_io_out ? io_r_117_b : _GEN_3616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3618 = 8'h76 == r_count_16_io_out ? io_r_118_b : _GEN_3617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3619 = 8'h77 == r_count_16_io_out ? io_r_119_b : _GEN_3618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3620 = 8'h78 == r_count_16_io_out ? io_r_120_b : _GEN_3619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3621 = 8'h79 == r_count_16_io_out ? io_r_121_b : _GEN_3620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3622 = 8'h7a == r_count_16_io_out ? io_r_122_b : _GEN_3621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3623 = 8'h7b == r_count_16_io_out ? io_r_123_b : _GEN_3622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3624 = 8'h7c == r_count_16_io_out ? io_r_124_b : _GEN_3623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3625 = 8'h7d == r_count_16_io_out ? io_r_125_b : _GEN_3624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3626 = 8'h7e == r_count_16_io_out ? io_r_126_b : _GEN_3625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3627 = 8'h7f == r_count_16_io_out ? io_r_127_b : _GEN_3626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3628 = 8'h80 == r_count_16_io_out ? io_r_128_b : _GEN_3627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3629 = 8'h81 == r_count_16_io_out ? io_r_129_b : _GEN_3628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3630 = 8'h82 == r_count_16_io_out ? io_r_130_b : _GEN_3629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3631 = 8'h83 == r_count_16_io_out ? io_r_131_b : _GEN_3630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3632 = 8'h84 == r_count_16_io_out ? io_r_132_b : _GEN_3631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3633 = 8'h85 == r_count_16_io_out ? io_r_133_b : _GEN_3632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3634 = 8'h86 == r_count_16_io_out ? io_r_134_b : _GEN_3633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3635 = 8'h87 == r_count_16_io_out ? io_r_135_b : _GEN_3634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3636 = 8'h88 == r_count_16_io_out ? io_r_136_b : _GEN_3635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3637 = 8'h89 == r_count_16_io_out ? io_r_137_b : _GEN_3636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3638 = 8'h8a == r_count_16_io_out ? io_r_138_b : _GEN_3637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3639 = 8'h8b == r_count_16_io_out ? io_r_139_b : _GEN_3638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3640 = 8'h8c == r_count_16_io_out ? io_r_140_b : _GEN_3639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3641 = 8'h8d == r_count_16_io_out ? io_r_141_b : _GEN_3640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3642 = 8'h8e == r_count_16_io_out ? io_r_142_b : _GEN_3641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3643 = 8'h8f == r_count_16_io_out ? io_r_143_b : _GEN_3642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3644 = 8'h90 == r_count_16_io_out ? io_r_144_b : _GEN_3643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3645 = 8'h91 == r_count_16_io_out ? io_r_145_b : _GEN_3644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3646 = 8'h92 == r_count_16_io_out ? io_r_146_b : _GEN_3645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3647 = 8'h93 == r_count_16_io_out ? io_r_147_b : _GEN_3646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3648 = 8'h94 == r_count_16_io_out ? io_r_148_b : _GEN_3647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3649 = 8'h95 == r_count_16_io_out ? io_r_149_b : _GEN_3648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3650 = 8'h96 == r_count_16_io_out ? io_r_150_b : _GEN_3649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3651 = 8'h97 == r_count_16_io_out ? io_r_151_b : _GEN_3650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3652 = 8'h98 == r_count_16_io_out ? io_r_152_b : _GEN_3651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3653 = 8'h99 == r_count_16_io_out ? io_r_153_b : _GEN_3652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3654 = 8'h9a == r_count_16_io_out ? io_r_154_b : _GEN_3653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3655 = 8'h9b == r_count_16_io_out ? io_r_155_b : _GEN_3654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3656 = 8'h9c == r_count_16_io_out ? io_r_156_b : _GEN_3655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3657 = 8'h9d == r_count_16_io_out ? io_r_157_b : _GEN_3656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3658 = 8'h9e == r_count_16_io_out ? io_r_158_b : _GEN_3657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3659 = 8'h9f == r_count_16_io_out ? io_r_159_b : _GEN_3658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3660 = 8'ha0 == r_count_16_io_out ? io_r_160_b : _GEN_3659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3661 = 8'ha1 == r_count_16_io_out ? io_r_161_b : _GEN_3660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3662 = 8'ha2 == r_count_16_io_out ? io_r_162_b : _GEN_3661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3663 = 8'ha3 == r_count_16_io_out ? io_r_163_b : _GEN_3662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3664 = 8'ha4 == r_count_16_io_out ? io_r_164_b : _GEN_3663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3665 = 8'ha5 == r_count_16_io_out ? io_r_165_b : _GEN_3664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3666 = 8'ha6 == r_count_16_io_out ? io_r_166_b : _GEN_3665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3667 = 8'ha7 == r_count_16_io_out ? io_r_167_b : _GEN_3666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3668 = 8'ha8 == r_count_16_io_out ? io_r_168_b : _GEN_3667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3669 = 8'ha9 == r_count_16_io_out ? io_r_169_b : _GEN_3668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3670 = 8'haa == r_count_16_io_out ? io_r_170_b : _GEN_3669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3671 = 8'hab == r_count_16_io_out ? io_r_171_b : _GEN_3670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3672 = 8'hac == r_count_16_io_out ? io_r_172_b : _GEN_3671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3673 = 8'had == r_count_16_io_out ? io_r_173_b : _GEN_3672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3674 = 8'hae == r_count_16_io_out ? io_r_174_b : _GEN_3673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3675 = 8'haf == r_count_16_io_out ? io_r_175_b : _GEN_3674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3676 = 8'hb0 == r_count_16_io_out ? io_r_176_b : _GEN_3675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3677 = 8'hb1 == r_count_16_io_out ? io_r_177_b : _GEN_3676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3678 = 8'hb2 == r_count_16_io_out ? io_r_178_b : _GEN_3677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3679 = 8'hb3 == r_count_16_io_out ? io_r_179_b : _GEN_3678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3680 = 8'hb4 == r_count_16_io_out ? io_r_180_b : _GEN_3679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3681 = 8'hb5 == r_count_16_io_out ? io_r_181_b : _GEN_3680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3682 = 8'hb6 == r_count_16_io_out ? io_r_182_b : _GEN_3681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3683 = 8'hb7 == r_count_16_io_out ? io_r_183_b : _GEN_3682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3684 = 8'hb8 == r_count_16_io_out ? io_r_184_b : _GEN_3683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3685 = 8'hb9 == r_count_16_io_out ? io_r_185_b : _GEN_3684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3686 = 8'hba == r_count_16_io_out ? io_r_186_b : _GEN_3685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3687 = 8'hbb == r_count_16_io_out ? io_r_187_b : _GEN_3686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3688 = 8'hbc == r_count_16_io_out ? io_r_188_b : _GEN_3687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3689 = 8'hbd == r_count_16_io_out ? io_r_189_b : _GEN_3688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3690 = 8'hbe == r_count_16_io_out ? io_r_190_b : _GEN_3689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3691 = 8'hbf == r_count_16_io_out ? io_r_191_b : _GEN_3690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3692 = 8'hc0 == r_count_16_io_out ? io_r_192_b : _GEN_3691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3693 = 8'hc1 == r_count_16_io_out ? io_r_193_b : _GEN_3692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3694 = 8'hc2 == r_count_16_io_out ? io_r_194_b : _GEN_3693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3695 = 8'hc3 == r_count_16_io_out ? io_r_195_b : _GEN_3694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3696 = 8'hc4 == r_count_16_io_out ? io_r_196_b : _GEN_3695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3697 = 8'hc5 == r_count_16_io_out ? io_r_197_b : _GEN_3696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3698 = 8'hc6 == r_count_16_io_out ? io_r_198_b : _GEN_3697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3701 = 8'h1 == r_count_17_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3702 = 8'h2 == r_count_17_io_out ? io_r_2_b : _GEN_3701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3703 = 8'h3 == r_count_17_io_out ? io_r_3_b : _GEN_3702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3704 = 8'h4 == r_count_17_io_out ? io_r_4_b : _GEN_3703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3705 = 8'h5 == r_count_17_io_out ? io_r_5_b : _GEN_3704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3706 = 8'h6 == r_count_17_io_out ? io_r_6_b : _GEN_3705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3707 = 8'h7 == r_count_17_io_out ? io_r_7_b : _GEN_3706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3708 = 8'h8 == r_count_17_io_out ? io_r_8_b : _GEN_3707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3709 = 8'h9 == r_count_17_io_out ? io_r_9_b : _GEN_3708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3710 = 8'ha == r_count_17_io_out ? io_r_10_b : _GEN_3709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3711 = 8'hb == r_count_17_io_out ? io_r_11_b : _GEN_3710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3712 = 8'hc == r_count_17_io_out ? io_r_12_b : _GEN_3711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3713 = 8'hd == r_count_17_io_out ? io_r_13_b : _GEN_3712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3714 = 8'he == r_count_17_io_out ? io_r_14_b : _GEN_3713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3715 = 8'hf == r_count_17_io_out ? io_r_15_b : _GEN_3714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3716 = 8'h10 == r_count_17_io_out ? io_r_16_b : _GEN_3715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3717 = 8'h11 == r_count_17_io_out ? io_r_17_b : _GEN_3716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3718 = 8'h12 == r_count_17_io_out ? io_r_18_b : _GEN_3717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3719 = 8'h13 == r_count_17_io_out ? io_r_19_b : _GEN_3718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3720 = 8'h14 == r_count_17_io_out ? io_r_20_b : _GEN_3719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3721 = 8'h15 == r_count_17_io_out ? io_r_21_b : _GEN_3720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3722 = 8'h16 == r_count_17_io_out ? io_r_22_b : _GEN_3721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3723 = 8'h17 == r_count_17_io_out ? io_r_23_b : _GEN_3722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3724 = 8'h18 == r_count_17_io_out ? io_r_24_b : _GEN_3723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3725 = 8'h19 == r_count_17_io_out ? io_r_25_b : _GEN_3724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3726 = 8'h1a == r_count_17_io_out ? io_r_26_b : _GEN_3725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3727 = 8'h1b == r_count_17_io_out ? io_r_27_b : _GEN_3726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3728 = 8'h1c == r_count_17_io_out ? io_r_28_b : _GEN_3727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3729 = 8'h1d == r_count_17_io_out ? io_r_29_b : _GEN_3728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3730 = 8'h1e == r_count_17_io_out ? io_r_30_b : _GEN_3729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3731 = 8'h1f == r_count_17_io_out ? io_r_31_b : _GEN_3730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3732 = 8'h20 == r_count_17_io_out ? io_r_32_b : _GEN_3731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3733 = 8'h21 == r_count_17_io_out ? io_r_33_b : _GEN_3732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3734 = 8'h22 == r_count_17_io_out ? io_r_34_b : _GEN_3733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3735 = 8'h23 == r_count_17_io_out ? io_r_35_b : _GEN_3734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3736 = 8'h24 == r_count_17_io_out ? io_r_36_b : _GEN_3735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3737 = 8'h25 == r_count_17_io_out ? io_r_37_b : _GEN_3736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3738 = 8'h26 == r_count_17_io_out ? io_r_38_b : _GEN_3737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3739 = 8'h27 == r_count_17_io_out ? io_r_39_b : _GEN_3738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3740 = 8'h28 == r_count_17_io_out ? io_r_40_b : _GEN_3739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3741 = 8'h29 == r_count_17_io_out ? io_r_41_b : _GEN_3740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3742 = 8'h2a == r_count_17_io_out ? io_r_42_b : _GEN_3741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3743 = 8'h2b == r_count_17_io_out ? io_r_43_b : _GEN_3742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3744 = 8'h2c == r_count_17_io_out ? io_r_44_b : _GEN_3743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3745 = 8'h2d == r_count_17_io_out ? io_r_45_b : _GEN_3744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3746 = 8'h2e == r_count_17_io_out ? io_r_46_b : _GEN_3745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3747 = 8'h2f == r_count_17_io_out ? io_r_47_b : _GEN_3746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3748 = 8'h30 == r_count_17_io_out ? io_r_48_b : _GEN_3747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3749 = 8'h31 == r_count_17_io_out ? io_r_49_b : _GEN_3748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3750 = 8'h32 == r_count_17_io_out ? io_r_50_b : _GEN_3749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3751 = 8'h33 == r_count_17_io_out ? io_r_51_b : _GEN_3750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3752 = 8'h34 == r_count_17_io_out ? io_r_52_b : _GEN_3751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3753 = 8'h35 == r_count_17_io_out ? io_r_53_b : _GEN_3752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3754 = 8'h36 == r_count_17_io_out ? io_r_54_b : _GEN_3753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3755 = 8'h37 == r_count_17_io_out ? io_r_55_b : _GEN_3754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3756 = 8'h38 == r_count_17_io_out ? io_r_56_b : _GEN_3755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3757 = 8'h39 == r_count_17_io_out ? io_r_57_b : _GEN_3756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3758 = 8'h3a == r_count_17_io_out ? io_r_58_b : _GEN_3757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3759 = 8'h3b == r_count_17_io_out ? io_r_59_b : _GEN_3758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3760 = 8'h3c == r_count_17_io_out ? io_r_60_b : _GEN_3759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3761 = 8'h3d == r_count_17_io_out ? io_r_61_b : _GEN_3760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3762 = 8'h3e == r_count_17_io_out ? io_r_62_b : _GEN_3761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3763 = 8'h3f == r_count_17_io_out ? io_r_63_b : _GEN_3762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3764 = 8'h40 == r_count_17_io_out ? io_r_64_b : _GEN_3763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3765 = 8'h41 == r_count_17_io_out ? io_r_65_b : _GEN_3764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3766 = 8'h42 == r_count_17_io_out ? io_r_66_b : _GEN_3765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3767 = 8'h43 == r_count_17_io_out ? io_r_67_b : _GEN_3766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3768 = 8'h44 == r_count_17_io_out ? io_r_68_b : _GEN_3767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3769 = 8'h45 == r_count_17_io_out ? io_r_69_b : _GEN_3768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3770 = 8'h46 == r_count_17_io_out ? io_r_70_b : _GEN_3769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3771 = 8'h47 == r_count_17_io_out ? io_r_71_b : _GEN_3770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3772 = 8'h48 == r_count_17_io_out ? io_r_72_b : _GEN_3771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3773 = 8'h49 == r_count_17_io_out ? io_r_73_b : _GEN_3772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3774 = 8'h4a == r_count_17_io_out ? io_r_74_b : _GEN_3773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3775 = 8'h4b == r_count_17_io_out ? io_r_75_b : _GEN_3774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3776 = 8'h4c == r_count_17_io_out ? io_r_76_b : _GEN_3775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3777 = 8'h4d == r_count_17_io_out ? io_r_77_b : _GEN_3776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3778 = 8'h4e == r_count_17_io_out ? io_r_78_b : _GEN_3777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3779 = 8'h4f == r_count_17_io_out ? io_r_79_b : _GEN_3778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3780 = 8'h50 == r_count_17_io_out ? io_r_80_b : _GEN_3779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3781 = 8'h51 == r_count_17_io_out ? io_r_81_b : _GEN_3780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3782 = 8'h52 == r_count_17_io_out ? io_r_82_b : _GEN_3781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3783 = 8'h53 == r_count_17_io_out ? io_r_83_b : _GEN_3782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3784 = 8'h54 == r_count_17_io_out ? io_r_84_b : _GEN_3783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3785 = 8'h55 == r_count_17_io_out ? io_r_85_b : _GEN_3784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3786 = 8'h56 == r_count_17_io_out ? io_r_86_b : _GEN_3785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3787 = 8'h57 == r_count_17_io_out ? io_r_87_b : _GEN_3786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3788 = 8'h58 == r_count_17_io_out ? io_r_88_b : _GEN_3787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3789 = 8'h59 == r_count_17_io_out ? io_r_89_b : _GEN_3788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3790 = 8'h5a == r_count_17_io_out ? io_r_90_b : _GEN_3789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3791 = 8'h5b == r_count_17_io_out ? io_r_91_b : _GEN_3790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3792 = 8'h5c == r_count_17_io_out ? io_r_92_b : _GEN_3791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3793 = 8'h5d == r_count_17_io_out ? io_r_93_b : _GEN_3792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3794 = 8'h5e == r_count_17_io_out ? io_r_94_b : _GEN_3793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3795 = 8'h5f == r_count_17_io_out ? io_r_95_b : _GEN_3794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3796 = 8'h60 == r_count_17_io_out ? io_r_96_b : _GEN_3795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3797 = 8'h61 == r_count_17_io_out ? io_r_97_b : _GEN_3796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3798 = 8'h62 == r_count_17_io_out ? io_r_98_b : _GEN_3797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3799 = 8'h63 == r_count_17_io_out ? io_r_99_b : _GEN_3798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3800 = 8'h64 == r_count_17_io_out ? io_r_100_b : _GEN_3799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3801 = 8'h65 == r_count_17_io_out ? io_r_101_b : _GEN_3800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3802 = 8'h66 == r_count_17_io_out ? io_r_102_b : _GEN_3801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3803 = 8'h67 == r_count_17_io_out ? io_r_103_b : _GEN_3802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3804 = 8'h68 == r_count_17_io_out ? io_r_104_b : _GEN_3803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3805 = 8'h69 == r_count_17_io_out ? io_r_105_b : _GEN_3804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3806 = 8'h6a == r_count_17_io_out ? io_r_106_b : _GEN_3805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3807 = 8'h6b == r_count_17_io_out ? io_r_107_b : _GEN_3806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3808 = 8'h6c == r_count_17_io_out ? io_r_108_b : _GEN_3807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3809 = 8'h6d == r_count_17_io_out ? io_r_109_b : _GEN_3808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3810 = 8'h6e == r_count_17_io_out ? io_r_110_b : _GEN_3809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3811 = 8'h6f == r_count_17_io_out ? io_r_111_b : _GEN_3810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3812 = 8'h70 == r_count_17_io_out ? io_r_112_b : _GEN_3811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3813 = 8'h71 == r_count_17_io_out ? io_r_113_b : _GEN_3812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3814 = 8'h72 == r_count_17_io_out ? io_r_114_b : _GEN_3813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3815 = 8'h73 == r_count_17_io_out ? io_r_115_b : _GEN_3814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3816 = 8'h74 == r_count_17_io_out ? io_r_116_b : _GEN_3815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3817 = 8'h75 == r_count_17_io_out ? io_r_117_b : _GEN_3816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3818 = 8'h76 == r_count_17_io_out ? io_r_118_b : _GEN_3817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3819 = 8'h77 == r_count_17_io_out ? io_r_119_b : _GEN_3818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3820 = 8'h78 == r_count_17_io_out ? io_r_120_b : _GEN_3819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3821 = 8'h79 == r_count_17_io_out ? io_r_121_b : _GEN_3820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3822 = 8'h7a == r_count_17_io_out ? io_r_122_b : _GEN_3821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3823 = 8'h7b == r_count_17_io_out ? io_r_123_b : _GEN_3822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3824 = 8'h7c == r_count_17_io_out ? io_r_124_b : _GEN_3823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3825 = 8'h7d == r_count_17_io_out ? io_r_125_b : _GEN_3824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3826 = 8'h7e == r_count_17_io_out ? io_r_126_b : _GEN_3825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3827 = 8'h7f == r_count_17_io_out ? io_r_127_b : _GEN_3826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3828 = 8'h80 == r_count_17_io_out ? io_r_128_b : _GEN_3827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3829 = 8'h81 == r_count_17_io_out ? io_r_129_b : _GEN_3828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3830 = 8'h82 == r_count_17_io_out ? io_r_130_b : _GEN_3829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3831 = 8'h83 == r_count_17_io_out ? io_r_131_b : _GEN_3830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3832 = 8'h84 == r_count_17_io_out ? io_r_132_b : _GEN_3831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3833 = 8'h85 == r_count_17_io_out ? io_r_133_b : _GEN_3832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3834 = 8'h86 == r_count_17_io_out ? io_r_134_b : _GEN_3833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3835 = 8'h87 == r_count_17_io_out ? io_r_135_b : _GEN_3834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3836 = 8'h88 == r_count_17_io_out ? io_r_136_b : _GEN_3835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3837 = 8'h89 == r_count_17_io_out ? io_r_137_b : _GEN_3836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3838 = 8'h8a == r_count_17_io_out ? io_r_138_b : _GEN_3837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3839 = 8'h8b == r_count_17_io_out ? io_r_139_b : _GEN_3838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3840 = 8'h8c == r_count_17_io_out ? io_r_140_b : _GEN_3839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3841 = 8'h8d == r_count_17_io_out ? io_r_141_b : _GEN_3840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3842 = 8'h8e == r_count_17_io_out ? io_r_142_b : _GEN_3841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3843 = 8'h8f == r_count_17_io_out ? io_r_143_b : _GEN_3842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3844 = 8'h90 == r_count_17_io_out ? io_r_144_b : _GEN_3843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3845 = 8'h91 == r_count_17_io_out ? io_r_145_b : _GEN_3844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3846 = 8'h92 == r_count_17_io_out ? io_r_146_b : _GEN_3845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3847 = 8'h93 == r_count_17_io_out ? io_r_147_b : _GEN_3846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3848 = 8'h94 == r_count_17_io_out ? io_r_148_b : _GEN_3847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3849 = 8'h95 == r_count_17_io_out ? io_r_149_b : _GEN_3848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3850 = 8'h96 == r_count_17_io_out ? io_r_150_b : _GEN_3849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3851 = 8'h97 == r_count_17_io_out ? io_r_151_b : _GEN_3850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3852 = 8'h98 == r_count_17_io_out ? io_r_152_b : _GEN_3851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3853 = 8'h99 == r_count_17_io_out ? io_r_153_b : _GEN_3852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3854 = 8'h9a == r_count_17_io_out ? io_r_154_b : _GEN_3853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3855 = 8'h9b == r_count_17_io_out ? io_r_155_b : _GEN_3854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3856 = 8'h9c == r_count_17_io_out ? io_r_156_b : _GEN_3855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3857 = 8'h9d == r_count_17_io_out ? io_r_157_b : _GEN_3856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3858 = 8'h9e == r_count_17_io_out ? io_r_158_b : _GEN_3857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3859 = 8'h9f == r_count_17_io_out ? io_r_159_b : _GEN_3858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3860 = 8'ha0 == r_count_17_io_out ? io_r_160_b : _GEN_3859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3861 = 8'ha1 == r_count_17_io_out ? io_r_161_b : _GEN_3860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3862 = 8'ha2 == r_count_17_io_out ? io_r_162_b : _GEN_3861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3863 = 8'ha3 == r_count_17_io_out ? io_r_163_b : _GEN_3862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3864 = 8'ha4 == r_count_17_io_out ? io_r_164_b : _GEN_3863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3865 = 8'ha5 == r_count_17_io_out ? io_r_165_b : _GEN_3864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3866 = 8'ha6 == r_count_17_io_out ? io_r_166_b : _GEN_3865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3867 = 8'ha7 == r_count_17_io_out ? io_r_167_b : _GEN_3866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3868 = 8'ha8 == r_count_17_io_out ? io_r_168_b : _GEN_3867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3869 = 8'ha9 == r_count_17_io_out ? io_r_169_b : _GEN_3868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3870 = 8'haa == r_count_17_io_out ? io_r_170_b : _GEN_3869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3871 = 8'hab == r_count_17_io_out ? io_r_171_b : _GEN_3870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3872 = 8'hac == r_count_17_io_out ? io_r_172_b : _GEN_3871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3873 = 8'had == r_count_17_io_out ? io_r_173_b : _GEN_3872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3874 = 8'hae == r_count_17_io_out ? io_r_174_b : _GEN_3873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3875 = 8'haf == r_count_17_io_out ? io_r_175_b : _GEN_3874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3876 = 8'hb0 == r_count_17_io_out ? io_r_176_b : _GEN_3875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3877 = 8'hb1 == r_count_17_io_out ? io_r_177_b : _GEN_3876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3878 = 8'hb2 == r_count_17_io_out ? io_r_178_b : _GEN_3877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3879 = 8'hb3 == r_count_17_io_out ? io_r_179_b : _GEN_3878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3880 = 8'hb4 == r_count_17_io_out ? io_r_180_b : _GEN_3879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3881 = 8'hb5 == r_count_17_io_out ? io_r_181_b : _GEN_3880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3882 = 8'hb6 == r_count_17_io_out ? io_r_182_b : _GEN_3881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3883 = 8'hb7 == r_count_17_io_out ? io_r_183_b : _GEN_3882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3884 = 8'hb8 == r_count_17_io_out ? io_r_184_b : _GEN_3883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3885 = 8'hb9 == r_count_17_io_out ? io_r_185_b : _GEN_3884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3886 = 8'hba == r_count_17_io_out ? io_r_186_b : _GEN_3885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3887 = 8'hbb == r_count_17_io_out ? io_r_187_b : _GEN_3886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3888 = 8'hbc == r_count_17_io_out ? io_r_188_b : _GEN_3887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3889 = 8'hbd == r_count_17_io_out ? io_r_189_b : _GEN_3888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3890 = 8'hbe == r_count_17_io_out ? io_r_190_b : _GEN_3889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3891 = 8'hbf == r_count_17_io_out ? io_r_191_b : _GEN_3890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3892 = 8'hc0 == r_count_17_io_out ? io_r_192_b : _GEN_3891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3893 = 8'hc1 == r_count_17_io_out ? io_r_193_b : _GEN_3892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3894 = 8'hc2 == r_count_17_io_out ? io_r_194_b : _GEN_3893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3895 = 8'hc3 == r_count_17_io_out ? io_r_195_b : _GEN_3894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3896 = 8'hc4 == r_count_17_io_out ? io_r_196_b : _GEN_3895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3897 = 8'hc5 == r_count_17_io_out ? io_r_197_b : _GEN_3896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3898 = 8'hc6 == r_count_17_io_out ? io_r_198_b : _GEN_3897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3901 = 8'h1 == r_count_18_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3902 = 8'h2 == r_count_18_io_out ? io_r_2_b : _GEN_3901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3903 = 8'h3 == r_count_18_io_out ? io_r_3_b : _GEN_3902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3904 = 8'h4 == r_count_18_io_out ? io_r_4_b : _GEN_3903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3905 = 8'h5 == r_count_18_io_out ? io_r_5_b : _GEN_3904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3906 = 8'h6 == r_count_18_io_out ? io_r_6_b : _GEN_3905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3907 = 8'h7 == r_count_18_io_out ? io_r_7_b : _GEN_3906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3908 = 8'h8 == r_count_18_io_out ? io_r_8_b : _GEN_3907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3909 = 8'h9 == r_count_18_io_out ? io_r_9_b : _GEN_3908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3910 = 8'ha == r_count_18_io_out ? io_r_10_b : _GEN_3909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3911 = 8'hb == r_count_18_io_out ? io_r_11_b : _GEN_3910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3912 = 8'hc == r_count_18_io_out ? io_r_12_b : _GEN_3911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3913 = 8'hd == r_count_18_io_out ? io_r_13_b : _GEN_3912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3914 = 8'he == r_count_18_io_out ? io_r_14_b : _GEN_3913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3915 = 8'hf == r_count_18_io_out ? io_r_15_b : _GEN_3914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3916 = 8'h10 == r_count_18_io_out ? io_r_16_b : _GEN_3915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3917 = 8'h11 == r_count_18_io_out ? io_r_17_b : _GEN_3916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3918 = 8'h12 == r_count_18_io_out ? io_r_18_b : _GEN_3917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3919 = 8'h13 == r_count_18_io_out ? io_r_19_b : _GEN_3918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3920 = 8'h14 == r_count_18_io_out ? io_r_20_b : _GEN_3919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3921 = 8'h15 == r_count_18_io_out ? io_r_21_b : _GEN_3920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3922 = 8'h16 == r_count_18_io_out ? io_r_22_b : _GEN_3921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3923 = 8'h17 == r_count_18_io_out ? io_r_23_b : _GEN_3922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3924 = 8'h18 == r_count_18_io_out ? io_r_24_b : _GEN_3923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3925 = 8'h19 == r_count_18_io_out ? io_r_25_b : _GEN_3924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3926 = 8'h1a == r_count_18_io_out ? io_r_26_b : _GEN_3925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3927 = 8'h1b == r_count_18_io_out ? io_r_27_b : _GEN_3926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3928 = 8'h1c == r_count_18_io_out ? io_r_28_b : _GEN_3927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3929 = 8'h1d == r_count_18_io_out ? io_r_29_b : _GEN_3928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3930 = 8'h1e == r_count_18_io_out ? io_r_30_b : _GEN_3929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3931 = 8'h1f == r_count_18_io_out ? io_r_31_b : _GEN_3930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3932 = 8'h20 == r_count_18_io_out ? io_r_32_b : _GEN_3931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3933 = 8'h21 == r_count_18_io_out ? io_r_33_b : _GEN_3932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3934 = 8'h22 == r_count_18_io_out ? io_r_34_b : _GEN_3933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3935 = 8'h23 == r_count_18_io_out ? io_r_35_b : _GEN_3934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3936 = 8'h24 == r_count_18_io_out ? io_r_36_b : _GEN_3935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3937 = 8'h25 == r_count_18_io_out ? io_r_37_b : _GEN_3936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3938 = 8'h26 == r_count_18_io_out ? io_r_38_b : _GEN_3937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3939 = 8'h27 == r_count_18_io_out ? io_r_39_b : _GEN_3938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3940 = 8'h28 == r_count_18_io_out ? io_r_40_b : _GEN_3939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3941 = 8'h29 == r_count_18_io_out ? io_r_41_b : _GEN_3940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3942 = 8'h2a == r_count_18_io_out ? io_r_42_b : _GEN_3941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3943 = 8'h2b == r_count_18_io_out ? io_r_43_b : _GEN_3942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3944 = 8'h2c == r_count_18_io_out ? io_r_44_b : _GEN_3943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3945 = 8'h2d == r_count_18_io_out ? io_r_45_b : _GEN_3944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3946 = 8'h2e == r_count_18_io_out ? io_r_46_b : _GEN_3945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3947 = 8'h2f == r_count_18_io_out ? io_r_47_b : _GEN_3946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3948 = 8'h30 == r_count_18_io_out ? io_r_48_b : _GEN_3947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3949 = 8'h31 == r_count_18_io_out ? io_r_49_b : _GEN_3948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3950 = 8'h32 == r_count_18_io_out ? io_r_50_b : _GEN_3949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3951 = 8'h33 == r_count_18_io_out ? io_r_51_b : _GEN_3950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3952 = 8'h34 == r_count_18_io_out ? io_r_52_b : _GEN_3951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3953 = 8'h35 == r_count_18_io_out ? io_r_53_b : _GEN_3952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3954 = 8'h36 == r_count_18_io_out ? io_r_54_b : _GEN_3953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3955 = 8'h37 == r_count_18_io_out ? io_r_55_b : _GEN_3954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3956 = 8'h38 == r_count_18_io_out ? io_r_56_b : _GEN_3955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3957 = 8'h39 == r_count_18_io_out ? io_r_57_b : _GEN_3956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3958 = 8'h3a == r_count_18_io_out ? io_r_58_b : _GEN_3957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3959 = 8'h3b == r_count_18_io_out ? io_r_59_b : _GEN_3958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3960 = 8'h3c == r_count_18_io_out ? io_r_60_b : _GEN_3959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3961 = 8'h3d == r_count_18_io_out ? io_r_61_b : _GEN_3960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3962 = 8'h3e == r_count_18_io_out ? io_r_62_b : _GEN_3961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3963 = 8'h3f == r_count_18_io_out ? io_r_63_b : _GEN_3962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3964 = 8'h40 == r_count_18_io_out ? io_r_64_b : _GEN_3963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3965 = 8'h41 == r_count_18_io_out ? io_r_65_b : _GEN_3964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3966 = 8'h42 == r_count_18_io_out ? io_r_66_b : _GEN_3965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3967 = 8'h43 == r_count_18_io_out ? io_r_67_b : _GEN_3966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3968 = 8'h44 == r_count_18_io_out ? io_r_68_b : _GEN_3967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3969 = 8'h45 == r_count_18_io_out ? io_r_69_b : _GEN_3968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3970 = 8'h46 == r_count_18_io_out ? io_r_70_b : _GEN_3969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3971 = 8'h47 == r_count_18_io_out ? io_r_71_b : _GEN_3970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3972 = 8'h48 == r_count_18_io_out ? io_r_72_b : _GEN_3971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3973 = 8'h49 == r_count_18_io_out ? io_r_73_b : _GEN_3972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3974 = 8'h4a == r_count_18_io_out ? io_r_74_b : _GEN_3973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3975 = 8'h4b == r_count_18_io_out ? io_r_75_b : _GEN_3974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3976 = 8'h4c == r_count_18_io_out ? io_r_76_b : _GEN_3975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3977 = 8'h4d == r_count_18_io_out ? io_r_77_b : _GEN_3976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3978 = 8'h4e == r_count_18_io_out ? io_r_78_b : _GEN_3977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3979 = 8'h4f == r_count_18_io_out ? io_r_79_b : _GEN_3978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3980 = 8'h50 == r_count_18_io_out ? io_r_80_b : _GEN_3979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3981 = 8'h51 == r_count_18_io_out ? io_r_81_b : _GEN_3980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3982 = 8'h52 == r_count_18_io_out ? io_r_82_b : _GEN_3981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3983 = 8'h53 == r_count_18_io_out ? io_r_83_b : _GEN_3982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3984 = 8'h54 == r_count_18_io_out ? io_r_84_b : _GEN_3983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3985 = 8'h55 == r_count_18_io_out ? io_r_85_b : _GEN_3984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3986 = 8'h56 == r_count_18_io_out ? io_r_86_b : _GEN_3985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3987 = 8'h57 == r_count_18_io_out ? io_r_87_b : _GEN_3986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3988 = 8'h58 == r_count_18_io_out ? io_r_88_b : _GEN_3987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3989 = 8'h59 == r_count_18_io_out ? io_r_89_b : _GEN_3988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3990 = 8'h5a == r_count_18_io_out ? io_r_90_b : _GEN_3989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3991 = 8'h5b == r_count_18_io_out ? io_r_91_b : _GEN_3990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3992 = 8'h5c == r_count_18_io_out ? io_r_92_b : _GEN_3991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3993 = 8'h5d == r_count_18_io_out ? io_r_93_b : _GEN_3992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3994 = 8'h5e == r_count_18_io_out ? io_r_94_b : _GEN_3993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3995 = 8'h5f == r_count_18_io_out ? io_r_95_b : _GEN_3994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3996 = 8'h60 == r_count_18_io_out ? io_r_96_b : _GEN_3995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3997 = 8'h61 == r_count_18_io_out ? io_r_97_b : _GEN_3996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3998 = 8'h62 == r_count_18_io_out ? io_r_98_b : _GEN_3997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3999 = 8'h63 == r_count_18_io_out ? io_r_99_b : _GEN_3998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4000 = 8'h64 == r_count_18_io_out ? io_r_100_b : _GEN_3999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4001 = 8'h65 == r_count_18_io_out ? io_r_101_b : _GEN_4000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4002 = 8'h66 == r_count_18_io_out ? io_r_102_b : _GEN_4001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4003 = 8'h67 == r_count_18_io_out ? io_r_103_b : _GEN_4002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4004 = 8'h68 == r_count_18_io_out ? io_r_104_b : _GEN_4003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4005 = 8'h69 == r_count_18_io_out ? io_r_105_b : _GEN_4004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4006 = 8'h6a == r_count_18_io_out ? io_r_106_b : _GEN_4005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4007 = 8'h6b == r_count_18_io_out ? io_r_107_b : _GEN_4006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4008 = 8'h6c == r_count_18_io_out ? io_r_108_b : _GEN_4007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4009 = 8'h6d == r_count_18_io_out ? io_r_109_b : _GEN_4008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4010 = 8'h6e == r_count_18_io_out ? io_r_110_b : _GEN_4009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4011 = 8'h6f == r_count_18_io_out ? io_r_111_b : _GEN_4010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4012 = 8'h70 == r_count_18_io_out ? io_r_112_b : _GEN_4011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4013 = 8'h71 == r_count_18_io_out ? io_r_113_b : _GEN_4012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4014 = 8'h72 == r_count_18_io_out ? io_r_114_b : _GEN_4013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4015 = 8'h73 == r_count_18_io_out ? io_r_115_b : _GEN_4014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4016 = 8'h74 == r_count_18_io_out ? io_r_116_b : _GEN_4015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4017 = 8'h75 == r_count_18_io_out ? io_r_117_b : _GEN_4016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4018 = 8'h76 == r_count_18_io_out ? io_r_118_b : _GEN_4017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4019 = 8'h77 == r_count_18_io_out ? io_r_119_b : _GEN_4018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4020 = 8'h78 == r_count_18_io_out ? io_r_120_b : _GEN_4019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4021 = 8'h79 == r_count_18_io_out ? io_r_121_b : _GEN_4020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4022 = 8'h7a == r_count_18_io_out ? io_r_122_b : _GEN_4021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4023 = 8'h7b == r_count_18_io_out ? io_r_123_b : _GEN_4022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4024 = 8'h7c == r_count_18_io_out ? io_r_124_b : _GEN_4023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4025 = 8'h7d == r_count_18_io_out ? io_r_125_b : _GEN_4024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4026 = 8'h7e == r_count_18_io_out ? io_r_126_b : _GEN_4025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4027 = 8'h7f == r_count_18_io_out ? io_r_127_b : _GEN_4026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4028 = 8'h80 == r_count_18_io_out ? io_r_128_b : _GEN_4027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4029 = 8'h81 == r_count_18_io_out ? io_r_129_b : _GEN_4028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4030 = 8'h82 == r_count_18_io_out ? io_r_130_b : _GEN_4029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4031 = 8'h83 == r_count_18_io_out ? io_r_131_b : _GEN_4030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4032 = 8'h84 == r_count_18_io_out ? io_r_132_b : _GEN_4031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4033 = 8'h85 == r_count_18_io_out ? io_r_133_b : _GEN_4032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4034 = 8'h86 == r_count_18_io_out ? io_r_134_b : _GEN_4033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4035 = 8'h87 == r_count_18_io_out ? io_r_135_b : _GEN_4034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4036 = 8'h88 == r_count_18_io_out ? io_r_136_b : _GEN_4035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4037 = 8'h89 == r_count_18_io_out ? io_r_137_b : _GEN_4036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4038 = 8'h8a == r_count_18_io_out ? io_r_138_b : _GEN_4037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4039 = 8'h8b == r_count_18_io_out ? io_r_139_b : _GEN_4038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4040 = 8'h8c == r_count_18_io_out ? io_r_140_b : _GEN_4039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4041 = 8'h8d == r_count_18_io_out ? io_r_141_b : _GEN_4040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4042 = 8'h8e == r_count_18_io_out ? io_r_142_b : _GEN_4041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4043 = 8'h8f == r_count_18_io_out ? io_r_143_b : _GEN_4042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4044 = 8'h90 == r_count_18_io_out ? io_r_144_b : _GEN_4043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4045 = 8'h91 == r_count_18_io_out ? io_r_145_b : _GEN_4044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4046 = 8'h92 == r_count_18_io_out ? io_r_146_b : _GEN_4045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4047 = 8'h93 == r_count_18_io_out ? io_r_147_b : _GEN_4046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4048 = 8'h94 == r_count_18_io_out ? io_r_148_b : _GEN_4047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4049 = 8'h95 == r_count_18_io_out ? io_r_149_b : _GEN_4048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4050 = 8'h96 == r_count_18_io_out ? io_r_150_b : _GEN_4049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4051 = 8'h97 == r_count_18_io_out ? io_r_151_b : _GEN_4050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4052 = 8'h98 == r_count_18_io_out ? io_r_152_b : _GEN_4051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4053 = 8'h99 == r_count_18_io_out ? io_r_153_b : _GEN_4052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4054 = 8'h9a == r_count_18_io_out ? io_r_154_b : _GEN_4053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4055 = 8'h9b == r_count_18_io_out ? io_r_155_b : _GEN_4054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4056 = 8'h9c == r_count_18_io_out ? io_r_156_b : _GEN_4055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4057 = 8'h9d == r_count_18_io_out ? io_r_157_b : _GEN_4056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4058 = 8'h9e == r_count_18_io_out ? io_r_158_b : _GEN_4057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4059 = 8'h9f == r_count_18_io_out ? io_r_159_b : _GEN_4058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4060 = 8'ha0 == r_count_18_io_out ? io_r_160_b : _GEN_4059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4061 = 8'ha1 == r_count_18_io_out ? io_r_161_b : _GEN_4060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4062 = 8'ha2 == r_count_18_io_out ? io_r_162_b : _GEN_4061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4063 = 8'ha3 == r_count_18_io_out ? io_r_163_b : _GEN_4062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4064 = 8'ha4 == r_count_18_io_out ? io_r_164_b : _GEN_4063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4065 = 8'ha5 == r_count_18_io_out ? io_r_165_b : _GEN_4064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4066 = 8'ha6 == r_count_18_io_out ? io_r_166_b : _GEN_4065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4067 = 8'ha7 == r_count_18_io_out ? io_r_167_b : _GEN_4066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4068 = 8'ha8 == r_count_18_io_out ? io_r_168_b : _GEN_4067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4069 = 8'ha9 == r_count_18_io_out ? io_r_169_b : _GEN_4068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4070 = 8'haa == r_count_18_io_out ? io_r_170_b : _GEN_4069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4071 = 8'hab == r_count_18_io_out ? io_r_171_b : _GEN_4070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4072 = 8'hac == r_count_18_io_out ? io_r_172_b : _GEN_4071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4073 = 8'had == r_count_18_io_out ? io_r_173_b : _GEN_4072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4074 = 8'hae == r_count_18_io_out ? io_r_174_b : _GEN_4073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4075 = 8'haf == r_count_18_io_out ? io_r_175_b : _GEN_4074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4076 = 8'hb0 == r_count_18_io_out ? io_r_176_b : _GEN_4075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4077 = 8'hb1 == r_count_18_io_out ? io_r_177_b : _GEN_4076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4078 = 8'hb2 == r_count_18_io_out ? io_r_178_b : _GEN_4077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4079 = 8'hb3 == r_count_18_io_out ? io_r_179_b : _GEN_4078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4080 = 8'hb4 == r_count_18_io_out ? io_r_180_b : _GEN_4079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4081 = 8'hb5 == r_count_18_io_out ? io_r_181_b : _GEN_4080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4082 = 8'hb6 == r_count_18_io_out ? io_r_182_b : _GEN_4081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4083 = 8'hb7 == r_count_18_io_out ? io_r_183_b : _GEN_4082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4084 = 8'hb8 == r_count_18_io_out ? io_r_184_b : _GEN_4083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4085 = 8'hb9 == r_count_18_io_out ? io_r_185_b : _GEN_4084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4086 = 8'hba == r_count_18_io_out ? io_r_186_b : _GEN_4085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4087 = 8'hbb == r_count_18_io_out ? io_r_187_b : _GEN_4086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4088 = 8'hbc == r_count_18_io_out ? io_r_188_b : _GEN_4087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4089 = 8'hbd == r_count_18_io_out ? io_r_189_b : _GEN_4088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4090 = 8'hbe == r_count_18_io_out ? io_r_190_b : _GEN_4089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4091 = 8'hbf == r_count_18_io_out ? io_r_191_b : _GEN_4090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4092 = 8'hc0 == r_count_18_io_out ? io_r_192_b : _GEN_4091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4093 = 8'hc1 == r_count_18_io_out ? io_r_193_b : _GEN_4092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4094 = 8'hc2 == r_count_18_io_out ? io_r_194_b : _GEN_4093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4095 = 8'hc3 == r_count_18_io_out ? io_r_195_b : _GEN_4094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4096 = 8'hc4 == r_count_18_io_out ? io_r_196_b : _GEN_4095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4097 = 8'hc5 == r_count_18_io_out ? io_r_197_b : _GEN_4096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4098 = 8'hc6 == r_count_18_io_out ? io_r_198_b : _GEN_4097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4101 = 8'h1 == r_count_19_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4102 = 8'h2 == r_count_19_io_out ? io_r_2_b : _GEN_4101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4103 = 8'h3 == r_count_19_io_out ? io_r_3_b : _GEN_4102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4104 = 8'h4 == r_count_19_io_out ? io_r_4_b : _GEN_4103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4105 = 8'h5 == r_count_19_io_out ? io_r_5_b : _GEN_4104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4106 = 8'h6 == r_count_19_io_out ? io_r_6_b : _GEN_4105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4107 = 8'h7 == r_count_19_io_out ? io_r_7_b : _GEN_4106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4108 = 8'h8 == r_count_19_io_out ? io_r_8_b : _GEN_4107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4109 = 8'h9 == r_count_19_io_out ? io_r_9_b : _GEN_4108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4110 = 8'ha == r_count_19_io_out ? io_r_10_b : _GEN_4109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4111 = 8'hb == r_count_19_io_out ? io_r_11_b : _GEN_4110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4112 = 8'hc == r_count_19_io_out ? io_r_12_b : _GEN_4111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4113 = 8'hd == r_count_19_io_out ? io_r_13_b : _GEN_4112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4114 = 8'he == r_count_19_io_out ? io_r_14_b : _GEN_4113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4115 = 8'hf == r_count_19_io_out ? io_r_15_b : _GEN_4114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4116 = 8'h10 == r_count_19_io_out ? io_r_16_b : _GEN_4115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4117 = 8'h11 == r_count_19_io_out ? io_r_17_b : _GEN_4116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4118 = 8'h12 == r_count_19_io_out ? io_r_18_b : _GEN_4117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4119 = 8'h13 == r_count_19_io_out ? io_r_19_b : _GEN_4118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4120 = 8'h14 == r_count_19_io_out ? io_r_20_b : _GEN_4119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4121 = 8'h15 == r_count_19_io_out ? io_r_21_b : _GEN_4120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4122 = 8'h16 == r_count_19_io_out ? io_r_22_b : _GEN_4121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4123 = 8'h17 == r_count_19_io_out ? io_r_23_b : _GEN_4122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4124 = 8'h18 == r_count_19_io_out ? io_r_24_b : _GEN_4123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4125 = 8'h19 == r_count_19_io_out ? io_r_25_b : _GEN_4124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4126 = 8'h1a == r_count_19_io_out ? io_r_26_b : _GEN_4125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4127 = 8'h1b == r_count_19_io_out ? io_r_27_b : _GEN_4126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4128 = 8'h1c == r_count_19_io_out ? io_r_28_b : _GEN_4127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4129 = 8'h1d == r_count_19_io_out ? io_r_29_b : _GEN_4128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4130 = 8'h1e == r_count_19_io_out ? io_r_30_b : _GEN_4129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4131 = 8'h1f == r_count_19_io_out ? io_r_31_b : _GEN_4130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4132 = 8'h20 == r_count_19_io_out ? io_r_32_b : _GEN_4131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4133 = 8'h21 == r_count_19_io_out ? io_r_33_b : _GEN_4132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4134 = 8'h22 == r_count_19_io_out ? io_r_34_b : _GEN_4133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4135 = 8'h23 == r_count_19_io_out ? io_r_35_b : _GEN_4134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4136 = 8'h24 == r_count_19_io_out ? io_r_36_b : _GEN_4135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4137 = 8'h25 == r_count_19_io_out ? io_r_37_b : _GEN_4136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4138 = 8'h26 == r_count_19_io_out ? io_r_38_b : _GEN_4137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4139 = 8'h27 == r_count_19_io_out ? io_r_39_b : _GEN_4138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4140 = 8'h28 == r_count_19_io_out ? io_r_40_b : _GEN_4139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4141 = 8'h29 == r_count_19_io_out ? io_r_41_b : _GEN_4140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4142 = 8'h2a == r_count_19_io_out ? io_r_42_b : _GEN_4141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4143 = 8'h2b == r_count_19_io_out ? io_r_43_b : _GEN_4142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4144 = 8'h2c == r_count_19_io_out ? io_r_44_b : _GEN_4143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4145 = 8'h2d == r_count_19_io_out ? io_r_45_b : _GEN_4144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4146 = 8'h2e == r_count_19_io_out ? io_r_46_b : _GEN_4145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4147 = 8'h2f == r_count_19_io_out ? io_r_47_b : _GEN_4146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4148 = 8'h30 == r_count_19_io_out ? io_r_48_b : _GEN_4147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4149 = 8'h31 == r_count_19_io_out ? io_r_49_b : _GEN_4148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4150 = 8'h32 == r_count_19_io_out ? io_r_50_b : _GEN_4149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4151 = 8'h33 == r_count_19_io_out ? io_r_51_b : _GEN_4150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4152 = 8'h34 == r_count_19_io_out ? io_r_52_b : _GEN_4151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4153 = 8'h35 == r_count_19_io_out ? io_r_53_b : _GEN_4152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4154 = 8'h36 == r_count_19_io_out ? io_r_54_b : _GEN_4153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4155 = 8'h37 == r_count_19_io_out ? io_r_55_b : _GEN_4154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4156 = 8'h38 == r_count_19_io_out ? io_r_56_b : _GEN_4155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4157 = 8'h39 == r_count_19_io_out ? io_r_57_b : _GEN_4156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4158 = 8'h3a == r_count_19_io_out ? io_r_58_b : _GEN_4157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4159 = 8'h3b == r_count_19_io_out ? io_r_59_b : _GEN_4158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4160 = 8'h3c == r_count_19_io_out ? io_r_60_b : _GEN_4159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4161 = 8'h3d == r_count_19_io_out ? io_r_61_b : _GEN_4160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4162 = 8'h3e == r_count_19_io_out ? io_r_62_b : _GEN_4161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4163 = 8'h3f == r_count_19_io_out ? io_r_63_b : _GEN_4162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4164 = 8'h40 == r_count_19_io_out ? io_r_64_b : _GEN_4163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4165 = 8'h41 == r_count_19_io_out ? io_r_65_b : _GEN_4164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4166 = 8'h42 == r_count_19_io_out ? io_r_66_b : _GEN_4165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4167 = 8'h43 == r_count_19_io_out ? io_r_67_b : _GEN_4166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4168 = 8'h44 == r_count_19_io_out ? io_r_68_b : _GEN_4167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4169 = 8'h45 == r_count_19_io_out ? io_r_69_b : _GEN_4168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4170 = 8'h46 == r_count_19_io_out ? io_r_70_b : _GEN_4169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4171 = 8'h47 == r_count_19_io_out ? io_r_71_b : _GEN_4170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4172 = 8'h48 == r_count_19_io_out ? io_r_72_b : _GEN_4171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4173 = 8'h49 == r_count_19_io_out ? io_r_73_b : _GEN_4172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4174 = 8'h4a == r_count_19_io_out ? io_r_74_b : _GEN_4173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4175 = 8'h4b == r_count_19_io_out ? io_r_75_b : _GEN_4174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4176 = 8'h4c == r_count_19_io_out ? io_r_76_b : _GEN_4175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4177 = 8'h4d == r_count_19_io_out ? io_r_77_b : _GEN_4176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4178 = 8'h4e == r_count_19_io_out ? io_r_78_b : _GEN_4177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4179 = 8'h4f == r_count_19_io_out ? io_r_79_b : _GEN_4178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4180 = 8'h50 == r_count_19_io_out ? io_r_80_b : _GEN_4179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4181 = 8'h51 == r_count_19_io_out ? io_r_81_b : _GEN_4180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4182 = 8'h52 == r_count_19_io_out ? io_r_82_b : _GEN_4181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4183 = 8'h53 == r_count_19_io_out ? io_r_83_b : _GEN_4182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4184 = 8'h54 == r_count_19_io_out ? io_r_84_b : _GEN_4183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4185 = 8'h55 == r_count_19_io_out ? io_r_85_b : _GEN_4184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4186 = 8'h56 == r_count_19_io_out ? io_r_86_b : _GEN_4185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4187 = 8'h57 == r_count_19_io_out ? io_r_87_b : _GEN_4186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4188 = 8'h58 == r_count_19_io_out ? io_r_88_b : _GEN_4187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4189 = 8'h59 == r_count_19_io_out ? io_r_89_b : _GEN_4188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4190 = 8'h5a == r_count_19_io_out ? io_r_90_b : _GEN_4189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4191 = 8'h5b == r_count_19_io_out ? io_r_91_b : _GEN_4190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4192 = 8'h5c == r_count_19_io_out ? io_r_92_b : _GEN_4191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4193 = 8'h5d == r_count_19_io_out ? io_r_93_b : _GEN_4192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4194 = 8'h5e == r_count_19_io_out ? io_r_94_b : _GEN_4193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4195 = 8'h5f == r_count_19_io_out ? io_r_95_b : _GEN_4194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4196 = 8'h60 == r_count_19_io_out ? io_r_96_b : _GEN_4195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4197 = 8'h61 == r_count_19_io_out ? io_r_97_b : _GEN_4196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4198 = 8'h62 == r_count_19_io_out ? io_r_98_b : _GEN_4197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4199 = 8'h63 == r_count_19_io_out ? io_r_99_b : _GEN_4198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4200 = 8'h64 == r_count_19_io_out ? io_r_100_b : _GEN_4199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4201 = 8'h65 == r_count_19_io_out ? io_r_101_b : _GEN_4200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4202 = 8'h66 == r_count_19_io_out ? io_r_102_b : _GEN_4201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4203 = 8'h67 == r_count_19_io_out ? io_r_103_b : _GEN_4202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4204 = 8'h68 == r_count_19_io_out ? io_r_104_b : _GEN_4203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4205 = 8'h69 == r_count_19_io_out ? io_r_105_b : _GEN_4204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4206 = 8'h6a == r_count_19_io_out ? io_r_106_b : _GEN_4205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4207 = 8'h6b == r_count_19_io_out ? io_r_107_b : _GEN_4206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4208 = 8'h6c == r_count_19_io_out ? io_r_108_b : _GEN_4207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4209 = 8'h6d == r_count_19_io_out ? io_r_109_b : _GEN_4208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4210 = 8'h6e == r_count_19_io_out ? io_r_110_b : _GEN_4209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4211 = 8'h6f == r_count_19_io_out ? io_r_111_b : _GEN_4210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4212 = 8'h70 == r_count_19_io_out ? io_r_112_b : _GEN_4211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4213 = 8'h71 == r_count_19_io_out ? io_r_113_b : _GEN_4212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4214 = 8'h72 == r_count_19_io_out ? io_r_114_b : _GEN_4213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4215 = 8'h73 == r_count_19_io_out ? io_r_115_b : _GEN_4214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4216 = 8'h74 == r_count_19_io_out ? io_r_116_b : _GEN_4215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4217 = 8'h75 == r_count_19_io_out ? io_r_117_b : _GEN_4216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4218 = 8'h76 == r_count_19_io_out ? io_r_118_b : _GEN_4217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4219 = 8'h77 == r_count_19_io_out ? io_r_119_b : _GEN_4218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4220 = 8'h78 == r_count_19_io_out ? io_r_120_b : _GEN_4219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4221 = 8'h79 == r_count_19_io_out ? io_r_121_b : _GEN_4220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4222 = 8'h7a == r_count_19_io_out ? io_r_122_b : _GEN_4221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4223 = 8'h7b == r_count_19_io_out ? io_r_123_b : _GEN_4222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4224 = 8'h7c == r_count_19_io_out ? io_r_124_b : _GEN_4223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4225 = 8'h7d == r_count_19_io_out ? io_r_125_b : _GEN_4224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4226 = 8'h7e == r_count_19_io_out ? io_r_126_b : _GEN_4225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4227 = 8'h7f == r_count_19_io_out ? io_r_127_b : _GEN_4226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4228 = 8'h80 == r_count_19_io_out ? io_r_128_b : _GEN_4227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4229 = 8'h81 == r_count_19_io_out ? io_r_129_b : _GEN_4228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4230 = 8'h82 == r_count_19_io_out ? io_r_130_b : _GEN_4229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4231 = 8'h83 == r_count_19_io_out ? io_r_131_b : _GEN_4230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4232 = 8'h84 == r_count_19_io_out ? io_r_132_b : _GEN_4231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4233 = 8'h85 == r_count_19_io_out ? io_r_133_b : _GEN_4232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4234 = 8'h86 == r_count_19_io_out ? io_r_134_b : _GEN_4233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4235 = 8'h87 == r_count_19_io_out ? io_r_135_b : _GEN_4234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4236 = 8'h88 == r_count_19_io_out ? io_r_136_b : _GEN_4235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4237 = 8'h89 == r_count_19_io_out ? io_r_137_b : _GEN_4236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4238 = 8'h8a == r_count_19_io_out ? io_r_138_b : _GEN_4237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4239 = 8'h8b == r_count_19_io_out ? io_r_139_b : _GEN_4238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4240 = 8'h8c == r_count_19_io_out ? io_r_140_b : _GEN_4239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4241 = 8'h8d == r_count_19_io_out ? io_r_141_b : _GEN_4240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4242 = 8'h8e == r_count_19_io_out ? io_r_142_b : _GEN_4241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4243 = 8'h8f == r_count_19_io_out ? io_r_143_b : _GEN_4242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4244 = 8'h90 == r_count_19_io_out ? io_r_144_b : _GEN_4243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4245 = 8'h91 == r_count_19_io_out ? io_r_145_b : _GEN_4244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4246 = 8'h92 == r_count_19_io_out ? io_r_146_b : _GEN_4245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4247 = 8'h93 == r_count_19_io_out ? io_r_147_b : _GEN_4246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4248 = 8'h94 == r_count_19_io_out ? io_r_148_b : _GEN_4247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4249 = 8'h95 == r_count_19_io_out ? io_r_149_b : _GEN_4248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4250 = 8'h96 == r_count_19_io_out ? io_r_150_b : _GEN_4249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4251 = 8'h97 == r_count_19_io_out ? io_r_151_b : _GEN_4250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4252 = 8'h98 == r_count_19_io_out ? io_r_152_b : _GEN_4251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4253 = 8'h99 == r_count_19_io_out ? io_r_153_b : _GEN_4252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4254 = 8'h9a == r_count_19_io_out ? io_r_154_b : _GEN_4253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4255 = 8'h9b == r_count_19_io_out ? io_r_155_b : _GEN_4254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4256 = 8'h9c == r_count_19_io_out ? io_r_156_b : _GEN_4255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4257 = 8'h9d == r_count_19_io_out ? io_r_157_b : _GEN_4256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4258 = 8'h9e == r_count_19_io_out ? io_r_158_b : _GEN_4257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4259 = 8'h9f == r_count_19_io_out ? io_r_159_b : _GEN_4258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4260 = 8'ha0 == r_count_19_io_out ? io_r_160_b : _GEN_4259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4261 = 8'ha1 == r_count_19_io_out ? io_r_161_b : _GEN_4260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4262 = 8'ha2 == r_count_19_io_out ? io_r_162_b : _GEN_4261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4263 = 8'ha3 == r_count_19_io_out ? io_r_163_b : _GEN_4262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4264 = 8'ha4 == r_count_19_io_out ? io_r_164_b : _GEN_4263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4265 = 8'ha5 == r_count_19_io_out ? io_r_165_b : _GEN_4264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4266 = 8'ha6 == r_count_19_io_out ? io_r_166_b : _GEN_4265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4267 = 8'ha7 == r_count_19_io_out ? io_r_167_b : _GEN_4266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4268 = 8'ha8 == r_count_19_io_out ? io_r_168_b : _GEN_4267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4269 = 8'ha9 == r_count_19_io_out ? io_r_169_b : _GEN_4268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4270 = 8'haa == r_count_19_io_out ? io_r_170_b : _GEN_4269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4271 = 8'hab == r_count_19_io_out ? io_r_171_b : _GEN_4270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4272 = 8'hac == r_count_19_io_out ? io_r_172_b : _GEN_4271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4273 = 8'had == r_count_19_io_out ? io_r_173_b : _GEN_4272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4274 = 8'hae == r_count_19_io_out ? io_r_174_b : _GEN_4273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4275 = 8'haf == r_count_19_io_out ? io_r_175_b : _GEN_4274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4276 = 8'hb0 == r_count_19_io_out ? io_r_176_b : _GEN_4275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4277 = 8'hb1 == r_count_19_io_out ? io_r_177_b : _GEN_4276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4278 = 8'hb2 == r_count_19_io_out ? io_r_178_b : _GEN_4277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4279 = 8'hb3 == r_count_19_io_out ? io_r_179_b : _GEN_4278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4280 = 8'hb4 == r_count_19_io_out ? io_r_180_b : _GEN_4279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4281 = 8'hb5 == r_count_19_io_out ? io_r_181_b : _GEN_4280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4282 = 8'hb6 == r_count_19_io_out ? io_r_182_b : _GEN_4281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4283 = 8'hb7 == r_count_19_io_out ? io_r_183_b : _GEN_4282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4284 = 8'hb8 == r_count_19_io_out ? io_r_184_b : _GEN_4283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4285 = 8'hb9 == r_count_19_io_out ? io_r_185_b : _GEN_4284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4286 = 8'hba == r_count_19_io_out ? io_r_186_b : _GEN_4285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4287 = 8'hbb == r_count_19_io_out ? io_r_187_b : _GEN_4286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4288 = 8'hbc == r_count_19_io_out ? io_r_188_b : _GEN_4287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4289 = 8'hbd == r_count_19_io_out ? io_r_189_b : _GEN_4288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4290 = 8'hbe == r_count_19_io_out ? io_r_190_b : _GEN_4289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4291 = 8'hbf == r_count_19_io_out ? io_r_191_b : _GEN_4290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4292 = 8'hc0 == r_count_19_io_out ? io_r_192_b : _GEN_4291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4293 = 8'hc1 == r_count_19_io_out ? io_r_193_b : _GEN_4292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4294 = 8'hc2 == r_count_19_io_out ? io_r_194_b : _GEN_4293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4295 = 8'hc3 == r_count_19_io_out ? io_r_195_b : _GEN_4294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4296 = 8'hc4 == r_count_19_io_out ? io_r_196_b : _GEN_4295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4297 = 8'hc5 == r_count_19_io_out ? io_r_197_b : _GEN_4296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4298 = 8'hc6 == r_count_19_io_out ? io_r_198_b : _GEN_4297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4301 = 8'h1 == r_count_20_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4302 = 8'h2 == r_count_20_io_out ? io_r_2_b : _GEN_4301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4303 = 8'h3 == r_count_20_io_out ? io_r_3_b : _GEN_4302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4304 = 8'h4 == r_count_20_io_out ? io_r_4_b : _GEN_4303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4305 = 8'h5 == r_count_20_io_out ? io_r_5_b : _GEN_4304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4306 = 8'h6 == r_count_20_io_out ? io_r_6_b : _GEN_4305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4307 = 8'h7 == r_count_20_io_out ? io_r_7_b : _GEN_4306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4308 = 8'h8 == r_count_20_io_out ? io_r_8_b : _GEN_4307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4309 = 8'h9 == r_count_20_io_out ? io_r_9_b : _GEN_4308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4310 = 8'ha == r_count_20_io_out ? io_r_10_b : _GEN_4309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4311 = 8'hb == r_count_20_io_out ? io_r_11_b : _GEN_4310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4312 = 8'hc == r_count_20_io_out ? io_r_12_b : _GEN_4311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4313 = 8'hd == r_count_20_io_out ? io_r_13_b : _GEN_4312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4314 = 8'he == r_count_20_io_out ? io_r_14_b : _GEN_4313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4315 = 8'hf == r_count_20_io_out ? io_r_15_b : _GEN_4314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4316 = 8'h10 == r_count_20_io_out ? io_r_16_b : _GEN_4315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4317 = 8'h11 == r_count_20_io_out ? io_r_17_b : _GEN_4316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4318 = 8'h12 == r_count_20_io_out ? io_r_18_b : _GEN_4317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4319 = 8'h13 == r_count_20_io_out ? io_r_19_b : _GEN_4318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4320 = 8'h14 == r_count_20_io_out ? io_r_20_b : _GEN_4319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4321 = 8'h15 == r_count_20_io_out ? io_r_21_b : _GEN_4320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4322 = 8'h16 == r_count_20_io_out ? io_r_22_b : _GEN_4321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4323 = 8'h17 == r_count_20_io_out ? io_r_23_b : _GEN_4322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4324 = 8'h18 == r_count_20_io_out ? io_r_24_b : _GEN_4323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4325 = 8'h19 == r_count_20_io_out ? io_r_25_b : _GEN_4324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4326 = 8'h1a == r_count_20_io_out ? io_r_26_b : _GEN_4325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4327 = 8'h1b == r_count_20_io_out ? io_r_27_b : _GEN_4326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4328 = 8'h1c == r_count_20_io_out ? io_r_28_b : _GEN_4327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4329 = 8'h1d == r_count_20_io_out ? io_r_29_b : _GEN_4328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4330 = 8'h1e == r_count_20_io_out ? io_r_30_b : _GEN_4329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4331 = 8'h1f == r_count_20_io_out ? io_r_31_b : _GEN_4330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4332 = 8'h20 == r_count_20_io_out ? io_r_32_b : _GEN_4331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4333 = 8'h21 == r_count_20_io_out ? io_r_33_b : _GEN_4332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4334 = 8'h22 == r_count_20_io_out ? io_r_34_b : _GEN_4333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4335 = 8'h23 == r_count_20_io_out ? io_r_35_b : _GEN_4334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4336 = 8'h24 == r_count_20_io_out ? io_r_36_b : _GEN_4335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4337 = 8'h25 == r_count_20_io_out ? io_r_37_b : _GEN_4336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4338 = 8'h26 == r_count_20_io_out ? io_r_38_b : _GEN_4337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4339 = 8'h27 == r_count_20_io_out ? io_r_39_b : _GEN_4338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4340 = 8'h28 == r_count_20_io_out ? io_r_40_b : _GEN_4339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4341 = 8'h29 == r_count_20_io_out ? io_r_41_b : _GEN_4340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4342 = 8'h2a == r_count_20_io_out ? io_r_42_b : _GEN_4341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4343 = 8'h2b == r_count_20_io_out ? io_r_43_b : _GEN_4342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4344 = 8'h2c == r_count_20_io_out ? io_r_44_b : _GEN_4343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4345 = 8'h2d == r_count_20_io_out ? io_r_45_b : _GEN_4344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4346 = 8'h2e == r_count_20_io_out ? io_r_46_b : _GEN_4345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4347 = 8'h2f == r_count_20_io_out ? io_r_47_b : _GEN_4346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4348 = 8'h30 == r_count_20_io_out ? io_r_48_b : _GEN_4347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4349 = 8'h31 == r_count_20_io_out ? io_r_49_b : _GEN_4348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4350 = 8'h32 == r_count_20_io_out ? io_r_50_b : _GEN_4349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4351 = 8'h33 == r_count_20_io_out ? io_r_51_b : _GEN_4350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4352 = 8'h34 == r_count_20_io_out ? io_r_52_b : _GEN_4351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4353 = 8'h35 == r_count_20_io_out ? io_r_53_b : _GEN_4352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4354 = 8'h36 == r_count_20_io_out ? io_r_54_b : _GEN_4353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4355 = 8'h37 == r_count_20_io_out ? io_r_55_b : _GEN_4354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4356 = 8'h38 == r_count_20_io_out ? io_r_56_b : _GEN_4355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4357 = 8'h39 == r_count_20_io_out ? io_r_57_b : _GEN_4356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4358 = 8'h3a == r_count_20_io_out ? io_r_58_b : _GEN_4357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4359 = 8'h3b == r_count_20_io_out ? io_r_59_b : _GEN_4358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4360 = 8'h3c == r_count_20_io_out ? io_r_60_b : _GEN_4359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4361 = 8'h3d == r_count_20_io_out ? io_r_61_b : _GEN_4360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4362 = 8'h3e == r_count_20_io_out ? io_r_62_b : _GEN_4361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4363 = 8'h3f == r_count_20_io_out ? io_r_63_b : _GEN_4362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4364 = 8'h40 == r_count_20_io_out ? io_r_64_b : _GEN_4363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4365 = 8'h41 == r_count_20_io_out ? io_r_65_b : _GEN_4364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4366 = 8'h42 == r_count_20_io_out ? io_r_66_b : _GEN_4365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4367 = 8'h43 == r_count_20_io_out ? io_r_67_b : _GEN_4366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4368 = 8'h44 == r_count_20_io_out ? io_r_68_b : _GEN_4367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4369 = 8'h45 == r_count_20_io_out ? io_r_69_b : _GEN_4368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4370 = 8'h46 == r_count_20_io_out ? io_r_70_b : _GEN_4369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4371 = 8'h47 == r_count_20_io_out ? io_r_71_b : _GEN_4370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4372 = 8'h48 == r_count_20_io_out ? io_r_72_b : _GEN_4371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4373 = 8'h49 == r_count_20_io_out ? io_r_73_b : _GEN_4372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4374 = 8'h4a == r_count_20_io_out ? io_r_74_b : _GEN_4373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4375 = 8'h4b == r_count_20_io_out ? io_r_75_b : _GEN_4374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4376 = 8'h4c == r_count_20_io_out ? io_r_76_b : _GEN_4375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4377 = 8'h4d == r_count_20_io_out ? io_r_77_b : _GEN_4376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4378 = 8'h4e == r_count_20_io_out ? io_r_78_b : _GEN_4377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4379 = 8'h4f == r_count_20_io_out ? io_r_79_b : _GEN_4378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4380 = 8'h50 == r_count_20_io_out ? io_r_80_b : _GEN_4379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4381 = 8'h51 == r_count_20_io_out ? io_r_81_b : _GEN_4380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4382 = 8'h52 == r_count_20_io_out ? io_r_82_b : _GEN_4381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4383 = 8'h53 == r_count_20_io_out ? io_r_83_b : _GEN_4382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4384 = 8'h54 == r_count_20_io_out ? io_r_84_b : _GEN_4383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4385 = 8'h55 == r_count_20_io_out ? io_r_85_b : _GEN_4384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4386 = 8'h56 == r_count_20_io_out ? io_r_86_b : _GEN_4385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4387 = 8'h57 == r_count_20_io_out ? io_r_87_b : _GEN_4386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4388 = 8'h58 == r_count_20_io_out ? io_r_88_b : _GEN_4387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4389 = 8'h59 == r_count_20_io_out ? io_r_89_b : _GEN_4388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4390 = 8'h5a == r_count_20_io_out ? io_r_90_b : _GEN_4389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4391 = 8'h5b == r_count_20_io_out ? io_r_91_b : _GEN_4390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4392 = 8'h5c == r_count_20_io_out ? io_r_92_b : _GEN_4391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4393 = 8'h5d == r_count_20_io_out ? io_r_93_b : _GEN_4392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4394 = 8'h5e == r_count_20_io_out ? io_r_94_b : _GEN_4393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4395 = 8'h5f == r_count_20_io_out ? io_r_95_b : _GEN_4394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4396 = 8'h60 == r_count_20_io_out ? io_r_96_b : _GEN_4395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4397 = 8'h61 == r_count_20_io_out ? io_r_97_b : _GEN_4396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4398 = 8'h62 == r_count_20_io_out ? io_r_98_b : _GEN_4397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4399 = 8'h63 == r_count_20_io_out ? io_r_99_b : _GEN_4398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4400 = 8'h64 == r_count_20_io_out ? io_r_100_b : _GEN_4399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4401 = 8'h65 == r_count_20_io_out ? io_r_101_b : _GEN_4400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4402 = 8'h66 == r_count_20_io_out ? io_r_102_b : _GEN_4401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4403 = 8'h67 == r_count_20_io_out ? io_r_103_b : _GEN_4402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4404 = 8'h68 == r_count_20_io_out ? io_r_104_b : _GEN_4403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4405 = 8'h69 == r_count_20_io_out ? io_r_105_b : _GEN_4404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4406 = 8'h6a == r_count_20_io_out ? io_r_106_b : _GEN_4405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4407 = 8'h6b == r_count_20_io_out ? io_r_107_b : _GEN_4406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4408 = 8'h6c == r_count_20_io_out ? io_r_108_b : _GEN_4407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4409 = 8'h6d == r_count_20_io_out ? io_r_109_b : _GEN_4408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4410 = 8'h6e == r_count_20_io_out ? io_r_110_b : _GEN_4409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4411 = 8'h6f == r_count_20_io_out ? io_r_111_b : _GEN_4410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4412 = 8'h70 == r_count_20_io_out ? io_r_112_b : _GEN_4411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4413 = 8'h71 == r_count_20_io_out ? io_r_113_b : _GEN_4412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4414 = 8'h72 == r_count_20_io_out ? io_r_114_b : _GEN_4413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4415 = 8'h73 == r_count_20_io_out ? io_r_115_b : _GEN_4414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4416 = 8'h74 == r_count_20_io_out ? io_r_116_b : _GEN_4415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4417 = 8'h75 == r_count_20_io_out ? io_r_117_b : _GEN_4416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4418 = 8'h76 == r_count_20_io_out ? io_r_118_b : _GEN_4417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4419 = 8'h77 == r_count_20_io_out ? io_r_119_b : _GEN_4418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4420 = 8'h78 == r_count_20_io_out ? io_r_120_b : _GEN_4419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4421 = 8'h79 == r_count_20_io_out ? io_r_121_b : _GEN_4420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4422 = 8'h7a == r_count_20_io_out ? io_r_122_b : _GEN_4421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4423 = 8'h7b == r_count_20_io_out ? io_r_123_b : _GEN_4422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4424 = 8'h7c == r_count_20_io_out ? io_r_124_b : _GEN_4423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4425 = 8'h7d == r_count_20_io_out ? io_r_125_b : _GEN_4424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4426 = 8'h7e == r_count_20_io_out ? io_r_126_b : _GEN_4425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4427 = 8'h7f == r_count_20_io_out ? io_r_127_b : _GEN_4426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4428 = 8'h80 == r_count_20_io_out ? io_r_128_b : _GEN_4427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4429 = 8'h81 == r_count_20_io_out ? io_r_129_b : _GEN_4428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4430 = 8'h82 == r_count_20_io_out ? io_r_130_b : _GEN_4429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4431 = 8'h83 == r_count_20_io_out ? io_r_131_b : _GEN_4430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4432 = 8'h84 == r_count_20_io_out ? io_r_132_b : _GEN_4431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4433 = 8'h85 == r_count_20_io_out ? io_r_133_b : _GEN_4432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4434 = 8'h86 == r_count_20_io_out ? io_r_134_b : _GEN_4433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4435 = 8'h87 == r_count_20_io_out ? io_r_135_b : _GEN_4434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4436 = 8'h88 == r_count_20_io_out ? io_r_136_b : _GEN_4435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4437 = 8'h89 == r_count_20_io_out ? io_r_137_b : _GEN_4436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4438 = 8'h8a == r_count_20_io_out ? io_r_138_b : _GEN_4437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4439 = 8'h8b == r_count_20_io_out ? io_r_139_b : _GEN_4438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4440 = 8'h8c == r_count_20_io_out ? io_r_140_b : _GEN_4439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4441 = 8'h8d == r_count_20_io_out ? io_r_141_b : _GEN_4440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4442 = 8'h8e == r_count_20_io_out ? io_r_142_b : _GEN_4441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4443 = 8'h8f == r_count_20_io_out ? io_r_143_b : _GEN_4442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4444 = 8'h90 == r_count_20_io_out ? io_r_144_b : _GEN_4443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4445 = 8'h91 == r_count_20_io_out ? io_r_145_b : _GEN_4444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4446 = 8'h92 == r_count_20_io_out ? io_r_146_b : _GEN_4445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4447 = 8'h93 == r_count_20_io_out ? io_r_147_b : _GEN_4446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4448 = 8'h94 == r_count_20_io_out ? io_r_148_b : _GEN_4447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4449 = 8'h95 == r_count_20_io_out ? io_r_149_b : _GEN_4448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4450 = 8'h96 == r_count_20_io_out ? io_r_150_b : _GEN_4449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4451 = 8'h97 == r_count_20_io_out ? io_r_151_b : _GEN_4450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4452 = 8'h98 == r_count_20_io_out ? io_r_152_b : _GEN_4451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4453 = 8'h99 == r_count_20_io_out ? io_r_153_b : _GEN_4452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4454 = 8'h9a == r_count_20_io_out ? io_r_154_b : _GEN_4453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4455 = 8'h9b == r_count_20_io_out ? io_r_155_b : _GEN_4454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4456 = 8'h9c == r_count_20_io_out ? io_r_156_b : _GEN_4455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4457 = 8'h9d == r_count_20_io_out ? io_r_157_b : _GEN_4456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4458 = 8'h9e == r_count_20_io_out ? io_r_158_b : _GEN_4457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4459 = 8'h9f == r_count_20_io_out ? io_r_159_b : _GEN_4458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4460 = 8'ha0 == r_count_20_io_out ? io_r_160_b : _GEN_4459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4461 = 8'ha1 == r_count_20_io_out ? io_r_161_b : _GEN_4460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4462 = 8'ha2 == r_count_20_io_out ? io_r_162_b : _GEN_4461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4463 = 8'ha3 == r_count_20_io_out ? io_r_163_b : _GEN_4462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4464 = 8'ha4 == r_count_20_io_out ? io_r_164_b : _GEN_4463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4465 = 8'ha5 == r_count_20_io_out ? io_r_165_b : _GEN_4464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4466 = 8'ha6 == r_count_20_io_out ? io_r_166_b : _GEN_4465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4467 = 8'ha7 == r_count_20_io_out ? io_r_167_b : _GEN_4466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4468 = 8'ha8 == r_count_20_io_out ? io_r_168_b : _GEN_4467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4469 = 8'ha9 == r_count_20_io_out ? io_r_169_b : _GEN_4468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4470 = 8'haa == r_count_20_io_out ? io_r_170_b : _GEN_4469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4471 = 8'hab == r_count_20_io_out ? io_r_171_b : _GEN_4470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4472 = 8'hac == r_count_20_io_out ? io_r_172_b : _GEN_4471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4473 = 8'had == r_count_20_io_out ? io_r_173_b : _GEN_4472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4474 = 8'hae == r_count_20_io_out ? io_r_174_b : _GEN_4473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4475 = 8'haf == r_count_20_io_out ? io_r_175_b : _GEN_4474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4476 = 8'hb0 == r_count_20_io_out ? io_r_176_b : _GEN_4475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4477 = 8'hb1 == r_count_20_io_out ? io_r_177_b : _GEN_4476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4478 = 8'hb2 == r_count_20_io_out ? io_r_178_b : _GEN_4477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4479 = 8'hb3 == r_count_20_io_out ? io_r_179_b : _GEN_4478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4480 = 8'hb4 == r_count_20_io_out ? io_r_180_b : _GEN_4479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4481 = 8'hb5 == r_count_20_io_out ? io_r_181_b : _GEN_4480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4482 = 8'hb6 == r_count_20_io_out ? io_r_182_b : _GEN_4481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4483 = 8'hb7 == r_count_20_io_out ? io_r_183_b : _GEN_4482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4484 = 8'hb8 == r_count_20_io_out ? io_r_184_b : _GEN_4483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4485 = 8'hb9 == r_count_20_io_out ? io_r_185_b : _GEN_4484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4486 = 8'hba == r_count_20_io_out ? io_r_186_b : _GEN_4485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4487 = 8'hbb == r_count_20_io_out ? io_r_187_b : _GEN_4486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4488 = 8'hbc == r_count_20_io_out ? io_r_188_b : _GEN_4487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4489 = 8'hbd == r_count_20_io_out ? io_r_189_b : _GEN_4488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4490 = 8'hbe == r_count_20_io_out ? io_r_190_b : _GEN_4489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4491 = 8'hbf == r_count_20_io_out ? io_r_191_b : _GEN_4490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4492 = 8'hc0 == r_count_20_io_out ? io_r_192_b : _GEN_4491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4493 = 8'hc1 == r_count_20_io_out ? io_r_193_b : _GEN_4492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4494 = 8'hc2 == r_count_20_io_out ? io_r_194_b : _GEN_4493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4495 = 8'hc3 == r_count_20_io_out ? io_r_195_b : _GEN_4494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4496 = 8'hc4 == r_count_20_io_out ? io_r_196_b : _GEN_4495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4497 = 8'hc5 == r_count_20_io_out ? io_r_197_b : _GEN_4496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4498 = 8'hc6 == r_count_20_io_out ? io_r_198_b : _GEN_4497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4501 = 8'h1 == r_count_21_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4502 = 8'h2 == r_count_21_io_out ? io_r_2_b : _GEN_4501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4503 = 8'h3 == r_count_21_io_out ? io_r_3_b : _GEN_4502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4504 = 8'h4 == r_count_21_io_out ? io_r_4_b : _GEN_4503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4505 = 8'h5 == r_count_21_io_out ? io_r_5_b : _GEN_4504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4506 = 8'h6 == r_count_21_io_out ? io_r_6_b : _GEN_4505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4507 = 8'h7 == r_count_21_io_out ? io_r_7_b : _GEN_4506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4508 = 8'h8 == r_count_21_io_out ? io_r_8_b : _GEN_4507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4509 = 8'h9 == r_count_21_io_out ? io_r_9_b : _GEN_4508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4510 = 8'ha == r_count_21_io_out ? io_r_10_b : _GEN_4509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4511 = 8'hb == r_count_21_io_out ? io_r_11_b : _GEN_4510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4512 = 8'hc == r_count_21_io_out ? io_r_12_b : _GEN_4511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4513 = 8'hd == r_count_21_io_out ? io_r_13_b : _GEN_4512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4514 = 8'he == r_count_21_io_out ? io_r_14_b : _GEN_4513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4515 = 8'hf == r_count_21_io_out ? io_r_15_b : _GEN_4514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4516 = 8'h10 == r_count_21_io_out ? io_r_16_b : _GEN_4515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4517 = 8'h11 == r_count_21_io_out ? io_r_17_b : _GEN_4516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4518 = 8'h12 == r_count_21_io_out ? io_r_18_b : _GEN_4517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4519 = 8'h13 == r_count_21_io_out ? io_r_19_b : _GEN_4518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4520 = 8'h14 == r_count_21_io_out ? io_r_20_b : _GEN_4519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4521 = 8'h15 == r_count_21_io_out ? io_r_21_b : _GEN_4520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4522 = 8'h16 == r_count_21_io_out ? io_r_22_b : _GEN_4521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4523 = 8'h17 == r_count_21_io_out ? io_r_23_b : _GEN_4522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4524 = 8'h18 == r_count_21_io_out ? io_r_24_b : _GEN_4523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4525 = 8'h19 == r_count_21_io_out ? io_r_25_b : _GEN_4524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4526 = 8'h1a == r_count_21_io_out ? io_r_26_b : _GEN_4525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4527 = 8'h1b == r_count_21_io_out ? io_r_27_b : _GEN_4526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4528 = 8'h1c == r_count_21_io_out ? io_r_28_b : _GEN_4527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4529 = 8'h1d == r_count_21_io_out ? io_r_29_b : _GEN_4528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4530 = 8'h1e == r_count_21_io_out ? io_r_30_b : _GEN_4529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4531 = 8'h1f == r_count_21_io_out ? io_r_31_b : _GEN_4530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4532 = 8'h20 == r_count_21_io_out ? io_r_32_b : _GEN_4531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4533 = 8'h21 == r_count_21_io_out ? io_r_33_b : _GEN_4532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4534 = 8'h22 == r_count_21_io_out ? io_r_34_b : _GEN_4533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4535 = 8'h23 == r_count_21_io_out ? io_r_35_b : _GEN_4534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4536 = 8'h24 == r_count_21_io_out ? io_r_36_b : _GEN_4535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4537 = 8'h25 == r_count_21_io_out ? io_r_37_b : _GEN_4536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4538 = 8'h26 == r_count_21_io_out ? io_r_38_b : _GEN_4537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4539 = 8'h27 == r_count_21_io_out ? io_r_39_b : _GEN_4538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4540 = 8'h28 == r_count_21_io_out ? io_r_40_b : _GEN_4539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4541 = 8'h29 == r_count_21_io_out ? io_r_41_b : _GEN_4540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4542 = 8'h2a == r_count_21_io_out ? io_r_42_b : _GEN_4541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4543 = 8'h2b == r_count_21_io_out ? io_r_43_b : _GEN_4542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4544 = 8'h2c == r_count_21_io_out ? io_r_44_b : _GEN_4543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4545 = 8'h2d == r_count_21_io_out ? io_r_45_b : _GEN_4544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4546 = 8'h2e == r_count_21_io_out ? io_r_46_b : _GEN_4545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4547 = 8'h2f == r_count_21_io_out ? io_r_47_b : _GEN_4546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4548 = 8'h30 == r_count_21_io_out ? io_r_48_b : _GEN_4547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4549 = 8'h31 == r_count_21_io_out ? io_r_49_b : _GEN_4548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4550 = 8'h32 == r_count_21_io_out ? io_r_50_b : _GEN_4549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4551 = 8'h33 == r_count_21_io_out ? io_r_51_b : _GEN_4550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4552 = 8'h34 == r_count_21_io_out ? io_r_52_b : _GEN_4551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4553 = 8'h35 == r_count_21_io_out ? io_r_53_b : _GEN_4552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4554 = 8'h36 == r_count_21_io_out ? io_r_54_b : _GEN_4553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4555 = 8'h37 == r_count_21_io_out ? io_r_55_b : _GEN_4554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4556 = 8'h38 == r_count_21_io_out ? io_r_56_b : _GEN_4555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4557 = 8'h39 == r_count_21_io_out ? io_r_57_b : _GEN_4556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4558 = 8'h3a == r_count_21_io_out ? io_r_58_b : _GEN_4557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4559 = 8'h3b == r_count_21_io_out ? io_r_59_b : _GEN_4558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4560 = 8'h3c == r_count_21_io_out ? io_r_60_b : _GEN_4559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4561 = 8'h3d == r_count_21_io_out ? io_r_61_b : _GEN_4560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4562 = 8'h3e == r_count_21_io_out ? io_r_62_b : _GEN_4561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4563 = 8'h3f == r_count_21_io_out ? io_r_63_b : _GEN_4562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4564 = 8'h40 == r_count_21_io_out ? io_r_64_b : _GEN_4563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4565 = 8'h41 == r_count_21_io_out ? io_r_65_b : _GEN_4564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4566 = 8'h42 == r_count_21_io_out ? io_r_66_b : _GEN_4565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4567 = 8'h43 == r_count_21_io_out ? io_r_67_b : _GEN_4566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4568 = 8'h44 == r_count_21_io_out ? io_r_68_b : _GEN_4567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4569 = 8'h45 == r_count_21_io_out ? io_r_69_b : _GEN_4568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4570 = 8'h46 == r_count_21_io_out ? io_r_70_b : _GEN_4569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4571 = 8'h47 == r_count_21_io_out ? io_r_71_b : _GEN_4570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4572 = 8'h48 == r_count_21_io_out ? io_r_72_b : _GEN_4571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4573 = 8'h49 == r_count_21_io_out ? io_r_73_b : _GEN_4572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4574 = 8'h4a == r_count_21_io_out ? io_r_74_b : _GEN_4573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4575 = 8'h4b == r_count_21_io_out ? io_r_75_b : _GEN_4574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4576 = 8'h4c == r_count_21_io_out ? io_r_76_b : _GEN_4575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4577 = 8'h4d == r_count_21_io_out ? io_r_77_b : _GEN_4576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4578 = 8'h4e == r_count_21_io_out ? io_r_78_b : _GEN_4577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4579 = 8'h4f == r_count_21_io_out ? io_r_79_b : _GEN_4578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4580 = 8'h50 == r_count_21_io_out ? io_r_80_b : _GEN_4579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4581 = 8'h51 == r_count_21_io_out ? io_r_81_b : _GEN_4580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4582 = 8'h52 == r_count_21_io_out ? io_r_82_b : _GEN_4581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4583 = 8'h53 == r_count_21_io_out ? io_r_83_b : _GEN_4582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4584 = 8'h54 == r_count_21_io_out ? io_r_84_b : _GEN_4583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4585 = 8'h55 == r_count_21_io_out ? io_r_85_b : _GEN_4584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4586 = 8'h56 == r_count_21_io_out ? io_r_86_b : _GEN_4585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4587 = 8'h57 == r_count_21_io_out ? io_r_87_b : _GEN_4586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4588 = 8'h58 == r_count_21_io_out ? io_r_88_b : _GEN_4587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4589 = 8'h59 == r_count_21_io_out ? io_r_89_b : _GEN_4588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4590 = 8'h5a == r_count_21_io_out ? io_r_90_b : _GEN_4589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4591 = 8'h5b == r_count_21_io_out ? io_r_91_b : _GEN_4590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4592 = 8'h5c == r_count_21_io_out ? io_r_92_b : _GEN_4591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4593 = 8'h5d == r_count_21_io_out ? io_r_93_b : _GEN_4592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4594 = 8'h5e == r_count_21_io_out ? io_r_94_b : _GEN_4593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4595 = 8'h5f == r_count_21_io_out ? io_r_95_b : _GEN_4594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4596 = 8'h60 == r_count_21_io_out ? io_r_96_b : _GEN_4595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4597 = 8'h61 == r_count_21_io_out ? io_r_97_b : _GEN_4596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4598 = 8'h62 == r_count_21_io_out ? io_r_98_b : _GEN_4597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4599 = 8'h63 == r_count_21_io_out ? io_r_99_b : _GEN_4598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4600 = 8'h64 == r_count_21_io_out ? io_r_100_b : _GEN_4599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4601 = 8'h65 == r_count_21_io_out ? io_r_101_b : _GEN_4600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4602 = 8'h66 == r_count_21_io_out ? io_r_102_b : _GEN_4601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4603 = 8'h67 == r_count_21_io_out ? io_r_103_b : _GEN_4602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4604 = 8'h68 == r_count_21_io_out ? io_r_104_b : _GEN_4603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4605 = 8'h69 == r_count_21_io_out ? io_r_105_b : _GEN_4604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4606 = 8'h6a == r_count_21_io_out ? io_r_106_b : _GEN_4605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4607 = 8'h6b == r_count_21_io_out ? io_r_107_b : _GEN_4606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4608 = 8'h6c == r_count_21_io_out ? io_r_108_b : _GEN_4607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4609 = 8'h6d == r_count_21_io_out ? io_r_109_b : _GEN_4608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4610 = 8'h6e == r_count_21_io_out ? io_r_110_b : _GEN_4609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4611 = 8'h6f == r_count_21_io_out ? io_r_111_b : _GEN_4610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4612 = 8'h70 == r_count_21_io_out ? io_r_112_b : _GEN_4611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4613 = 8'h71 == r_count_21_io_out ? io_r_113_b : _GEN_4612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4614 = 8'h72 == r_count_21_io_out ? io_r_114_b : _GEN_4613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4615 = 8'h73 == r_count_21_io_out ? io_r_115_b : _GEN_4614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4616 = 8'h74 == r_count_21_io_out ? io_r_116_b : _GEN_4615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4617 = 8'h75 == r_count_21_io_out ? io_r_117_b : _GEN_4616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4618 = 8'h76 == r_count_21_io_out ? io_r_118_b : _GEN_4617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4619 = 8'h77 == r_count_21_io_out ? io_r_119_b : _GEN_4618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4620 = 8'h78 == r_count_21_io_out ? io_r_120_b : _GEN_4619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4621 = 8'h79 == r_count_21_io_out ? io_r_121_b : _GEN_4620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4622 = 8'h7a == r_count_21_io_out ? io_r_122_b : _GEN_4621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4623 = 8'h7b == r_count_21_io_out ? io_r_123_b : _GEN_4622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4624 = 8'h7c == r_count_21_io_out ? io_r_124_b : _GEN_4623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4625 = 8'h7d == r_count_21_io_out ? io_r_125_b : _GEN_4624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4626 = 8'h7e == r_count_21_io_out ? io_r_126_b : _GEN_4625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4627 = 8'h7f == r_count_21_io_out ? io_r_127_b : _GEN_4626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4628 = 8'h80 == r_count_21_io_out ? io_r_128_b : _GEN_4627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4629 = 8'h81 == r_count_21_io_out ? io_r_129_b : _GEN_4628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4630 = 8'h82 == r_count_21_io_out ? io_r_130_b : _GEN_4629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4631 = 8'h83 == r_count_21_io_out ? io_r_131_b : _GEN_4630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4632 = 8'h84 == r_count_21_io_out ? io_r_132_b : _GEN_4631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4633 = 8'h85 == r_count_21_io_out ? io_r_133_b : _GEN_4632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4634 = 8'h86 == r_count_21_io_out ? io_r_134_b : _GEN_4633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4635 = 8'h87 == r_count_21_io_out ? io_r_135_b : _GEN_4634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4636 = 8'h88 == r_count_21_io_out ? io_r_136_b : _GEN_4635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4637 = 8'h89 == r_count_21_io_out ? io_r_137_b : _GEN_4636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4638 = 8'h8a == r_count_21_io_out ? io_r_138_b : _GEN_4637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4639 = 8'h8b == r_count_21_io_out ? io_r_139_b : _GEN_4638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4640 = 8'h8c == r_count_21_io_out ? io_r_140_b : _GEN_4639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4641 = 8'h8d == r_count_21_io_out ? io_r_141_b : _GEN_4640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4642 = 8'h8e == r_count_21_io_out ? io_r_142_b : _GEN_4641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4643 = 8'h8f == r_count_21_io_out ? io_r_143_b : _GEN_4642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4644 = 8'h90 == r_count_21_io_out ? io_r_144_b : _GEN_4643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4645 = 8'h91 == r_count_21_io_out ? io_r_145_b : _GEN_4644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4646 = 8'h92 == r_count_21_io_out ? io_r_146_b : _GEN_4645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4647 = 8'h93 == r_count_21_io_out ? io_r_147_b : _GEN_4646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4648 = 8'h94 == r_count_21_io_out ? io_r_148_b : _GEN_4647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4649 = 8'h95 == r_count_21_io_out ? io_r_149_b : _GEN_4648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4650 = 8'h96 == r_count_21_io_out ? io_r_150_b : _GEN_4649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4651 = 8'h97 == r_count_21_io_out ? io_r_151_b : _GEN_4650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4652 = 8'h98 == r_count_21_io_out ? io_r_152_b : _GEN_4651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4653 = 8'h99 == r_count_21_io_out ? io_r_153_b : _GEN_4652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4654 = 8'h9a == r_count_21_io_out ? io_r_154_b : _GEN_4653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4655 = 8'h9b == r_count_21_io_out ? io_r_155_b : _GEN_4654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4656 = 8'h9c == r_count_21_io_out ? io_r_156_b : _GEN_4655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4657 = 8'h9d == r_count_21_io_out ? io_r_157_b : _GEN_4656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4658 = 8'h9e == r_count_21_io_out ? io_r_158_b : _GEN_4657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4659 = 8'h9f == r_count_21_io_out ? io_r_159_b : _GEN_4658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4660 = 8'ha0 == r_count_21_io_out ? io_r_160_b : _GEN_4659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4661 = 8'ha1 == r_count_21_io_out ? io_r_161_b : _GEN_4660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4662 = 8'ha2 == r_count_21_io_out ? io_r_162_b : _GEN_4661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4663 = 8'ha3 == r_count_21_io_out ? io_r_163_b : _GEN_4662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4664 = 8'ha4 == r_count_21_io_out ? io_r_164_b : _GEN_4663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4665 = 8'ha5 == r_count_21_io_out ? io_r_165_b : _GEN_4664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4666 = 8'ha6 == r_count_21_io_out ? io_r_166_b : _GEN_4665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4667 = 8'ha7 == r_count_21_io_out ? io_r_167_b : _GEN_4666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4668 = 8'ha8 == r_count_21_io_out ? io_r_168_b : _GEN_4667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4669 = 8'ha9 == r_count_21_io_out ? io_r_169_b : _GEN_4668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4670 = 8'haa == r_count_21_io_out ? io_r_170_b : _GEN_4669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4671 = 8'hab == r_count_21_io_out ? io_r_171_b : _GEN_4670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4672 = 8'hac == r_count_21_io_out ? io_r_172_b : _GEN_4671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4673 = 8'had == r_count_21_io_out ? io_r_173_b : _GEN_4672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4674 = 8'hae == r_count_21_io_out ? io_r_174_b : _GEN_4673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4675 = 8'haf == r_count_21_io_out ? io_r_175_b : _GEN_4674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4676 = 8'hb0 == r_count_21_io_out ? io_r_176_b : _GEN_4675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4677 = 8'hb1 == r_count_21_io_out ? io_r_177_b : _GEN_4676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4678 = 8'hb2 == r_count_21_io_out ? io_r_178_b : _GEN_4677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4679 = 8'hb3 == r_count_21_io_out ? io_r_179_b : _GEN_4678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4680 = 8'hb4 == r_count_21_io_out ? io_r_180_b : _GEN_4679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4681 = 8'hb5 == r_count_21_io_out ? io_r_181_b : _GEN_4680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4682 = 8'hb6 == r_count_21_io_out ? io_r_182_b : _GEN_4681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4683 = 8'hb7 == r_count_21_io_out ? io_r_183_b : _GEN_4682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4684 = 8'hb8 == r_count_21_io_out ? io_r_184_b : _GEN_4683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4685 = 8'hb9 == r_count_21_io_out ? io_r_185_b : _GEN_4684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4686 = 8'hba == r_count_21_io_out ? io_r_186_b : _GEN_4685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4687 = 8'hbb == r_count_21_io_out ? io_r_187_b : _GEN_4686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4688 = 8'hbc == r_count_21_io_out ? io_r_188_b : _GEN_4687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4689 = 8'hbd == r_count_21_io_out ? io_r_189_b : _GEN_4688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4690 = 8'hbe == r_count_21_io_out ? io_r_190_b : _GEN_4689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4691 = 8'hbf == r_count_21_io_out ? io_r_191_b : _GEN_4690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4692 = 8'hc0 == r_count_21_io_out ? io_r_192_b : _GEN_4691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4693 = 8'hc1 == r_count_21_io_out ? io_r_193_b : _GEN_4692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4694 = 8'hc2 == r_count_21_io_out ? io_r_194_b : _GEN_4693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4695 = 8'hc3 == r_count_21_io_out ? io_r_195_b : _GEN_4694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4696 = 8'hc4 == r_count_21_io_out ? io_r_196_b : _GEN_4695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4697 = 8'hc5 == r_count_21_io_out ? io_r_197_b : _GEN_4696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4698 = 8'hc6 == r_count_21_io_out ? io_r_198_b : _GEN_4697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4701 = 8'h1 == r_count_22_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4702 = 8'h2 == r_count_22_io_out ? io_r_2_b : _GEN_4701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4703 = 8'h3 == r_count_22_io_out ? io_r_3_b : _GEN_4702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4704 = 8'h4 == r_count_22_io_out ? io_r_4_b : _GEN_4703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4705 = 8'h5 == r_count_22_io_out ? io_r_5_b : _GEN_4704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4706 = 8'h6 == r_count_22_io_out ? io_r_6_b : _GEN_4705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4707 = 8'h7 == r_count_22_io_out ? io_r_7_b : _GEN_4706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4708 = 8'h8 == r_count_22_io_out ? io_r_8_b : _GEN_4707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4709 = 8'h9 == r_count_22_io_out ? io_r_9_b : _GEN_4708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4710 = 8'ha == r_count_22_io_out ? io_r_10_b : _GEN_4709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4711 = 8'hb == r_count_22_io_out ? io_r_11_b : _GEN_4710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4712 = 8'hc == r_count_22_io_out ? io_r_12_b : _GEN_4711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4713 = 8'hd == r_count_22_io_out ? io_r_13_b : _GEN_4712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4714 = 8'he == r_count_22_io_out ? io_r_14_b : _GEN_4713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4715 = 8'hf == r_count_22_io_out ? io_r_15_b : _GEN_4714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4716 = 8'h10 == r_count_22_io_out ? io_r_16_b : _GEN_4715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4717 = 8'h11 == r_count_22_io_out ? io_r_17_b : _GEN_4716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4718 = 8'h12 == r_count_22_io_out ? io_r_18_b : _GEN_4717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4719 = 8'h13 == r_count_22_io_out ? io_r_19_b : _GEN_4718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4720 = 8'h14 == r_count_22_io_out ? io_r_20_b : _GEN_4719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4721 = 8'h15 == r_count_22_io_out ? io_r_21_b : _GEN_4720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4722 = 8'h16 == r_count_22_io_out ? io_r_22_b : _GEN_4721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4723 = 8'h17 == r_count_22_io_out ? io_r_23_b : _GEN_4722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4724 = 8'h18 == r_count_22_io_out ? io_r_24_b : _GEN_4723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4725 = 8'h19 == r_count_22_io_out ? io_r_25_b : _GEN_4724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4726 = 8'h1a == r_count_22_io_out ? io_r_26_b : _GEN_4725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4727 = 8'h1b == r_count_22_io_out ? io_r_27_b : _GEN_4726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4728 = 8'h1c == r_count_22_io_out ? io_r_28_b : _GEN_4727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4729 = 8'h1d == r_count_22_io_out ? io_r_29_b : _GEN_4728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4730 = 8'h1e == r_count_22_io_out ? io_r_30_b : _GEN_4729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4731 = 8'h1f == r_count_22_io_out ? io_r_31_b : _GEN_4730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4732 = 8'h20 == r_count_22_io_out ? io_r_32_b : _GEN_4731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4733 = 8'h21 == r_count_22_io_out ? io_r_33_b : _GEN_4732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4734 = 8'h22 == r_count_22_io_out ? io_r_34_b : _GEN_4733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4735 = 8'h23 == r_count_22_io_out ? io_r_35_b : _GEN_4734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4736 = 8'h24 == r_count_22_io_out ? io_r_36_b : _GEN_4735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4737 = 8'h25 == r_count_22_io_out ? io_r_37_b : _GEN_4736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4738 = 8'h26 == r_count_22_io_out ? io_r_38_b : _GEN_4737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4739 = 8'h27 == r_count_22_io_out ? io_r_39_b : _GEN_4738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4740 = 8'h28 == r_count_22_io_out ? io_r_40_b : _GEN_4739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4741 = 8'h29 == r_count_22_io_out ? io_r_41_b : _GEN_4740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4742 = 8'h2a == r_count_22_io_out ? io_r_42_b : _GEN_4741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4743 = 8'h2b == r_count_22_io_out ? io_r_43_b : _GEN_4742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4744 = 8'h2c == r_count_22_io_out ? io_r_44_b : _GEN_4743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4745 = 8'h2d == r_count_22_io_out ? io_r_45_b : _GEN_4744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4746 = 8'h2e == r_count_22_io_out ? io_r_46_b : _GEN_4745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4747 = 8'h2f == r_count_22_io_out ? io_r_47_b : _GEN_4746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4748 = 8'h30 == r_count_22_io_out ? io_r_48_b : _GEN_4747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4749 = 8'h31 == r_count_22_io_out ? io_r_49_b : _GEN_4748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4750 = 8'h32 == r_count_22_io_out ? io_r_50_b : _GEN_4749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4751 = 8'h33 == r_count_22_io_out ? io_r_51_b : _GEN_4750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4752 = 8'h34 == r_count_22_io_out ? io_r_52_b : _GEN_4751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4753 = 8'h35 == r_count_22_io_out ? io_r_53_b : _GEN_4752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4754 = 8'h36 == r_count_22_io_out ? io_r_54_b : _GEN_4753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4755 = 8'h37 == r_count_22_io_out ? io_r_55_b : _GEN_4754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4756 = 8'h38 == r_count_22_io_out ? io_r_56_b : _GEN_4755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4757 = 8'h39 == r_count_22_io_out ? io_r_57_b : _GEN_4756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4758 = 8'h3a == r_count_22_io_out ? io_r_58_b : _GEN_4757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4759 = 8'h3b == r_count_22_io_out ? io_r_59_b : _GEN_4758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4760 = 8'h3c == r_count_22_io_out ? io_r_60_b : _GEN_4759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4761 = 8'h3d == r_count_22_io_out ? io_r_61_b : _GEN_4760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4762 = 8'h3e == r_count_22_io_out ? io_r_62_b : _GEN_4761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4763 = 8'h3f == r_count_22_io_out ? io_r_63_b : _GEN_4762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4764 = 8'h40 == r_count_22_io_out ? io_r_64_b : _GEN_4763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4765 = 8'h41 == r_count_22_io_out ? io_r_65_b : _GEN_4764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4766 = 8'h42 == r_count_22_io_out ? io_r_66_b : _GEN_4765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4767 = 8'h43 == r_count_22_io_out ? io_r_67_b : _GEN_4766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4768 = 8'h44 == r_count_22_io_out ? io_r_68_b : _GEN_4767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4769 = 8'h45 == r_count_22_io_out ? io_r_69_b : _GEN_4768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4770 = 8'h46 == r_count_22_io_out ? io_r_70_b : _GEN_4769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4771 = 8'h47 == r_count_22_io_out ? io_r_71_b : _GEN_4770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4772 = 8'h48 == r_count_22_io_out ? io_r_72_b : _GEN_4771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4773 = 8'h49 == r_count_22_io_out ? io_r_73_b : _GEN_4772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4774 = 8'h4a == r_count_22_io_out ? io_r_74_b : _GEN_4773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4775 = 8'h4b == r_count_22_io_out ? io_r_75_b : _GEN_4774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4776 = 8'h4c == r_count_22_io_out ? io_r_76_b : _GEN_4775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4777 = 8'h4d == r_count_22_io_out ? io_r_77_b : _GEN_4776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4778 = 8'h4e == r_count_22_io_out ? io_r_78_b : _GEN_4777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4779 = 8'h4f == r_count_22_io_out ? io_r_79_b : _GEN_4778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4780 = 8'h50 == r_count_22_io_out ? io_r_80_b : _GEN_4779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4781 = 8'h51 == r_count_22_io_out ? io_r_81_b : _GEN_4780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4782 = 8'h52 == r_count_22_io_out ? io_r_82_b : _GEN_4781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4783 = 8'h53 == r_count_22_io_out ? io_r_83_b : _GEN_4782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4784 = 8'h54 == r_count_22_io_out ? io_r_84_b : _GEN_4783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4785 = 8'h55 == r_count_22_io_out ? io_r_85_b : _GEN_4784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4786 = 8'h56 == r_count_22_io_out ? io_r_86_b : _GEN_4785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4787 = 8'h57 == r_count_22_io_out ? io_r_87_b : _GEN_4786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4788 = 8'h58 == r_count_22_io_out ? io_r_88_b : _GEN_4787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4789 = 8'h59 == r_count_22_io_out ? io_r_89_b : _GEN_4788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4790 = 8'h5a == r_count_22_io_out ? io_r_90_b : _GEN_4789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4791 = 8'h5b == r_count_22_io_out ? io_r_91_b : _GEN_4790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4792 = 8'h5c == r_count_22_io_out ? io_r_92_b : _GEN_4791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4793 = 8'h5d == r_count_22_io_out ? io_r_93_b : _GEN_4792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4794 = 8'h5e == r_count_22_io_out ? io_r_94_b : _GEN_4793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4795 = 8'h5f == r_count_22_io_out ? io_r_95_b : _GEN_4794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4796 = 8'h60 == r_count_22_io_out ? io_r_96_b : _GEN_4795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4797 = 8'h61 == r_count_22_io_out ? io_r_97_b : _GEN_4796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4798 = 8'h62 == r_count_22_io_out ? io_r_98_b : _GEN_4797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4799 = 8'h63 == r_count_22_io_out ? io_r_99_b : _GEN_4798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4800 = 8'h64 == r_count_22_io_out ? io_r_100_b : _GEN_4799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4801 = 8'h65 == r_count_22_io_out ? io_r_101_b : _GEN_4800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4802 = 8'h66 == r_count_22_io_out ? io_r_102_b : _GEN_4801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4803 = 8'h67 == r_count_22_io_out ? io_r_103_b : _GEN_4802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4804 = 8'h68 == r_count_22_io_out ? io_r_104_b : _GEN_4803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4805 = 8'h69 == r_count_22_io_out ? io_r_105_b : _GEN_4804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4806 = 8'h6a == r_count_22_io_out ? io_r_106_b : _GEN_4805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4807 = 8'h6b == r_count_22_io_out ? io_r_107_b : _GEN_4806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4808 = 8'h6c == r_count_22_io_out ? io_r_108_b : _GEN_4807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4809 = 8'h6d == r_count_22_io_out ? io_r_109_b : _GEN_4808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4810 = 8'h6e == r_count_22_io_out ? io_r_110_b : _GEN_4809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4811 = 8'h6f == r_count_22_io_out ? io_r_111_b : _GEN_4810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4812 = 8'h70 == r_count_22_io_out ? io_r_112_b : _GEN_4811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4813 = 8'h71 == r_count_22_io_out ? io_r_113_b : _GEN_4812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4814 = 8'h72 == r_count_22_io_out ? io_r_114_b : _GEN_4813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4815 = 8'h73 == r_count_22_io_out ? io_r_115_b : _GEN_4814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4816 = 8'h74 == r_count_22_io_out ? io_r_116_b : _GEN_4815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4817 = 8'h75 == r_count_22_io_out ? io_r_117_b : _GEN_4816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4818 = 8'h76 == r_count_22_io_out ? io_r_118_b : _GEN_4817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4819 = 8'h77 == r_count_22_io_out ? io_r_119_b : _GEN_4818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4820 = 8'h78 == r_count_22_io_out ? io_r_120_b : _GEN_4819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4821 = 8'h79 == r_count_22_io_out ? io_r_121_b : _GEN_4820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4822 = 8'h7a == r_count_22_io_out ? io_r_122_b : _GEN_4821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4823 = 8'h7b == r_count_22_io_out ? io_r_123_b : _GEN_4822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4824 = 8'h7c == r_count_22_io_out ? io_r_124_b : _GEN_4823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4825 = 8'h7d == r_count_22_io_out ? io_r_125_b : _GEN_4824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4826 = 8'h7e == r_count_22_io_out ? io_r_126_b : _GEN_4825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4827 = 8'h7f == r_count_22_io_out ? io_r_127_b : _GEN_4826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4828 = 8'h80 == r_count_22_io_out ? io_r_128_b : _GEN_4827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4829 = 8'h81 == r_count_22_io_out ? io_r_129_b : _GEN_4828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4830 = 8'h82 == r_count_22_io_out ? io_r_130_b : _GEN_4829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4831 = 8'h83 == r_count_22_io_out ? io_r_131_b : _GEN_4830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4832 = 8'h84 == r_count_22_io_out ? io_r_132_b : _GEN_4831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4833 = 8'h85 == r_count_22_io_out ? io_r_133_b : _GEN_4832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4834 = 8'h86 == r_count_22_io_out ? io_r_134_b : _GEN_4833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4835 = 8'h87 == r_count_22_io_out ? io_r_135_b : _GEN_4834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4836 = 8'h88 == r_count_22_io_out ? io_r_136_b : _GEN_4835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4837 = 8'h89 == r_count_22_io_out ? io_r_137_b : _GEN_4836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4838 = 8'h8a == r_count_22_io_out ? io_r_138_b : _GEN_4837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4839 = 8'h8b == r_count_22_io_out ? io_r_139_b : _GEN_4838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4840 = 8'h8c == r_count_22_io_out ? io_r_140_b : _GEN_4839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4841 = 8'h8d == r_count_22_io_out ? io_r_141_b : _GEN_4840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4842 = 8'h8e == r_count_22_io_out ? io_r_142_b : _GEN_4841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4843 = 8'h8f == r_count_22_io_out ? io_r_143_b : _GEN_4842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4844 = 8'h90 == r_count_22_io_out ? io_r_144_b : _GEN_4843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4845 = 8'h91 == r_count_22_io_out ? io_r_145_b : _GEN_4844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4846 = 8'h92 == r_count_22_io_out ? io_r_146_b : _GEN_4845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4847 = 8'h93 == r_count_22_io_out ? io_r_147_b : _GEN_4846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4848 = 8'h94 == r_count_22_io_out ? io_r_148_b : _GEN_4847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4849 = 8'h95 == r_count_22_io_out ? io_r_149_b : _GEN_4848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4850 = 8'h96 == r_count_22_io_out ? io_r_150_b : _GEN_4849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4851 = 8'h97 == r_count_22_io_out ? io_r_151_b : _GEN_4850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4852 = 8'h98 == r_count_22_io_out ? io_r_152_b : _GEN_4851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4853 = 8'h99 == r_count_22_io_out ? io_r_153_b : _GEN_4852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4854 = 8'h9a == r_count_22_io_out ? io_r_154_b : _GEN_4853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4855 = 8'h9b == r_count_22_io_out ? io_r_155_b : _GEN_4854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4856 = 8'h9c == r_count_22_io_out ? io_r_156_b : _GEN_4855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4857 = 8'h9d == r_count_22_io_out ? io_r_157_b : _GEN_4856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4858 = 8'h9e == r_count_22_io_out ? io_r_158_b : _GEN_4857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4859 = 8'h9f == r_count_22_io_out ? io_r_159_b : _GEN_4858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4860 = 8'ha0 == r_count_22_io_out ? io_r_160_b : _GEN_4859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4861 = 8'ha1 == r_count_22_io_out ? io_r_161_b : _GEN_4860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4862 = 8'ha2 == r_count_22_io_out ? io_r_162_b : _GEN_4861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4863 = 8'ha3 == r_count_22_io_out ? io_r_163_b : _GEN_4862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4864 = 8'ha4 == r_count_22_io_out ? io_r_164_b : _GEN_4863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4865 = 8'ha5 == r_count_22_io_out ? io_r_165_b : _GEN_4864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4866 = 8'ha6 == r_count_22_io_out ? io_r_166_b : _GEN_4865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4867 = 8'ha7 == r_count_22_io_out ? io_r_167_b : _GEN_4866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4868 = 8'ha8 == r_count_22_io_out ? io_r_168_b : _GEN_4867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4869 = 8'ha9 == r_count_22_io_out ? io_r_169_b : _GEN_4868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4870 = 8'haa == r_count_22_io_out ? io_r_170_b : _GEN_4869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4871 = 8'hab == r_count_22_io_out ? io_r_171_b : _GEN_4870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4872 = 8'hac == r_count_22_io_out ? io_r_172_b : _GEN_4871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4873 = 8'had == r_count_22_io_out ? io_r_173_b : _GEN_4872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4874 = 8'hae == r_count_22_io_out ? io_r_174_b : _GEN_4873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4875 = 8'haf == r_count_22_io_out ? io_r_175_b : _GEN_4874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4876 = 8'hb0 == r_count_22_io_out ? io_r_176_b : _GEN_4875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4877 = 8'hb1 == r_count_22_io_out ? io_r_177_b : _GEN_4876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4878 = 8'hb2 == r_count_22_io_out ? io_r_178_b : _GEN_4877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4879 = 8'hb3 == r_count_22_io_out ? io_r_179_b : _GEN_4878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4880 = 8'hb4 == r_count_22_io_out ? io_r_180_b : _GEN_4879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4881 = 8'hb5 == r_count_22_io_out ? io_r_181_b : _GEN_4880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4882 = 8'hb6 == r_count_22_io_out ? io_r_182_b : _GEN_4881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4883 = 8'hb7 == r_count_22_io_out ? io_r_183_b : _GEN_4882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4884 = 8'hb8 == r_count_22_io_out ? io_r_184_b : _GEN_4883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4885 = 8'hb9 == r_count_22_io_out ? io_r_185_b : _GEN_4884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4886 = 8'hba == r_count_22_io_out ? io_r_186_b : _GEN_4885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4887 = 8'hbb == r_count_22_io_out ? io_r_187_b : _GEN_4886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4888 = 8'hbc == r_count_22_io_out ? io_r_188_b : _GEN_4887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4889 = 8'hbd == r_count_22_io_out ? io_r_189_b : _GEN_4888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4890 = 8'hbe == r_count_22_io_out ? io_r_190_b : _GEN_4889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4891 = 8'hbf == r_count_22_io_out ? io_r_191_b : _GEN_4890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4892 = 8'hc0 == r_count_22_io_out ? io_r_192_b : _GEN_4891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4893 = 8'hc1 == r_count_22_io_out ? io_r_193_b : _GEN_4892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4894 = 8'hc2 == r_count_22_io_out ? io_r_194_b : _GEN_4893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4895 = 8'hc3 == r_count_22_io_out ? io_r_195_b : _GEN_4894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4896 = 8'hc4 == r_count_22_io_out ? io_r_196_b : _GEN_4895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4897 = 8'hc5 == r_count_22_io_out ? io_r_197_b : _GEN_4896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4898 = 8'hc6 == r_count_22_io_out ? io_r_198_b : _GEN_4897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4901 = 8'h1 == r_count_23_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4902 = 8'h2 == r_count_23_io_out ? io_r_2_b : _GEN_4901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4903 = 8'h3 == r_count_23_io_out ? io_r_3_b : _GEN_4902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4904 = 8'h4 == r_count_23_io_out ? io_r_4_b : _GEN_4903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4905 = 8'h5 == r_count_23_io_out ? io_r_5_b : _GEN_4904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4906 = 8'h6 == r_count_23_io_out ? io_r_6_b : _GEN_4905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4907 = 8'h7 == r_count_23_io_out ? io_r_7_b : _GEN_4906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4908 = 8'h8 == r_count_23_io_out ? io_r_8_b : _GEN_4907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4909 = 8'h9 == r_count_23_io_out ? io_r_9_b : _GEN_4908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4910 = 8'ha == r_count_23_io_out ? io_r_10_b : _GEN_4909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4911 = 8'hb == r_count_23_io_out ? io_r_11_b : _GEN_4910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4912 = 8'hc == r_count_23_io_out ? io_r_12_b : _GEN_4911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4913 = 8'hd == r_count_23_io_out ? io_r_13_b : _GEN_4912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4914 = 8'he == r_count_23_io_out ? io_r_14_b : _GEN_4913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4915 = 8'hf == r_count_23_io_out ? io_r_15_b : _GEN_4914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4916 = 8'h10 == r_count_23_io_out ? io_r_16_b : _GEN_4915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4917 = 8'h11 == r_count_23_io_out ? io_r_17_b : _GEN_4916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4918 = 8'h12 == r_count_23_io_out ? io_r_18_b : _GEN_4917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4919 = 8'h13 == r_count_23_io_out ? io_r_19_b : _GEN_4918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4920 = 8'h14 == r_count_23_io_out ? io_r_20_b : _GEN_4919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4921 = 8'h15 == r_count_23_io_out ? io_r_21_b : _GEN_4920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4922 = 8'h16 == r_count_23_io_out ? io_r_22_b : _GEN_4921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4923 = 8'h17 == r_count_23_io_out ? io_r_23_b : _GEN_4922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4924 = 8'h18 == r_count_23_io_out ? io_r_24_b : _GEN_4923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4925 = 8'h19 == r_count_23_io_out ? io_r_25_b : _GEN_4924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4926 = 8'h1a == r_count_23_io_out ? io_r_26_b : _GEN_4925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4927 = 8'h1b == r_count_23_io_out ? io_r_27_b : _GEN_4926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4928 = 8'h1c == r_count_23_io_out ? io_r_28_b : _GEN_4927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4929 = 8'h1d == r_count_23_io_out ? io_r_29_b : _GEN_4928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4930 = 8'h1e == r_count_23_io_out ? io_r_30_b : _GEN_4929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4931 = 8'h1f == r_count_23_io_out ? io_r_31_b : _GEN_4930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4932 = 8'h20 == r_count_23_io_out ? io_r_32_b : _GEN_4931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4933 = 8'h21 == r_count_23_io_out ? io_r_33_b : _GEN_4932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4934 = 8'h22 == r_count_23_io_out ? io_r_34_b : _GEN_4933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4935 = 8'h23 == r_count_23_io_out ? io_r_35_b : _GEN_4934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4936 = 8'h24 == r_count_23_io_out ? io_r_36_b : _GEN_4935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4937 = 8'h25 == r_count_23_io_out ? io_r_37_b : _GEN_4936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4938 = 8'h26 == r_count_23_io_out ? io_r_38_b : _GEN_4937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4939 = 8'h27 == r_count_23_io_out ? io_r_39_b : _GEN_4938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4940 = 8'h28 == r_count_23_io_out ? io_r_40_b : _GEN_4939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4941 = 8'h29 == r_count_23_io_out ? io_r_41_b : _GEN_4940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4942 = 8'h2a == r_count_23_io_out ? io_r_42_b : _GEN_4941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4943 = 8'h2b == r_count_23_io_out ? io_r_43_b : _GEN_4942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4944 = 8'h2c == r_count_23_io_out ? io_r_44_b : _GEN_4943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4945 = 8'h2d == r_count_23_io_out ? io_r_45_b : _GEN_4944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4946 = 8'h2e == r_count_23_io_out ? io_r_46_b : _GEN_4945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4947 = 8'h2f == r_count_23_io_out ? io_r_47_b : _GEN_4946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4948 = 8'h30 == r_count_23_io_out ? io_r_48_b : _GEN_4947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4949 = 8'h31 == r_count_23_io_out ? io_r_49_b : _GEN_4948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4950 = 8'h32 == r_count_23_io_out ? io_r_50_b : _GEN_4949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4951 = 8'h33 == r_count_23_io_out ? io_r_51_b : _GEN_4950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4952 = 8'h34 == r_count_23_io_out ? io_r_52_b : _GEN_4951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4953 = 8'h35 == r_count_23_io_out ? io_r_53_b : _GEN_4952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4954 = 8'h36 == r_count_23_io_out ? io_r_54_b : _GEN_4953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4955 = 8'h37 == r_count_23_io_out ? io_r_55_b : _GEN_4954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4956 = 8'h38 == r_count_23_io_out ? io_r_56_b : _GEN_4955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4957 = 8'h39 == r_count_23_io_out ? io_r_57_b : _GEN_4956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4958 = 8'h3a == r_count_23_io_out ? io_r_58_b : _GEN_4957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4959 = 8'h3b == r_count_23_io_out ? io_r_59_b : _GEN_4958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4960 = 8'h3c == r_count_23_io_out ? io_r_60_b : _GEN_4959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4961 = 8'h3d == r_count_23_io_out ? io_r_61_b : _GEN_4960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4962 = 8'h3e == r_count_23_io_out ? io_r_62_b : _GEN_4961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4963 = 8'h3f == r_count_23_io_out ? io_r_63_b : _GEN_4962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4964 = 8'h40 == r_count_23_io_out ? io_r_64_b : _GEN_4963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4965 = 8'h41 == r_count_23_io_out ? io_r_65_b : _GEN_4964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4966 = 8'h42 == r_count_23_io_out ? io_r_66_b : _GEN_4965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4967 = 8'h43 == r_count_23_io_out ? io_r_67_b : _GEN_4966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4968 = 8'h44 == r_count_23_io_out ? io_r_68_b : _GEN_4967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4969 = 8'h45 == r_count_23_io_out ? io_r_69_b : _GEN_4968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4970 = 8'h46 == r_count_23_io_out ? io_r_70_b : _GEN_4969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4971 = 8'h47 == r_count_23_io_out ? io_r_71_b : _GEN_4970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4972 = 8'h48 == r_count_23_io_out ? io_r_72_b : _GEN_4971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4973 = 8'h49 == r_count_23_io_out ? io_r_73_b : _GEN_4972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4974 = 8'h4a == r_count_23_io_out ? io_r_74_b : _GEN_4973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4975 = 8'h4b == r_count_23_io_out ? io_r_75_b : _GEN_4974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4976 = 8'h4c == r_count_23_io_out ? io_r_76_b : _GEN_4975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4977 = 8'h4d == r_count_23_io_out ? io_r_77_b : _GEN_4976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4978 = 8'h4e == r_count_23_io_out ? io_r_78_b : _GEN_4977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4979 = 8'h4f == r_count_23_io_out ? io_r_79_b : _GEN_4978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4980 = 8'h50 == r_count_23_io_out ? io_r_80_b : _GEN_4979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4981 = 8'h51 == r_count_23_io_out ? io_r_81_b : _GEN_4980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4982 = 8'h52 == r_count_23_io_out ? io_r_82_b : _GEN_4981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4983 = 8'h53 == r_count_23_io_out ? io_r_83_b : _GEN_4982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4984 = 8'h54 == r_count_23_io_out ? io_r_84_b : _GEN_4983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4985 = 8'h55 == r_count_23_io_out ? io_r_85_b : _GEN_4984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4986 = 8'h56 == r_count_23_io_out ? io_r_86_b : _GEN_4985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4987 = 8'h57 == r_count_23_io_out ? io_r_87_b : _GEN_4986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4988 = 8'h58 == r_count_23_io_out ? io_r_88_b : _GEN_4987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4989 = 8'h59 == r_count_23_io_out ? io_r_89_b : _GEN_4988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4990 = 8'h5a == r_count_23_io_out ? io_r_90_b : _GEN_4989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4991 = 8'h5b == r_count_23_io_out ? io_r_91_b : _GEN_4990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4992 = 8'h5c == r_count_23_io_out ? io_r_92_b : _GEN_4991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4993 = 8'h5d == r_count_23_io_out ? io_r_93_b : _GEN_4992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4994 = 8'h5e == r_count_23_io_out ? io_r_94_b : _GEN_4993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4995 = 8'h5f == r_count_23_io_out ? io_r_95_b : _GEN_4994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4996 = 8'h60 == r_count_23_io_out ? io_r_96_b : _GEN_4995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4997 = 8'h61 == r_count_23_io_out ? io_r_97_b : _GEN_4996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4998 = 8'h62 == r_count_23_io_out ? io_r_98_b : _GEN_4997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4999 = 8'h63 == r_count_23_io_out ? io_r_99_b : _GEN_4998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5000 = 8'h64 == r_count_23_io_out ? io_r_100_b : _GEN_4999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5001 = 8'h65 == r_count_23_io_out ? io_r_101_b : _GEN_5000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5002 = 8'h66 == r_count_23_io_out ? io_r_102_b : _GEN_5001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5003 = 8'h67 == r_count_23_io_out ? io_r_103_b : _GEN_5002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5004 = 8'h68 == r_count_23_io_out ? io_r_104_b : _GEN_5003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5005 = 8'h69 == r_count_23_io_out ? io_r_105_b : _GEN_5004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5006 = 8'h6a == r_count_23_io_out ? io_r_106_b : _GEN_5005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5007 = 8'h6b == r_count_23_io_out ? io_r_107_b : _GEN_5006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5008 = 8'h6c == r_count_23_io_out ? io_r_108_b : _GEN_5007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5009 = 8'h6d == r_count_23_io_out ? io_r_109_b : _GEN_5008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5010 = 8'h6e == r_count_23_io_out ? io_r_110_b : _GEN_5009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5011 = 8'h6f == r_count_23_io_out ? io_r_111_b : _GEN_5010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5012 = 8'h70 == r_count_23_io_out ? io_r_112_b : _GEN_5011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5013 = 8'h71 == r_count_23_io_out ? io_r_113_b : _GEN_5012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5014 = 8'h72 == r_count_23_io_out ? io_r_114_b : _GEN_5013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5015 = 8'h73 == r_count_23_io_out ? io_r_115_b : _GEN_5014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5016 = 8'h74 == r_count_23_io_out ? io_r_116_b : _GEN_5015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5017 = 8'h75 == r_count_23_io_out ? io_r_117_b : _GEN_5016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5018 = 8'h76 == r_count_23_io_out ? io_r_118_b : _GEN_5017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5019 = 8'h77 == r_count_23_io_out ? io_r_119_b : _GEN_5018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5020 = 8'h78 == r_count_23_io_out ? io_r_120_b : _GEN_5019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5021 = 8'h79 == r_count_23_io_out ? io_r_121_b : _GEN_5020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5022 = 8'h7a == r_count_23_io_out ? io_r_122_b : _GEN_5021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5023 = 8'h7b == r_count_23_io_out ? io_r_123_b : _GEN_5022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5024 = 8'h7c == r_count_23_io_out ? io_r_124_b : _GEN_5023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5025 = 8'h7d == r_count_23_io_out ? io_r_125_b : _GEN_5024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5026 = 8'h7e == r_count_23_io_out ? io_r_126_b : _GEN_5025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5027 = 8'h7f == r_count_23_io_out ? io_r_127_b : _GEN_5026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5028 = 8'h80 == r_count_23_io_out ? io_r_128_b : _GEN_5027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5029 = 8'h81 == r_count_23_io_out ? io_r_129_b : _GEN_5028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5030 = 8'h82 == r_count_23_io_out ? io_r_130_b : _GEN_5029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5031 = 8'h83 == r_count_23_io_out ? io_r_131_b : _GEN_5030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5032 = 8'h84 == r_count_23_io_out ? io_r_132_b : _GEN_5031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5033 = 8'h85 == r_count_23_io_out ? io_r_133_b : _GEN_5032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5034 = 8'h86 == r_count_23_io_out ? io_r_134_b : _GEN_5033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5035 = 8'h87 == r_count_23_io_out ? io_r_135_b : _GEN_5034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5036 = 8'h88 == r_count_23_io_out ? io_r_136_b : _GEN_5035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5037 = 8'h89 == r_count_23_io_out ? io_r_137_b : _GEN_5036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5038 = 8'h8a == r_count_23_io_out ? io_r_138_b : _GEN_5037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5039 = 8'h8b == r_count_23_io_out ? io_r_139_b : _GEN_5038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5040 = 8'h8c == r_count_23_io_out ? io_r_140_b : _GEN_5039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5041 = 8'h8d == r_count_23_io_out ? io_r_141_b : _GEN_5040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5042 = 8'h8e == r_count_23_io_out ? io_r_142_b : _GEN_5041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5043 = 8'h8f == r_count_23_io_out ? io_r_143_b : _GEN_5042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5044 = 8'h90 == r_count_23_io_out ? io_r_144_b : _GEN_5043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5045 = 8'h91 == r_count_23_io_out ? io_r_145_b : _GEN_5044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5046 = 8'h92 == r_count_23_io_out ? io_r_146_b : _GEN_5045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5047 = 8'h93 == r_count_23_io_out ? io_r_147_b : _GEN_5046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5048 = 8'h94 == r_count_23_io_out ? io_r_148_b : _GEN_5047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5049 = 8'h95 == r_count_23_io_out ? io_r_149_b : _GEN_5048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5050 = 8'h96 == r_count_23_io_out ? io_r_150_b : _GEN_5049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5051 = 8'h97 == r_count_23_io_out ? io_r_151_b : _GEN_5050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5052 = 8'h98 == r_count_23_io_out ? io_r_152_b : _GEN_5051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5053 = 8'h99 == r_count_23_io_out ? io_r_153_b : _GEN_5052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5054 = 8'h9a == r_count_23_io_out ? io_r_154_b : _GEN_5053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5055 = 8'h9b == r_count_23_io_out ? io_r_155_b : _GEN_5054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5056 = 8'h9c == r_count_23_io_out ? io_r_156_b : _GEN_5055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5057 = 8'h9d == r_count_23_io_out ? io_r_157_b : _GEN_5056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5058 = 8'h9e == r_count_23_io_out ? io_r_158_b : _GEN_5057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5059 = 8'h9f == r_count_23_io_out ? io_r_159_b : _GEN_5058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5060 = 8'ha0 == r_count_23_io_out ? io_r_160_b : _GEN_5059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5061 = 8'ha1 == r_count_23_io_out ? io_r_161_b : _GEN_5060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5062 = 8'ha2 == r_count_23_io_out ? io_r_162_b : _GEN_5061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5063 = 8'ha3 == r_count_23_io_out ? io_r_163_b : _GEN_5062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5064 = 8'ha4 == r_count_23_io_out ? io_r_164_b : _GEN_5063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5065 = 8'ha5 == r_count_23_io_out ? io_r_165_b : _GEN_5064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5066 = 8'ha6 == r_count_23_io_out ? io_r_166_b : _GEN_5065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5067 = 8'ha7 == r_count_23_io_out ? io_r_167_b : _GEN_5066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5068 = 8'ha8 == r_count_23_io_out ? io_r_168_b : _GEN_5067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5069 = 8'ha9 == r_count_23_io_out ? io_r_169_b : _GEN_5068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5070 = 8'haa == r_count_23_io_out ? io_r_170_b : _GEN_5069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5071 = 8'hab == r_count_23_io_out ? io_r_171_b : _GEN_5070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5072 = 8'hac == r_count_23_io_out ? io_r_172_b : _GEN_5071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5073 = 8'had == r_count_23_io_out ? io_r_173_b : _GEN_5072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5074 = 8'hae == r_count_23_io_out ? io_r_174_b : _GEN_5073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5075 = 8'haf == r_count_23_io_out ? io_r_175_b : _GEN_5074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5076 = 8'hb0 == r_count_23_io_out ? io_r_176_b : _GEN_5075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5077 = 8'hb1 == r_count_23_io_out ? io_r_177_b : _GEN_5076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5078 = 8'hb2 == r_count_23_io_out ? io_r_178_b : _GEN_5077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5079 = 8'hb3 == r_count_23_io_out ? io_r_179_b : _GEN_5078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5080 = 8'hb4 == r_count_23_io_out ? io_r_180_b : _GEN_5079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5081 = 8'hb5 == r_count_23_io_out ? io_r_181_b : _GEN_5080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5082 = 8'hb6 == r_count_23_io_out ? io_r_182_b : _GEN_5081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5083 = 8'hb7 == r_count_23_io_out ? io_r_183_b : _GEN_5082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5084 = 8'hb8 == r_count_23_io_out ? io_r_184_b : _GEN_5083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5085 = 8'hb9 == r_count_23_io_out ? io_r_185_b : _GEN_5084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5086 = 8'hba == r_count_23_io_out ? io_r_186_b : _GEN_5085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5087 = 8'hbb == r_count_23_io_out ? io_r_187_b : _GEN_5086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5088 = 8'hbc == r_count_23_io_out ? io_r_188_b : _GEN_5087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5089 = 8'hbd == r_count_23_io_out ? io_r_189_b : _GEN_5088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5090 = 8'hbe == r_count_23_io_out ? io_r_190_b : _GEN_5089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5091 = 8'hbf == r_count_23_io_out ? io_r_191_b : _GEN_5090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5092 = 8'hc0 == r_count_23_io_out ? io_r_192_b : _GEN_5091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5093 = 8'hc1 == r_count_23_io_out ? io_r_193_b : _GEN_5092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5094 = 8'hc2 == r_count_23_io_out ? io_r_194_b : _GEN_5093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5095 = 8'hc3 == r_count_23_io_out ? io_r_195_b : _GEN_5094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5096 = 8'hc4 == r_count_23_io_out ? io_r_196_b : _GEN_5095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5097 = 8'hc5 == r_count_23_io_out ? io_r_197_b : _GEN_5096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5098 = 8'hc6 == r_count_23_io_out ? io_r_198_b : _GEN_5097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5101 = 8'h1 == r_count_24_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5102 = 8'h2 == r_count_24_io_out ? io_r_2_b : _GEN_5101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5103 = 8'h3 == r_count_24_io_out ? io_r_3_b : _GEN_5102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5104 = 8'h4 == r_count_24_io_out ? io_r_4_b : _GEN_5103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5105 = 8'h5 == r_count_24_io_out ? io_r_5_b : _GEN_5104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5106 = 8'h6 == r_count_24_io_out ? io_r_6_b : _GEN_5105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5107 = 8'h7 == r_count_24_io_out ? io_r_7_b : _GEN_5106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5108 = 8'h8 == r_count_24_io_out ? io_r_8_b : _GEN_5107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5109 = 8'h9 == r_count_24_io_out ? io_r_9_b : _GEN_5108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5110 = 8'ha == r_count_24_io_out ? io_r_10_b : _GEN_5109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5111 = 8'hb == r_count_24_io_out ? io_r_11_b : _GEN_5110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5112 = 8'hc == r_count_24_io_out ? io_r_12_b : _GEN_5111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5113 = 8'hd == r_count_24_io_out ? io_r_13_b : _GEN_5112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5114 = 8'he == r_count_24_io_out ? io_r_14_b : _GEN_5113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5115 = 8'hf == r_count_24_io_out ? io_r_15_b : _GEN_5114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5116 = 8'h10 == r_count_24_io_out ? io_r_16_b : _GEN_5115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5117 = 8'h11 == r_count_24_io_out ? io_r_17_b : _GEN_5116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5118 = 8'h12 == r_count_24_io_out ? io_r_18_b : _GEN_5117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5119 = 8'h13 == r_count_24_io_out ? io_r_19_b : _GEN_5118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5120 = 8'h14 == r_count_24_io_out ? io_r_20_b : _GEN_5119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5121 = 8'h15 == r_count_24_io_out ? io_r_21_b : _GEN_5120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5122 = 8'h16 == r_count_24_io_out ? io_r_22_b : _GEN_5121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5123 = 8'h17 == r_count_24_io_out ? io_r_23_b : _GEN_5122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5124 = 8'h18 == r_count_24_io_out ? io_r_24_b : _GEN_5123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5125 = 8'h19 == r_count_24_io_out ? io_r_25_b : _GEN_5124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5126 = 8'h1a == r_count_24_io_out ? io_r_26_b : _GEN_5125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5127 = 8'h1b == r_count_24_io_out ? io_r_27_b : _GEN_5126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5128 = 8'h1c == r_count_24_io_out ? io_r_28_b : _GEN_5127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5129 = 8'h1d == r_count_24_io_out ? io_r_29_b : _GEN_5128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5130 = 8'h1e == r_count_24_io_out ? io_r_30_b : _GEN_5129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5131 = 8'h1f == r_count_24_io_out ? io_r_31_b : _GEN_5130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5132 = 8'h20 == r_count_24_io_out ? io_r_32_b : _GEN_5131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5133 = 8'h21 == r_count_24_io_out ? io_r_33_b : _GEN_5132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5134 = 8'h22 == r_count_24_io_out ? io_r_34_b : _GEN_5133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5135 = 8'h23 == r_count_24_io_out ? io_r_35_b : _GEN_5134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5136 = 8'h24 == r_count_24_io_out ? io_r_36_b : _GEN_5135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5137 = 8'h25 == r_count_24_io_out ? io_r_37_b : _GEN_5136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5138 = 8'h26 == r_count_24_io_out ? io_r_38_b : _GEN_5137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5139 = 8'h27 == r_count_24_io_out ? io_r_39_b : _GEN_5138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5140 = 8'h28 == r_count_24_io_out ? io_r_40_b : _GEN_5139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5141 = 8'h29 == r_count_24_io_out ? io_r_41_b : _GEN_5140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5142 = 8'h2a == r_count_24_io_out ? io_r_42_b : _GEN_5141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5143 = 8'h2b == r_count_24_io_out ? io_r_43_b : _GEN_5142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5144 = 8'h2c == r_count_24_io_out ? io_r_44_b : _GEN_5143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5145 = 8'h2d == r_count_24_io_out ? io_r_45_b : _GEN_5144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5146 = 8'h2e == r_count_24_io_out ? io_r_46_b : _GEN_5145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5147 = 8'h2f == r_count_24_io_out ? io_r_47_b : _GEN_5146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5148 = 8'h30 == r_count_24_io_out ? io_r_48_b : _GEN_5147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5149 = 8'h31 == r_count_24_io_out ? io_r_49_b : _GEN_5148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5150 = 8'h32 == r_count_24_io_out ? io_r_50_b : _GEN_5149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5151 = 8'h33 == r_count_24_io_out ? io_r_51_b : _GEN_5150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5152 = 8'h34 == r_count_24_io_out ? io_r_52_b : _GEN_5151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5153 = 8'h35 == r_count_24_io_out ? io_r_53_b : _GEN_5152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5154 = 8'h36 == r_count_24_io_out ? io_r_54_b : _GEN_5153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5155 = 8'h37 == r_count_24_io_out ? io_r_55_b : _GEN_5154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5156 = 8'h38 == r_count_24_io_out ? io_r_56_b : _GEN_5155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5157 = 8'h39 == r_count_24_io_out ? io_r_57_b : _GEN_5156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5158 = 8'h3a == r_count_24_io_out ? io_r_58_b : _GEN_5157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5159 = 8'h3b == r_count_24_io_out ? io_r_59_b : _GEN_5158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5160 = 8'h3c == r_count_24_io_out ? io_r_60_b : _GEN_5159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5161 = 8'h3d == r_count_24_io_out ? io_r_61_b : _GEN_5160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5162 = 8'h3e == r_count_24_io_out ? io_r_62_b : _GEN_5161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5163 = 8'h3f == r_count_24_io_out ? io_r_63_b : _GEN_5162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5164 = 8'h40 == r_count_24_io_out ? io_r_64_b : _GEN_5163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5165 = 8'h41 == r_count_24_io_out ? io_r_65_b : _GEN_5164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5166 = 8'h42 == r_count_24_io_out ? io_r_66_b : _GEN_5165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5167 = 8'h43 == r_count_24_io_out ? io_r_67_b : _GEN_5166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5168 = 8'h44 == r_count_24_io_out ? io_r_68_b : _GEN_5167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5169 = 8'h45 == r_count_24_io_out ? io_r_69_b : _GEN_5168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5170 = 8'h46 == r_count_24_io_out ? io_r_70_b : _GEN_5169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5171 = 8'h47 == r_count_24_io_out ? io_r_71_b : _GEN_5170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5172 = 8'h48 == r_count_24_io_out ? io_r_72_b : _GEN_5171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5173 = 8'h49 == r_count_24_io_out ? io_r_73_b : _GEN_5172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5174 = 8'h4a == r_count_24_io_out ? io_r_74_b : _GEN_5173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5175 = 8'h4b == r_count_24_io_out ? io_r_75_b : _GEN_5174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5176 = 8'h4c == r_count_24_io_out ? io_r_76_b : _GEN_5175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5177 = 8'h4d == r_count_24_io_out ? io_r_77_b : _GEN_5176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5178 = 8'h4e == r_count_24_io_out ? io_r_78_b : _GEN_5177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5179 = 8'h4f == r_count_24_io_out ? io_r_79_b : _GEN_5178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5180 = 8'h50 == r_count_24_io_out ? io_r_80_b : _GEN_5179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5181 = 8'h51 == r_count_24_io_out ? io_r_81_b : _GEN_5180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5182 = 8'h52 == r_count_24_io_out ? io_r_82_b : _GEN_5181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5183 = 8'h53 == r_count_24_io_out ? io_r_83_b : _GEN_5182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5184 = 8'h54 == r_count_24_io_out ? io_r_84_b : _GEN_5183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5185 = 8'h55 == r_count_24_io_out ? io_r_85_b : _GEN_5184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5186 = 8'h56 == r_count_24_io_out ? io_r_86_b : _GEN_5185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5187 = 8'h57 == r_count_24_io_out ? io_r_87_b : _GEN_5186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5188 = 8'h58 == r_count_24_io_out ? io_r_88_b : _GEN_5187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5189 = 8'h59 == r_count_24_io_out ? io_r_89_b : _GEN_5188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5190 = 8'h5a == r_count_24_io_out ? io_r_90_b : _GEN_5189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5191 = 8'h5b == r_count_24_io_out ? io_r_91_b : _GEN_5190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5192 = 8'h5c == r_count_24_io_out ? io_r_92_b : _GEN_5191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5193 = 8'h5d == r_count_24_io_out ? io_r_93_b : _GEN_5192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5194 = 8'h5e == r_count_24_io_out ? io_r_94_b : _GEN_5193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5195 = 8'h5f == r_count_24_io_out ? io_r_95_b : _GEN_5194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5196 = 8'h60 == r_count_24_io_out ? io_r_96_b : _GEN_5195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5197 = 8'h61 == r_count_24_io_out ? io_r_97_b : _GEN_5196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5198 = 8'h62 == r_count_24_io_out ? io_r_98_b : _GEN_5197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5199 = 8'h63 == r_count_24_io_out ? io_r_99_b : _GEN_5198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5200 = 8'h64 == r_count_24_io_out ? io_r_100_b : _GEN_5199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5201 = 8'h65 == r_count_24_io_out ? io_r_101_b : _GEN_5200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5202 = 8'h66 == r_count_24_io_out ? io_r_102_b : _GEN_5201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5203 = 8'h67 == r_count_24_io_out ? io_r_103_b : _GEN_5202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5204 = 8'h68 == r_count_24_io_out ? io_r_104_b : _GEN_5203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5205 = 8'h69 == r_count_24_io_out ? io_r_105_b : _GEN_5204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5206 = 8'h6a == r_count_24_io_out ? io_r_106_b : _GEN_5205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5207 = 8'h6b == r_count_24_io_out ? io_r_107_b : _GEN_5206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5208 = 8'h6c == r_count_24_io_out ? io_r_108_b : _GEN_5207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5209 = 8'h6d == r_count_24_io_out ? io_r_109_b : _GEN_5208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5210 = 8'h6e == r_count_24_io_out ? io_r_110_b : _GEN_5209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5211 = 8'h6f == r_count_24_io_out ? io_r_111_b : _GEN_5210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5212 = 8'h70 == r_count_24_io_out ? io_r_112_b : _GEN_5211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5213 = 8'h71 == r_count_24_io_out ? io_r_113_b : _GEN_5212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5214 = 8'h72 == r_count_24_io_out ? io_r_114_b : _GEN_5213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5215 = 8'h73 == r_count_24_io_out ? io_r_115_b : _GEN_5214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5216 = 8'h74 == r_count_24_io_out ? io_r_116_b : _GEN_5215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5217 = 8'h75 == r_count_24_io_out ? io_r_117_b : _GEN_5216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5218 = 8'h76 == r_count_24_io_out ? io_r_118_b : _GEN_5217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5219 = 8'h77 == r_count_24_io_out ? io_r_119_b : _GEN_5218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5220 = 8'h78 == r_count_24_io_out ? io_r_120_b : _GEN_5219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5221 = 8'h79 == r_count_24_io_out ? io_r_121_b : _GEN_5220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5222 = 8'h7a == r_count_24_io_out ? io_r_122_b : _GEN_5221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5223 = 8'h7b == r_count_24_io_out ? io_r_123_b : _GEN_5222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5224 = 8'h7c == r_count_24_io_out ? io_r_124_b : _GEN_5223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5225 = 8'h7d == r_count_24_io_out ? io_r_125_b : _GEN_5224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5226 = 8'h7e == r_count_24_io_out ? io_r_126_b : _GEN_5225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5227 = 8'h7f == r_count_24_io_out ? io_r_127_b : _GEN_5226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5228 = 8'h80 == r_count_24_io_out ? io_r_128_b : _GEN_5227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5229 = 8'h81 == r_count_24_io_out ? io_r_129_b : _GEN_5228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5230 = 8'h82 == r_count_24_io_out ? io_r_130_b : _GEN_5229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5231 = 8'h83 == r_count_24_io_out ? io_r_131_b : _GEN_5230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5232 = 8'h84 == r_count_24_io_out ? io_r_132_b : _GEN_5231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5233 = 8'h85 == r_count_24_io_out ? io_r_133_b : _GEN_5232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5234 = 8'h86 == r_count_24_io_out ? io_r_134_b : _GEN_5233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5235 = 8'h87 == r_count_24_io_out ? io_r_135_b : _GEN_5234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5236 = 8'h88 == r_count_24_io_out ? io_r_136_b : _GEN_5235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5237 = 8'h89 == r_count_24_io_out ? io_r_137_b : _GEN_5236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5238 = 8'h8a == r_count_24_io_out ? io_r_138_b : _GEN_5237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5239 = 8'h8b == r_count_24_io_out ? io_r_139_b : _GEN_5238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5240 = 8'h8c == r_count_24_io_out ? io_r_140_b : _GEN_5239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5241 = 8'h8d == r_count_24_io_out ? io_r_141_b : _GEN_5240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5242 = 8'h8e == r_count_24_io_out ? io_r_142_b : _GEN_5241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5243 = 8'h8f == r_count_24_io_out ? io_r_143_b : _GEN_5242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5244 = 8'h90 == r_count_24_io_out ? io_r_144_b : _GEN_5243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5245 = 8'h91 == r_count_24_io_out ? io_r_145_b : _GEN_5244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5246 = 8'h92 == r_count_24_io_out ? io_r_146_b : _GEN_5245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5247 = 8'h93 == r_count_24_io_out ? io_r_147_b : _GEN_5246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5248 = 8'h94 == r_count_24_io_out ? io_r_148_b : _GEN_5247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5249 = 8'h95 == r_count_24_io_out ? io_r_149_b : _GEN_5248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5250 = 8'h96 == r_count_24_io_out ? io_r_150_b : _GEN_5249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5251 = 8'h97 == r_count_24_io_out ? io_r_151_b : _GEN_5250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5252 = 8'h98 == r_count_24_io_out ? io_r_152_b : _GEN_5251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5253 = 8'h99 == r_count_24_io_out ? io_r_153_b : _GEN_5252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5254 = 8'h9a == r_count_24_io_out ? io_r_154_b : _GEN_5253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5255 = 8'h9b == r_count_24_io_out ? io_r_155_b : _GEN_5254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5256 = 8'h9c == r_count_24_io_out ? io_r_156_b : _GEN_5255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5257 = 8'h9d == r_count_24_io_out ? io_r_157_b : _GEN_5256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5258 = 8'h9e == r_count_24_io_out ? io_r_158_b : _GEN_5257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5259 = 8'h9f == r_count_24_io_out ? io_r_159_b : _GEN_5258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5260 = 8'ha0 == r_count_24_io_out ? io_r_160_b : _GEN_5259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5261 = 8'ha1 == r_count_24_io_out ? io_r_161_b : _GEN_5260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5262 = 8'ha2 == r_count_24_io_out ? io_r_162_b : _GEN_5261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5263 = 8'ha3 == r_count_24_io_out ? io_r_163_b : _GEN_5262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5264 = 8'ha4 == r_count_24_io_out ? io_r_164_b : _GEN_5263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5265 = 8'ha5 == r_count_24_io_out ? io_r_165_b : _GEN_5264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5266 = 8'ha6 == r_count_24_io_out ? io_r_166_b : _GEN_5265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5267 = 8'ha7 == r_count_24_io_out ? io_r_167_b : _GEN_5266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5268 = 8'ha8 == r_count_24_io_out ? io_r_168_b : _GEN_5267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5269 = 8'ha9 == r_count_24_io_out ? io_r_169_b : _GEN_5268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5270 = 8'haa == r_count_24_io_out ? io_r_170_b : _GEN_5269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5271 = 8'hab == r_count_24_io_out ? io_r_171_b : _GEN_5270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5272 = 8'hac == r_count_24_io_out ? io_r_172_b : _GEN_5271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5273 = 8'had == r_count_24_io_out ? io_r_173_b : _GEN_5272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5274 = 8'hae == r_count_24_io_out ? io_r_174_b : _GEN_5273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5275 = 8'haf == r_count_24_io_out ? io_r_175_b : _GEN_5274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5276 = 8'hb0 == r_count_24_io_out ? io_r_176_b : _GEN_5275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5277 = 8'hb1 == r_count_24_io_out ? io_r_177_b : _GEN_5276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5278 = 8'hb2 == r_count_24_io_out ? io_r_178_b : _GEN_5277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5279 = 8'hb3 == r_count_24_io_out ? io_r_179_b : _GEN_5278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5280 = 8'hb4 == r_count_24_io_out ? io_r_180_b : _GEN_5279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5281 = 8'hb5 == r_count_24_io_out ? io_r_181_b : _GEN_5280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5282 = 8'hb6 == r_count_24_io_out ? io_r_182_b : _GEN_5281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5283 = 8'hb7 == r_count_24_io_out ? io_r_183_b : _GEN_5282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5284 = 8'hb8 == r_count_24_io_out ? io_r_184_b : _GEN_5283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5285 = 8'hb9 == r_count_24_io_out ? io_r_185_b : _GEN_5284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5286 = 8'hba == r_count_24_io_out ? io_r_186_b : _GEN_5285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5287 = 8'hbb == r_count_24_io_out ? io_r_187_b : _GEN_5286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5288 = 8'hbc == r_count_24_io_out ? io_r_188_b : _GEN_5287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5289 = 8'hbd == r_count_24_io_out ? io_r_189_b : _GEN_5288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5290 = 8'hbe == r_count_24_io_out ? io_r_190_b : _GEN_5289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5291 = 8'hbf == r_count_24_io_out ? io_r_191_b : _GEN_5290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5292 = 8'hc0 == r_count_24_io_out ? io_r_192_b : _GEN_5291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5293 = 8'hc1 == r_count_24_io_out ? io_r_193_b : _GEN_5292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5294 = 8'hc2 == r_count_24_io_out ? io_r_194_b : _GEN_5293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5295 = 8'hc3 == r_count_24_io_out ? io_r_195_b : _GEN_5294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5296 = 8'hc4 == r_count_24_io_out ? io_r_196_b : _GEN_5295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5297 = 8'hc5 == r_count_24_io_out ? io_r_197_b : _GEN_5296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5298 = 8'hc6 == r_count_24_io_out ? io_r_198_b : _GEN_5297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5301 = 8'h1 == r_count_25_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5302 = 8'h2 == r_count_25_io_out ? io_r_2_b : _GEN_5301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5303 = 8'h3 == r_count_25_io_out ? io_r_3_b : _GEN_5302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5304 = 8'h4 == r_count_25_io_out ? io_r_4_b : _GEN_5303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5305 = 8'h5 == r_count_25_io_out ? io_r_5_b : _GEN_5304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5306 = 8'h6 == r_count_25_io_out ? io_r_6_b : _GEN_5305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5307 = 8'h7 == r_count_25_io_out ? io_r_7_b : _GEN_5306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5308 = 8'h8 == r_count_25_io_out ? io_r_8_b : _GEN_5307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5309 = 8'h9 == r_count_25_io_out ? io_r_9_b : _GEN_5308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5310 = 8'ha == r_count_25_io_out ? io_r_10_b : _GEN_5309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5311 = 8'hb == r_count_25_io_out ? io_r_11_b : _GEN_5310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5312 = 8'hc == r_count_25_io_out ? io_r_12_b : _GEN_5311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5313 = 8'hd == r_count_25_io_out ? io_r_13_b : _GEN_5312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5314 = 8'he == r_count_25_io_out ? io_r_14_b : _GEN_5313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5315 = 8'hf == r_count_25_io_out ? io_r_15_b : _GEN_5314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5316 = 8'h10 == r_count_25_io_out ? io_r_16_b : _GEN_5315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5317 = 8'h11 == r_count_25_io_out ? io_r_17_b : _GEN_5316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5318 = 8'h12 == r_count_25_io_out ? io_r_18_b : _GEN_5317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5319 = 8'h13 == r_count_25_io_out ? io_r_19_b : _GEN_5318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5320 = 8'h14 == r_count_25_io_out ? io_r_20_b : _GEN_5319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5321 = 8'h15 == r_count_25_io_out ? io_r_21_b : _GEN_5320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5322 = 8'h16 == r_count_25_io_out ? io_r_22_b : _GEN_5321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5323 = 8'h17 == r_count_25_io_out ? io_r_23_b : _GEN_5322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5324 = 8'h18 == r_count_25_io_out ? io_r_24_b : _GEN_5323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5325 = 8'h19 == r_count_25_io_out ? io_r_25_b : _GEN_5324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5326 = 8'h1a == r_count_25_io_out ? io_r_26_b : _GEN_5325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5327 = 8'h1b == r_count_25_io_out ? io_r_27_b : _GEN_5326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5328 = 8'h1c == r_count_25_io_out ? io_r_28_b : _GEN_5327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5329 = 8'h1d == r_count_25_io_out ? io_r_29_b : _GEN_5328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5330 = 8'h1e == r_count_25_io_out ? io_r_30_b : _GEN_5329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5331 = 8'h1f == r_count_25_io_out ? io_r_31_b : _GEN_5330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5332 = 8'h20 == r_count_25_io_out ? io_r_32_b : _GEN_5331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5333 = 8'h21 == r_count_25_io_out ? io_r_33_b : _GEN_5332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5334 = 8'h22 == r_count_25_io_out ? io_r_34_b : _GEN_5333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5335 = 8'h23 == r_count_25_io_out ? io_r_35_b : _GEN_5334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5336 = 8'h24 == r_count_25_io_out ? io_r_36_b : _GEN_5335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5337 = 8'h25 == r_count_25_io_out ? io_r_37_b : _GEN_5336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5338 = 8'h26 == r_count_25_io_out ? io_r_38_b : _GEN_5337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5339 = 8'h27 == r_count_25_io_out ? io_r_39_b : _GEN_5338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5340 = 8'h28 == r_count_25_io_out ? io_r_40_b : _GEN_5339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5341 = 8'h29 == r_count_25_io_out ? io_r_41_b : _GEN_5340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5342 = 8'h2a == r_count_25_io_out ? io_r_42_b : _GEN_5341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5343 = 8'h2b == r_count_25_io_out ? io_r_43_b : _GEN_5342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5344 = 8'h2c == r_count_25_io_out ? io_r_44_b : _GEN_5343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5345 = 8'h2d == r_count_25_io_out ? io_r_45_b : _GEN_5344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5346 = 8'h2e == r_count_25_io_out ? io_r_46_b : _GEN_5345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5347 = 8'h2f == r_count_25_io_out ? io_r_47_b : _GEN_5346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5348 = 8'h30 == r_count_25_io_out ? io_r_48_b : _GEN_5347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5349 = 8'h31 == r_count_25_io_out ? io_r_49_b : _GEN_5348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5350 = 8'h32 == r_count_25_io_out ? io_r_50_b : _GEN_5349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5351 = 8'h33 == r_count_25_io_out ? io_r_51_b : _GEN_5350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5352 = 8'h34 == r_count_25_io_out ? io_r_52_b : _GEN_5351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5353 = 8'h35 == r_count_25_io_out ? io_r_53_b : _GEN_5352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5354 = 8'h36 == r_count_25_io_out ? io_r_54_b : _GEN_5353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5355 = 8'h37 == r_count_25_io_out ? io_r_55_b : _GEN_5354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5356 = 8'h38 == r_count_25_io_out ? io_r_56_b : _GEN_5355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5357 = 8'h39 == r_count_25_io_out ? io_r_57_b : _GEN_5356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5358 = 8'h3a == r_count_25_io_out ? io_r_58_b : _GEN_5357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5359 = 8'h3b == r_count_25_io_out ? io_r_59_b : _GEN_5358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5360 = 8'h3c == r_count_25_io_out ? io_r_60_b : _GEN_5359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5361 = 8'h3d == r_count_25_io_out ? io_r_61_b : _GEN_5360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5362 = 8'h3e == r_count_25_io_out ? io_r_62_b : _GEN_5361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5363 = 8'h3f == r_count_25_io_out ? io_r_63_b : _GEN_5362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5364 = 8'h40 == r_count_25_io_out ? io_r_64_b : _GEN_5363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5365 = 8'h41 == r_count_25_io_out ? io_r_65_b : _GEN_5364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5366 = 8'h42 == r_count_25_io_out ? io_r_66_b : _GEN_5365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5367 = 8'h43 == r_count_25_io_out ? io_r_67_b : _GEN_5366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5368 = 8'h44 == r_count_25_io_out ? io_r_68_b : _GEN_5367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5369 = 8'h45 == r_count_25_io_out ? io_r_69_b : _GEN_5368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5370 = 8'h46 == r_count_25_io_out ? io_r_70_b : _GEN_5369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5371 = 8'h47 == r_count_25_io_out ? io_r_71_b : _GEN_5370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5372 = 8'h48 == r_count_25_io_out ? io_r_72_b : _GEN_5371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5373 = 8'h49 == r_count_25_io_out ? io_r_73_b : _GEN_5372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5374 = 8'h4a == r_count_25_io_out ? io_r_74_b : _GEN_5373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5375 = 8'h4b == r_count_25_io_out ? io_r_75_b : _GEN_5374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5376 = 8'h4c == r_count_25_io_out ? io_r_76_b : _GEN_5375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5377 = 8'h4d == r_count_25_io_out ? io_r_77_b : _GEN_5376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5378 = 8'h4e == r_count_25_io_out ? io_r_78_b : _GEN_5377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5379 = 8'h4f == r_count_25_io_out ? io_r_79_b : _GEN_5378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5380 = 8'h50 == r_count_25_io_out ? io_r_80_b : _GEN_5379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5381 = 8'h51 == r_count_25_io_out ? io_r_81_b : _GEN_5380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5382 = 8'h52 == r_count_25_io_out ? io_r_82_b : _GEN_5381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5383 = 8'h53 == r_count_25_io_out ? io_r_83_b : _GEN_5382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5384 = 8'h54 == r_count_25_io_out ? io_r_84_b : _GEN_5383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5385 = 8'h55 == r_count_25_io_out ? io_r_85_b : _GEN_5384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5386 = 8'h56 == r_count_25_io_out ? io_r_86_b : _GEN_5385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5387 = 8'h57 == r_count_25_io_out ? io_r_87_b : _GEN_5386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5388 = 8'h58 == r_count_25_io_out ? io_r_88_b : _GEN_5387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5389 = 8'h59 == r_count_25_io_out ? io_r_89_b : _GEN_5388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5390 = 8'h5a == r_count_25_io_out ? io_r_90_b : _GEN_5389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5391 = 8'h5b == r_count_25_io_out ? io_r_91_b : _GEN_5390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5392 = 8'h5c == r_count_25_io_out ? io_r_92_b : _GEN_5391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5393 = 8'h5d == r_count_25_io_out ? io_r_93_b : _GEN_5392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5394 = 8'h5e == r_count_25_io_out ? io_r_94_b : _GEN_5393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5395 = 8'h5f == r_count_25_io_out ? io_r_95_b : _GEN_5394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5396 = 8'h60 == r_count_25_io_out ? io_r_96_b : _GEN_5395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5397 = 8'h61 == r_count_25_io_out ? io_r_97_b : _GEN_5396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5398 = 8'h62 == r_count_25_io_out ? io_r_98_b : _GEN_5397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5399 = 8'h63 == r_count_25_io_out ? io_r_99_b : _GEN_5398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5400 = 8'h64 == r_count_25_io_out ? io_r_100_b : _GEN_5399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5401 = 8'h65 == r_count_25_io_out ? io_r_101_b : _GEN_5400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5402 = 8'h66 == r_count_25_io_out ? io_r_102_b : _GEN_5401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5403 = 8'h67 == r_count_25_io_out ? io_r_103_b : _GEN_5402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5404 = 8'h68 == r_count_25_io_out ? io_r_104_b : _GEN_5403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5405 = 8'h69 == r_count_25_io_out ? io_r_105_b : _GEN_5404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5406 = 8'h6a == r_count_25_io_out ? io_r_106_b : _GEN_5405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5407 = 8'h6b == r_count_25_io_out ? io_r_107_b : _GEN_5406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5408 = 8'h6c == r_count_25_io_out ? io_r_108_b : _GEN_5407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5409 = 8'h6d == r_count_25_io_out ? io_r_109_b : _GEN_5408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5410 = 8'h6e == r_count_25_io_out ? io_r_110_b : _GEN_5409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5411 = 8'h6f == r_count_25_io_out ? io_r_111_b : _GEN_5410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5412 = 8'h70 == r_count_25_io_out ? io_r_112_b : _GEN_5411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5413 = 8'h71 == r_count_25_io_out ? io_r_113_b : _GEN_5412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5414 = 8'h72 == r_count_25_io_out ? io_r_114_b : _GEN_5413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5415 = 8'h73 == r_count_25_io_out ? io_r_115_b : _GEN_5414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5416 = 8'h74 == r_count_25_io_out ? io_r_116_b : _GEN_5415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5417 = 8'h75 == r_count_25_io_out ? io_r_117_b : _GEN_5416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5418 = 8'h76 == r_count_25_io_out ? io_r_118_b : _GEN_5417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5419 = 8'h77 == r_count_25_io_out ? io_r_119_b : _GEN_5418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5420 = 8'h78 == r_count_25_io_out ? io_r_120_b : _GEN_5419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5421 = 8'h79 == r_count_25_io_out ? io_r_121_b : _GEN_5420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5422 = 8'h7a == r_count_25_io_out ? io_r_122_b : _GEN_5421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5423 = 8'h7b == r_count_25_io_out ? io_r_123_b : _GEN_5422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5424 = 8'h7c == r_count_25_io_out ? io_r_124_b : _GEN_5423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5425 = 8'h7d == r_count_25_io_out ? io_r_125_b : _GEN_5424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5426 = 8'h7e == r_count_25_io_out ? io_r_126_b : _GEN_5425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5427 = 8'h7f == r_count_25_io_out ? io_r_127_b : _GEN_5426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5428 = 8'h80 == r_count_25_io_out ? io_r_128_b : _GEN_5427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5429 = 8'h81 == r_count_25_io_out ? io_r_129_b : _GEN_5428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5430 = 8'h82 == r_count_25_io_out ? io_r_130_b : _GEN_5429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5431 = 8'h83 == r_count_25_io_out ? io_r_131_b : _GEN_5430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5432 = 8'h84 == r_count_25_io_out ? io_r_132_b : _GEN_5431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5433 = 8'h85 == r_count_25_io_out ? io_r_133_b : _GEN_5432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5434 = 8'h86 == r_count_25_io_out ? io_r_134_b : _GEN_5433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5435 = 8'h87 == r_count_25_io_out ? io_r_135_b : _GEN_5434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5436 = 8'h88 == r_count_25_io_out ? io_r_136_b : _GEN_5435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5437 = 8'h89 == r_count_25_io_out ? io_r_137_b : _GEN_5436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5438 = 8'h8a == r_count_25_io_out ? io_r_138_b : _GEN_5437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5439 = 8'h8b == r_count_25_io_out ? io_r_139_b : _GEN_5438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5440 = 8'h8c == r_count_25_io_out ? io_r_140_b : _GEN_5439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5441 = 8'h8d == r_count_25_io_out ? io_r_141_b : _GEN_5440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5442 = 8'h8e == r_count_25_io_out ? io_r_142_b : _GEN_5441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5443 = 8'h8f == r_count_25_io_out ? io_r_143_b : _GEN_5442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5444 = 8'h90 == r_count_25_io_out ? io_r_144_b : _GEN_5443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5445 = 8'h91 == r_count_25_io_out ? io_r_145_b : _GEN_5444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5446 = 8'h92 == r_count_25_io_out ? io_r_146_b : _GEN_5445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5447 = 8'h93 == r_count_25_io_out ? io_r_147_b : _GEN_5446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5448 = 8'h94 == r_count_25_io_out ? io_r_148_b : _GEN_5447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5449 = 8'h95 == r_count_25_io_out ? io_r_149_b : _GEN_5448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5450 = 8'h96 == r_count_25_io_out ? io_r_150_b : _GEN_5449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5451 = 8'h97 == r_count_25_io_out ? io_r_151_b : _GEN_5450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5452 = 8'h98 == r_count_25_io_out ? io_r_152_b : _GEN_5451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5453 = 8'h99 == r_count_25_io_out ? io_r_153_b : _GEN_5452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5454 = 8'h9a == r_count_25_io_out ? io_r_154_b : _GEN_5453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5455 = 8'h9b == r_count_25_io_out ? io_r_155_b : _GEN_5454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5456 = 8'h9c == r_count_25_io_out ? io_r_156_b : _GEN_5455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5457 = 8'h9d == r_count_25_io_out ? io_r_157_b : _GEN_5456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5458 = 8'h9e == r_count_25_io_out ? io_r_158_b : _GEN_5457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5459 = 8'h9f == r_count_25_io_out ? io_r_159_b : _GEN_5458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5460 = 8'ha0 == r_count_25_io_out ? io_r_160_b : _GEN_5459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5461 = 8'ha1 == r_count_25_io_out ? io_r_161_b : _GEN_5460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5462 = 8'ha2 == r_count_25_io_out ? io_r_162_b : _GEN_5461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5463 = 8'ha3 == r_count_25_io_out ? io_r_163_b : _GEN_5462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5464 = 8'ha4 == r_count_25_io_out ? io_r_164_b : _GEN_5463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5465 = 8'ha5 == r_count_25_io_out ? io_r_165_b : _GEN_5464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5466 = 8'ha6 == r_count_25_io_out ? io_r_166_b : _GEN_5465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5467 = 8'ha7 == r_count_25_io_out ? io_r_167_b : _GEN_5466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5468 = 8'ha8 == r_count_25_io_out ? io_r_168_b : _GEN_5467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5469 = 8'ha9 == r_count_25_io_out ? io_r_169_b : _GEN_5468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5470 = 8'haa == r_count_25_io_out ? io_r_170_b : _GEN_5469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5471 = 8'hab == r_count_25_io_out ? io_r_171_b : _GEN_5470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5472 = 8'hac == r_count_25_io_out ? io_r_172_b : _GEN_5471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5473 = 8'had == r_count_25_io_out ? io_r_173_b : _GEN_5472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5474 = 8'hae == r_count_25_io_out ? io_r_174_b : _GEN_5473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5475 = 8'haf == r_count_25_io_out ? io_r_175_b : _GEN_5474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5476 = 8'hb0 == r_count_25_io_out ? io_r_176_b : _GEN_5475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5477 = 8'hb1 == r_count_25_io_out ? io_r_177_b : _GEN_5476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5478 = 8'hb2 == r_count_25_io_out ? io_r_178_b : _GEN_5477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5479 = 8'hb3 == r_count_25_io_out ? io_r_179_b : _GEN_5478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5480 = 8'hb4 == r_count_25_io_out ? io_r_180_b : _GEN_5479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5481 = 8'hb5 == r_count_25_io_out ? io_r_181_b : _GEN_5480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5482 = 8'hb6 == r_count_25_io_out ? io_r_182_b : _GEN_5481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5483 = 8'hb7 == r_count_25_io_out ? io_r_183_b : _GEN_5482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5484 = 8'hb8 == r_count_25_io_out ? io_r_184_b : _GEN_5483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5485 = 8'hb9 == r_count_25_io_out ? io_r_185_b : _GEN_5484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5486 = 8'hba == r_count_25_io_out ? io_r_186_b : _GEN_5485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5487 = 8'hbb == r_count_25_io_out ? io_r_187_b : _GEN_5486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5488 = 8'hbc == r_count_25_io_out ? io_r_188_b : _GEN_5487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5489 = 8'hbd == r_count_25_io_out ? io_r_189_b : _GEN_5488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5490 = 8'hbe == r_count_25_io_out ? io_r_190_b : _GEN_5489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5491 = 8'hbf == r_count_25_io_out ? io_r_191_b : _GEN_5490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5492 = 8'hc0 == r_count_25_io_out ? io_r_192_b : _GEN_5491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5493 = 8'hc1 == r_count_25_io_out ? io_r_193_b : _GEN_5492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5494 = 8'hc2 == r_count_25_io_out ? io_r_194_b : _GEN_5493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5495 = 8'hc3 == r_count_25_io_out ? io_r_195_b : _GEN_5494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5496 = 8'hc4 == r_count_25_io_out ? io_r_196_b : _GEN_5495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5497 = 8'hc5 == r_count_25_io_out ? io_r_197_b : _GEN_5496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5498 = 8'hc6 == r_count_25_io_out ? io_r_198_b : _GEN_5497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5501 = 8'h1 == r_count_26_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5502 = 8'h2 == r_count_26_io_out ? io_r_2_b : _GEN_5501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5503 = 8'h3 == r_count_26_io_out ? io_r_3_b : _GEN_5502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5504 = 8'h4 == r_count_26_io_out ? io_r_4_b : _GEN_5503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5505 = 8'h5 == r_count_26_io_out ? io_r_5_b : _GEN_5504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5506 = 8'h6 == r_count_26_io_out ? io_r_6_b : _GEN_5505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5507 = 8'h7 == r_count_26_io_out ? io_r_7_b : _GEN_5506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5508 = 8'h8 == r_count_26_io_out ? io_r_8_b : _GEN_5507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5509 = 8'h9 == r_count_26_io_out ? io_r_9_b : _GEN_5508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5510 = 8'ha == r_count_26_io_out ? io_r_10_b : _GEN_5509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5511 = 8'hb == r_count_26_io_out ? io_r_11_b : _GEN_5510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5512 = 8'hc == r_count_26_io_out ? io_r_12_b : _GEN_5511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5513 = 8'hd == r_count_26_io_out ? io_r_13_b : _GEN_5512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5514 = 8'he == r_count_26_io_out ? io_r_14_b : _GEN_5513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5515 = 8'hf == r_count_26_io_out ? io_r_15_b : _GEN_5514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5516 = 8'h10 == r_count_26_io_out ? io_r_16_b : _GEN_5515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5517 = 8'h11 == r_count_26_io_out ? io_r_17_b : _GEN_5516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5518 = 8'h12 == r_count_26_io_out ? io_r_18_b : _GEN_5517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5519 = 8'h13 == r_count_26_io_out ? io_r_19_b : _GEN_5518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5520 = 8'h14 == r_count_26_io_out ? io_r_20_b : _GEN_5519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5521 = 8'h15 == r_count_26_io_out ? io_r_21_b : _GEN_5520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5522 = 8'h16 == r_count_26_io_out ? io_r_22_b : _GEN_5521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5523 = 8'h17 == r_count_26_io_out ? io_r_23_b : _GEN_5522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5524 = 8'h18 == r_count_26_io_out ? io_r_24_b : _GEN_5523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5525 = 8'h19 == r_count_26_io_out ? io_r_25_b : _GEN_5524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5526 = 8'h1a == r_count_26_io_out ? io_r_26_b : _GEN_5525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5527 = 8'h1b == r_count_26_io_out ? io_r_27_b : _GEN_5526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5528 = 8'h1c == r_count_26_io_out ? io_r_28_b : _GEN_5527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5529 = 8'h1d == r_count_26_io_out ? io_r_29_b : _GEN_5528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5530 = 8'h1e == r_count_26_io_out ? io_r_30_b : _GEN_5529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5531 = 8'h1f == r_count_26_io_out ? io_r_31_b : _GEN_5530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5532 = 8'h20 == r_count_26_io_out ? io_r_32_b : _GEN_5531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5533 = 8'h21 == r_count_26_io_out ? io_r_33_b : _GEN_5532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5534 = 8'h22 == r_count_26_io_out ? io_r_34_b : _GEN_5533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5535 = 8'h23 == r_count_26_io_out ? io_r_35_b : _GEN_5534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5536 = 8'h24 == r_count_26_io_out ? io_r_36_b : _GEN_5535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5537 = 8'h25 == r_count_26_io_out ? io_r_37_b : _GEN_5536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5538 = 8'h26 == r_count_26_io_out ? io_r_38_b : _GEN_5537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5539 = 8'h27 == r_count_26_io_out ? io_r_39_b : _GEN_5538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5540 = 8'h28 == r_count_26_io_out ? io_r_40_b : _GEN_5539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5541 = 8'h29 == r_count_26_io_out ? io_r_41_b : _GEN_5540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5542 = 8'h2a == r_count_26_io_out ? io_r_42_b : _GEN_5541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5543 = 8'h2b == r_count_26_io_out ? io_r_43_b : _GEN_5542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5544 = 8'h2c == r_count_26_io_out ? io_r_44_b : _GEN_5543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5545 = 8'h2d == r_count_26_io_out ? io_r_45_b : _GEN_5544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5546 = 8'h2e == r_count_26_io_out ? io_r_46_b : _GEN_5545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5547 = 8'h2f == r_count_26_io_out ? io_r_47_b : _GEN_5546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5548 = 8'h30 == r_count_26_io_out ? io_r_48_b : _GEN_5547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5549 = 8'h31 == r_count_26_io_out ? io_r_49_b : _GEN_5548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5550 = 8'h32 == r_count_26_io_out ? io_r_50_b : _GEN_5549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5551 = 8'h33 == r_count_26_io_out ? io_r_51_b : _GEN_5550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5552 = 8'h34 == r_count_26_io_out ? io_r_52_b : _GEN_5551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5553 = 8'h35 == r_count_26_io_out ? io_r_53_b : _GEN_5552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5554 = 8'h36 == r_count_26_io_out ? io_r_54_b : _GEN_5553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5555 = 8'h37 == r_count_26_io_out ? io_r_55_b : _GEN_5554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5556 = 8'h38 == r_count_26_io_out ? io_r_56_b : _GEN_5555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5557 = 8'h39 == r_count_26_io_out ? io_r_57_b : _GEN_5556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5558 = 8'h3a == r_count_26_io_out ? io_r_58_b : _GEN_5557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5559 = 8'h3b == r_count_26_io_out ? io_r_59_b : _GEN_5558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5560 = 8'h3c == r_count_26_io_out ? io_r_60_b : _GEN_5559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5561 = 8'h3d == r_count_26_io_out ? io_r_61_b : _GEN_5560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5562 = 8'h3e == r_count_26_io_out ? io_r_62_b : _GEN_5561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5563 = 8'h3f == r_count_26_io_out ? io_r_63_b : _GEN_5562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5564 = 8'h40 == r_count_26_io_out ? io_r_64_b : _GEN_5563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5565 = 8'h41 == r_count_26_io_out ? io_r_65_b : _GEN_5564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5566 = 8'h42 == r_count_26_io_out ? io_r_66_b : _GEN_5565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5567 = 8'h43 == r_count_26_io_out ? io_r_67_b : _GEN_5566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5568 = 8'h44 == r_count_26_io_out ? io_r_68_b : _GEN_5567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5569 = 8'h45 == r_count_26_io_out ? io_r_69_b : _GEN_5568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5570 = 8'h46 == r_count_26_io_out ? io_r_70_b : _GEN_5569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5571 = 8'h47 == r_count_26_io_out ? io_r_71_b : _GEN_5570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5572 = 8'h48 == r_count_26_io_out ? io_r_72_b : _GEN_5571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5573 = 8'h49 == r_count_26_io_out ? io_r_73_b : _GEN_5572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5574 = 8'h4a == r_count_26_io_out ? io_r_74_b : _GEN_5573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5575 = 8'h4b == r_count_26_io_out ? io_r_75_b : _GEN_5574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5576 = 8'h4c == r_count_26_io_out ? io_r_76_b : _GEN_5575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5577 = 8'h4d == r_count_26_io_out ? io_r_77_b : _GEN_5576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5578 = 8'h4e == r_count_26_io_out ? io_r_78_b : _GEN_5577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5579 = 8'h4f == r_count_26_io_out ? io_r_79_b : _GEN_5578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5580 = 8'h50 == r_count_26_io_out ? io_r_80_b : _GEN_5579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5581 = 8'h51 == r_count_26_io_out ? io_r_81_b : _GEN_5580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5582 = 8'h52 == r_count_26_io_out ? io_r_82_b : _GEN_5581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5583 = 8'h53 == r_count_26_io_out ? io_r_83_b : _GEN_5582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5584 = 8'h54 == r_count_26_io_out ? io_r_84_b : _GEN_5583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5585 = 8'h55 == r_count_26_io_out ? io_r_85_b : _GEN_5584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5586 = 8'h56 == r_count_26_io_out ? io_r_86_b : _GEN_5585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5587 = 8'h57 == r_count_26_io_out ? io_r_87_b : _GEN_5586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5588 = 8'h58 == r_count_26_io_out ? io_r_88_b : _GEN_5587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5589 = 8'h59 == r_count_26_io_out ? io_r_89_b : _GEN_5588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5590 = 8'h5a == r_count_26_io_out ? io_r_90_b : _GEN_5589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5591 = 8'h5b == r_count_26_io_out ? io_r_91_b : _GEN_5590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5592 = 8'h5c == r_count_26_io_out ? io_r_92_b : _GEN_5591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5593 = 8'h5d == r_count_26_io_out ? io_r_93_b : _GEN_5592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5594 = 8'h5e == r_count_26_io_out ? io_r_94_b : _GEN_5593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5595 = 8'h5f == r_count_26_io_out ? io_r_95_b : _GEN_5594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5596 = 8'h60 == r_count_26_io_out ? io_r_96_b : _GEN_5595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5597 = 8'h61 == r_count_26_io_out ? io_r_97_b : _GEN_5596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5598 = 8'h62 == r_count_26_io_out ? io_r_98_b : _GEN_5597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5599 = 8'h63 == r_count_26_io_out ? io_r_99_b : _GEN_5598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5600 = 8'h64 == r_count_26_io_out ? io_r_100_b : _GEN_5599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5601 = 8'h65 == r_count_26_io_out ? io_r_101_b : _GEN_5600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5602 = 8'h66 == r_count_26_io_out ? io_r_102_b : _GEN_5601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5603 = 8'h67 == r_count_26_io_out ? io_r_103_b : _GEN_5602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5604 = 8'h68 == r_count_26_io_out ? io_r_104_b : _GEN_5603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5605 = 8'h69 == r_count_26_io_out ? io_r_105_b : _GEN_5604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5606 = 8'h6a == r_count_26_io_out ? io_r_106_b : _GEN_5605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5607 = 8'h6b == r_count_26_io_out ? io_r_107_b : _GEN_5606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5608 = 8'h6c == r_count_26_io_out ? io_r_108_b : _GEN_5607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5609 = 8'h6d == r_count_26_io_out ? io_r_109_b : _GEN_5608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5610 = 8'h6e == r_count_26_io_out ? io_r_110_b : _GEN_5609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5611 = 8'h6f == r_count_26_io_out ? io_r_111_b : _GEN_5610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5612 = 8'h70 == r_count_26_io_out ? io_r_112_b : _GEN_5611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5613 = 8'h71 == r_count_26_io_out ? io_r_113_b : _GEN_5612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5614 = 8'h72 == r_count_26_io_out ? io_r_114_b : _GEN_5613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5615 = 8'h73 == r_count_26_io_out ? io_r_115_b : _GEN_5614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5616 = 8'h74 == r_count_26_io_out ? io_r_116_b : _GEN_5615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5617 = 8'h75 == r_count_26_io_out ? io_r_117_b : _GEN_5616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5618 = 8'h76 == r_count_26_io_out ? io_r_118_b : _GEN_5617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5619 = 8'h77 == r_count_26_io_out ? io_r_119_b : _GEN_5618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5620 = 8'h78 == r_count_26_io_out ? io_r_120_b : _GEN_5619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5621 = 8'h79 == r_count_26_io_out ? io_r_121_b : _GEN_5620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5622 = 8'h7a == r_count_26_io_out ? io_r_122_b : _GEN_5621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5623 = 8'h7b == r_count_26_io_out ? io_r_123_b : _GEN_5622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5624 = 8'h7c == r_count_26_io_out ? io_r_124_b : _GEN_5623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5625 = 8'h7d == r_count_26_io_out ? io_r_125_b : _GEN_5624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5626 = 8'h7e == r_count_26_io_out ? io_r_126_b : _GEN_5625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5627 = 8'h7f == r_count_26_io_out ? io_r_127_b : _GEN_5626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5628 = 8'h80 == r_count_26_io_out ? io_r_128_b : _GEN_5627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5629 = 8'h81 == r_count_26_io_out ? io_r_129_b : _GEN_5628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5630 = 8'h82 == r_count_26_io_out ? io_r_130_b : _GEN_5629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5631 = 8'h83 == r_count_26_io_out ? io_r_131_b : _GEN_5630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5632 = 8'h84 == r_count_26_io_out ? io_r_132_b : _GEN_5631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5633 = 8'h85 == r_count_26_io_out ? io_r_133_b : _GEN_5632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5634 = 8'h86 == r_count_26_io_out ? io_r_134_b : _GEN_5633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5635 = 8'h87 == r_count_26_io_out ? io_r_135_b : _GEN_5634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5636 = 8'h88 == r_count_26_io_out ? io_r_136_b : _GEN_5635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5637 = 8'h89 == r_count_26_io_out ? io_r_137_b : _GEN_5636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5638 = 8'h8a == r_count_26_io_out ? io_r_138_b : _GEN_5637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5639 = 8'h8b == r_count_26_io_out ? io_r_139_b : _GEN_5638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5640 = 8'h8c == r_count_26_io_out ? io_r_140_b : _GEN_5639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5641 = 8'h8d == r_count_26_io_out ? io_r_141_b : _GEN_5640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5642 = 8'h8e == r_count_26_io_out ? io_r_142_b : _GEN_5641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5643 = 8'h8f == r_count_26_io_out ? io_r_143_b : _GEN_5642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5644 = 8'h90 == r_count_26_io_out ? io_r_144_b : _GEN_5643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5645 = 8'h91 == r_count_26_io_out ? io_r_145_b : _GEN_5644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5646 = 8'h92 == r_count_26_io_out ? io_r_146_b : _GEN_5645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5647 = 8'h93 == r_count_26_io_out ? io_r_147_b : _GEN_5646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5648 = 8'h94 == r_count_26_io_out ? io_r_148_b : _GEN_5647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5649 = 8'h95 == r_count_26_io_out ? io_r_149_b : _GEN_5648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5650 = 8'h96 == r_count_26_io_out ? io_r_150_b : _GEN_5649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5651 = 8'h97 == r_count_26_io_out ? io_r_151_b : _GEN_5650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5652 = 8'h98 == r_count_26_io_out ? io_r_152_b : _GEN_5651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5653 = 8'h99 == r_count_26_io_out ? io_r_153_b : _GEN_5652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5654 = 8'h9a == r_count_26_io_out ? io_r_154_b : _GEN_5653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5655 = 8'h9b == r_count_26_io_out ? io_r_155_b : _GEN_5654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5656 = 8'h9c == r_count_26_io_out ? io_r_156_b : _GEN_5655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5657 = 8'h9d == r_count_26_io_out ? io_r_157_b : _GEN_5656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5658 = 8'h9e == r_count_26_io_out ? io_r_158_b : _GEN_5657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5659 = 8'h9f == r_count_26_io_out ? io_r_159_b : _GEN_5658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5660 = 8'ha0 == r_count_26_io_out ? io_r_160_b : _GEN_5659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5661 = 8'ha1 == r_count_26_io_out ? io_r_161_b : _GEN_5660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5662 = 8'ha2 == r_count_26_io_out ? io_r_162_b : _GEN_5661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5663 = 8'ha3 == r_count_26_io_out ? io_r_163_b : _GEN_5662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5664 = 8'ha4 == r_count_26_io_out ? io_r_164_b : _GEN_5663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5665 = 8'ha5 == r_count_26_io_out ? io_r_165_b : _GEN_5664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5666 = 8'ha6 == r_count_26_io_out ? io_r_166_b : _GEN_5665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5667 = 8'ha7 == r_count_26_io_out ? io_r_167_b : _GEN_5666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5668 = 8'ha8 == r_count_26_io_out ? io_r_168_b : _GEN_5667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5669 = 8'ha9 == r_count_26_io_out ? io_r_169_b : _GEN_5668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5670 = 8'haa == r_count_26_io_out ? io_r_170_b : _GEN_5669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5671 = 8'hab == r_count_26_io_out ? io_r_171_b : _GEN_5670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5672 = 8'hac == r_count_26_io_out ? io_r_172_b : _GEN_5671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5673 = 8'had == r_count_26_io_out ? io_r_173_b : _GEN_5672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5674 = 8'hae == r_count_26_io_out ? io_r_174_b : _GEN_5673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5675 = 8'haf == r_count_26_io_out ? io_r_175_b : _GEN_5674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5676 = 8'hb0 == r_count_26_io_out ? io_r_176_b : _GEN_5675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5677 = 8'hb1 == r_count_26_io_out ? io_r_177_b : _GEN_5676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5678 = 8'hb2 == r_count_26_io_out ? io_r_178_b : _GEN_5677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5679 = 8'hb3 == r_count_26_io_out ? io_r_179_b : _GEN_5678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5680 = 8'hb4 == r_count_26_io_out ? io_r_180_b : _GEN_5679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5681 = 8'hb5 == r_count_26_io_out ? io_r_181_b : _GEN_5680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5682 = 8'hb6 == r_count_26_io_out ? io_r_182_b : _GEN_5681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5683 = 8'hb7 == r_count_26_io_out ? io_r_183_b : _GEN_5682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5684 = 8'hb8 == r_count_26_io_out ? io_r_184_b : _GEN_5683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5685 = 8'hb9 == r_count_26_io_out ? io_r_185_b : _GEN_5684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5686 = 8'hba == r_count_26_io_out ? io_r_186_b : _GEN_5685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5687 = 8'hbb == r_count_26_io_out ? io_r_187_b : _GEN_5686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5688 = 8'hbc == r_count_26_io_out ? io_r_188_b : _GEN_5687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5689 = 8'hbd == r_count_26_io_out ? io_r_189_b : _GEN_5688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5690 = 8'hbe == r_count_26_io_out ? io_r_190_b : _GEN_5689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5691 = 8'hbf == r_count_26_io_out ? io_r_191_b : _GEN_5690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5692 = 8'hc0 == r_count_26_io_out ? io_r_192_b : _GEN_5691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5693 = 8'hc1 == r_count_26_io_out ? io_r_193_b : _GEN_5692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5694 = 8'hc2 == r_count_26_io_out ? io_r_194_b : _GEN_5693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5695 = 8'hc3 == r_count_26_io_out ? io_r_195_b : _GEN_5694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5696 = 8'hc4 == r_count_26_io_out ? io_r_196_b : _GEN_5695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5697 = 8'hc5 == r_count_26_io_out ? io_r_197_b : _GEN_5696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5698 = 8'hc6 == r_count_26_io_out ? io_r_198_b : _GEN_5697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5701 = 8'h1 == r_count_27_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5702 = 8'h2 == r_count_27_io_out ? io_r_2_b : _GEN_5701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5703 = 8'h3 == r_count_27_io_out ? io_r_3_b : _GEN_5702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5704 = 8'h4 == r_count_27_io_out ? io_r_4_b : _GEN_5703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5705 = 8'h5 == r_count_27_io_out ? io_r_5_b : _GEN_5704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5706 = 8'h6 == r_count_27_io_out ? io_r_6_b : _GEN_5705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5707 = 8'h7 == r_count_27_io_out ? io_r_7_b : _GEN_5706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5708 = 8'h8 == r_count_27_io_out ? io_r_8_b : _GEN_5707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5709 = 8'h9 == r_count_27_io_out ? io_r_9_b : _GEN_5708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5710 = 8'ha == r_count_27_io_out ? io_r_10_b : _GEN_5709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5711 = 8'hb == r_count_27_io_out ? io_r_11_b : _GEN_5710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5712 = 8'hc == r_count_27_io_out ? io_r_12_b : _GEN_5711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5713 = 8'hd == r_count_27_io_out ? io_r_13_b : _GEN_5712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5714 = 8'he == r_count_27_io_out ? io_r_14_b : _GEN_5713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5715 = 8'hf == r_count_27_io_out ? io_r_15_b : _GEN_5714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5716 = 8'h10 == r_count_27_io_out ? io_r_16_b : _GEN_5715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5717 = 8'h11 == r_count_27_io_out ? io_r_17_b : _GEN_5716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5718 = 8'h12 == r_count_27_io_out ? io_r_18_b : _GEN_5717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5719 = 8'h13 == r_count_27_io_out ? io_r_19_b : _GEN_5718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5720 = 8'h14 == r_count_27_io_out ? io_r_20_b : _GEN_5719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5721 = 8'h15 == r_count_27_io_out ? io_r_21_b : _GEN_5720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5722 = 8'h16 == r_count_27_io_out ? io_r_22_b : _GEN_5721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5723 = 8'h17 == r_count_27_io_out ? io_r_23_b : _GEN_5722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5724 = 8'h18 == r_count_27_io_out ? io_r_24_b : _GEN_5723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5725 = 8'h19 == r_count_27_io_out ? io_r_25_b : _GEN_5724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5726 = 8'h1a == r_count_27_io_out ? io_r_26_b : _GEN_5725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5727 = 8'h1b == r_count_27_io_out ? io_r_27_b : _GEN_5726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5728 = 8'h1c == r_count_27_io_out ? io_r_28_b : _GEN_5727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5729 = 8'h1d == r_count_27_io_out ? io_r_29_b : _GEN_5728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5730 = 8'h1e == r_count_27_io_out ? io_r_30_b : _GEN_5729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5731 = 8'h1f == r_count_27_io_out ? io_r_31_b : _GEN_5730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5732 = 8'h20 == r_count_27_io_out ? io_r_32_b : _GEN_5731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5733 = 8'h21 == r_count_27_io_out ? io_r_33_b : _GEN_5732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5734 = 8'h22 == r_count_27_io_out ? io_r_34_b : _GEN_5733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5735 = 8'h23 == r_count_27_io_out ? io_r_35_b : _GEN_5734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5736 = 8'h24 == r_count_27_io_out ? io_r_36_b : _GEN_5735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5737 = 8'h25 == r_count_27_io_out ? io_r_37_b : _GEN_5736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5738 = 8'h26 == r_count_27_io_out ? io_r_38_b : _GEN_5737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5739 = 8'h27 == r_count_27_io_out ? io_r_39_b : _GEN_5738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5740 = 8'h28 == r_count_27_io_out ? io_r_40_b : _GEN_5739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5741 = 8'h29 == r_count_27_io_out ? io_r_41_b : _GEN_5740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5742 = 8'h2a == r_count_27_io_out ? io_r_42_b : _GEN_5741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5743 = 8'h2b == r_count_27_io_out ? io_r_43_b : _GEN_5742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5744 = 8'h2c == r_count_27_io_out ? io_r_44_b : _GEN_5743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5745 = 8'h2d == r_count_27_io_out ? io_r_45_b : _GEN_5744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5746 = 8'h2e == r_count_27_io_out ? io_r_46_b : _GEN_5745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5747 = 8'h2f == r_count_27_io_out ? io_r_47_b : _GEN_5746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5748 = 8'h30 == r_count_27_io_out ? io_r_48_b : _GEN_5747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5749 = 8'h31 == r_count_27_io_out ? io_r_49_b : _GEN_5748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5750 = 8'h32 == r_count_27_io_out ? io_r_50_b : _GEN_5749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5751 = 8'h33 == r_count_27_io_out ? io_r_51_b : _GEN_5750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5752 = 8'h34 == r_count_27_io_out ? io_r_52_b : _GEN_5751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5753 = 8'h35 == r_count_27_io_out ? io_r_53_b : _GEN_5752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5754 = 8'h36 == r_count_27_io_out ? io_r_54_b : _GEN_5753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5755 = 8'h37 == r_count_27_io_out ? io_r_55_b : _GEN_5754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5756 = 8'h38 == r_count_27_io_out ? io_r_56_b : _GEN_5755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5757 = 8'h39 == r_count_27_io_out ? io_r_57_b : _GEN_5756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5758 = 8'h3a == r_count_27_io_out ? io_r_58_b : _GEN_5757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5759 = 8'h3b == r_count_27_io_out ? io_r_59_b : _GEN_5758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5760 = 8'h3c == r_count_27_io_out ? io_r_60_b : _GEN_5759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5761 = 8'h3d == r_count_27_io_out ? io_r_61_b : _GEN_5760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5762 = 8'h3e == r_count_27_io_out ? io_r_62_b : _GEN_5761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5763 = 8'h3f == r_count_27_io_out ? io_r_63_b : _GEN_5762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5764 = 8'h40 == r_count_27_io_out ? io_r_64_b : _GEN_5763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5765 = 8'h41 == r_count_27_io_out ? io_r_65_b : _GEN_5764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5766 = 8'h42 == r_count_27_io_out ? io_r_66_b : _GEN_5765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5767 = 8'h43 == r_count_27_io_out ? io_r_67_b : _GEN_5766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5768 = 8'h44 == r_count_27_io_out ? io_r_68_b : _GEN_5767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5769 = 8'h45 == r_count_27_io_out ? io_r_69_b : _GEN_5768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5770 = 8'h46 == r_count_27_io_out ? io_r_70_b : _GEN_5769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5771 = 8'h47 == r_count_27_io_out ? io_r_71_b : _GEN_5770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5772 = 8'h48 == r_count_27_io_out ? io_r_72_b : _GEN_5771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5773 = 8'h49 == r_count_27_io_out ? io_r_73_b : _GEN_5772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5774 = 8'h4a == r_count_27_io_out ? io_r_74_b : _GEN_5773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5775 = 8'h4b == r_count_27_io_out ? io_r_75_b : _GEN_5774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5776 = 8'h4c == r_count_27_io_out ? io_r_76_b : _GEN_5775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5777 = 8'h4d == r_count_27_io_out ? io_r_77_b : _GEN_5776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5778 = 8'h4e == r_count_27_io_out ? io_r_78_b : _GEN_5777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5779 = 8'h4f == r_count_27_io_out ? io_r_79_b : _GEN_5778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5780 = 8'h50 == r_count_27_io_out ? io_r_80_b : _GEN_5779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5781 = 8'h51 == r_count_27_io_out ? io_r_81_b : _GEN_5780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5782 = 8'h52 == r_count_27_io_out ? io_r_82_b : _GEN_5781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5783 = 8'h53 == r_count_27_io_out ? io_r_83_b : _GEN_5782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5784 = 8'h54 == r_count_27_io_out ? io_r_84_b : _GEN_5783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5785 = 8'h55 == r_count_27_io_out ? io_r_85_b : _GEN_5784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5786 = 8'h56 == r_count_27_io_out ? io_r_86_b : _GEN_5785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5787 = 8'h57 == r_count_27_io_out ? io_r_87_b : _GEN_5786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5788 = 8'h58 == r_count_27_io_out ? io_r_88_b : _GEN_5787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5789 = 8'h59 == r_count_27_io_out ? io_r_89_b : _GEN_5788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5790 = 8'h5a == r_count_27_io_out ? io_r_90_b : _GEN_5789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5791 = 8'h5b == r_count_27_io_out ? io_r_91_b : _GEN_5790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5792 = 8'h5c == r_count_27_io_out ? io_r_92_b : _GEN_5791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5793 = 8'h5d == r_count_27_io_out ? io_r_93_b : _GEN_5792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5794 = 8'h5e == r_count_27_io_out ? io_r_94_b : _GEN_5793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5795 = 8'h5f == r_count_27_io_out ? io_r_95_b : _GEN_5794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5796 = 8'h60 == r_count_27_io_out ? io_r_96_b : _GEN_5795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5797 = 8'h61 == r_count_27_io_out ? io_r_97_b : _GEN_5796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5798 = 8'h62 == r_count_27_io_out ? io_r_98_b : _GEN_5797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5799 = 8'h63 == r_count_27_io_out ? io_r_99_b : _GEN_5798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5800 = 8'h64 == r_count_27_io_out ? io_r_100_b : _GEN_5799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5801 = 8'h65 == r_count_27_io_out ? io_r_101_b : _GEN_5800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5802 = 8'h66 == r_count_27_io_out ? io_r_102_b : _GEN_5801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5803 = 8'h67 == r_count_27_io_out ? io_r_103_b : _GEN_5802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5804 = 8'h68 == r_count_27_io_out ? io_r_104_b : _GEN_5803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5805 = 8'h69 == r_count_27_io_out ? io_r_105_b : _GEN_5804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5806 = 8'h6a == r_count_27_io_out ? io_r_106_b : _GEN_5805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5807 = 8'h6b == r_count_27_io_out ? io_r_107_b : _GEN_5806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5808 = 8'h6c == r_count_27_io_out ? io_r_108_b : _GEN_5807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5809 = 8'h6d == r_count_27_io_out ? io_r_109_b : _GEN_5808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5810 = 8'h6e == r_count_27_io_out ? io_r_110_b : _GEN_5809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5811 = 8'h6f == r_count_27_io_out ? io_r_111_b : _GEN_5810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5812 = 8'h70 == r_count_27_io_out ? io_r_112_b : _GEN_5811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5813 = 8'h71 == r_count_27_io_out ? io_r_113_b : _GEN_5812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5814 = 8'h72 == r_count_27_io_out ? io_r_114_b : _GEN_5813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5815 = 8'h73 == r_count_27_io_out ? io_r_115_b : _GEN_5814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5816 = 8'h74 == r_count_27_io_out ? io_r_116_b : _GEN_5815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5817 = 8'h75 == r_count_27_io_out ? io_r_117_b : _GEN_5816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5818 = 8'h76 == r_count_27_io_out ? io_r_118_b : _GEN_5817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5819 = 8'h77 == r_count_27_io_out ? io_r_119_b : _GEN_5818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5820 = 8'h78 == r_count_27_io_out ? io_r_120_b : _GEN_5819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5821 = 8'h79 == r_count_27_io_out ? io_r_121_b : _GEN_5820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5822 = 8'h7a == r_count_27_io_out ? io_r_122_b : _GEN_5821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5823 = 8'h7b == r_count_27_io_out ? io_r_123_b : _GEN_5822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5824 = 8'h7c == r_count_27_io_out ? io_r_124_b : _GEN_5823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5825 = 8'h7d == r_count_27_io_out ? io_r_125_b : _GEN_5824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5826 = 8'h7e == r_count_27_io_out ? io_r_126_b : _GEN_5825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5827 = 8'h7f == r_count_27_io_out ? io_r_127_b : _GEN_5826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5828 = 8'h80 == r_count_27_io_out ? io_r_128_b : _GEN_5827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5829 = 8'h81 == r_count_27_io_out ? io_r_129_b : _GEN_5828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5830 = 8'h82 == r_count_27_io_out ? io_r_130_b : _GEN_5829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5831 = 8'h83 == r_count_27_io_out ? io_r_131_b : _GEN_5830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5832 = 8'h84 == r_count_27_io_out ? io_r_132_b : _GEN_5831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5833 = 8'h85 == r_count_27_io_out ? io_r_133_b : _GEN_5832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5834 = 8'h86 == r_count_27_io_out ? io_r_134_b : _GEN_5833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5835 = 8'h87 == r_count_27_io_out ? io_r_135_b : _GEN_5834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5836 = 8'h88 == r_count_27_io_out ? io_r_136_b : _GEN_5835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5837 = 8'h89 == r_count_27_io_out ? io_r_137_b : _GEN_5836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5838 = 8'h8a == r_count_27_io_out ? io_r_138_b : _GEN_5837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5839 = 8'h8b == r_count_27_io_out ? io_r_139_b : _GEN_5838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5840 = 8'h8c == r_count_27_io_out ? io_r_140_b : _GEN_5839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5841 = 8'h8d == r_count_27_io_out ? io_r_141_b : _GEN_5840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5842 = 8'h8e == r_count_27_io_out ? io_r_142_b : _GEN_5841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5843 = 8'h8f == r_count_27_io_out ? io_r_143_b : _GEN_5842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5844 = 8'h90 == r_count_27_io_out ? io_r_144_b : _GEN_5843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5845 = 8'h91 == r_count_27_io_out ? io_r_145_b : _GEN_5844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5846 = 8'h92 == r_count_27_io_out ? io_r_146_b : _GEN_5845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5847 = 8'h93 == r_count_27_io_out ? io_r_147_b : _GEN_5846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5848 = 8'h94 == r_count_27_io_out ? io_r_148_b : _GEN_5847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5849 = 8'h95 == r_count_27_io_out ? io_r_149_b : _GEN_5848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5850 = 8'h96 == r_count_27_io_out ? io_r_150_b : _GEN_5849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5851 = 8'h97 == r_count_27_io_out ? io_r_151_b : _GEN_5850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5852 = 8'h98 == r_count_27_io_out ? io_r_152_b : _GEN_5851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5853 = 8'h99 == r_count_27_io_out ? io_r_153_b : _GEN_5852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5854 = 8'h9a == r_count_27_io_out ? io_r_154_b : _GEN_5853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5855 = 8'h9b == r_count_27_io_out ? io_r_155_b : _GEN_5854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5856 = 8'h9c == r_count_27_io_out ? io_r_156_b : _GEN_5855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5857 = 8'h9d == r_count_27_io_out ? io_r_157_b : _GEN_5856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5858 = 8'h9e == r_count_27_io_out ? io_r_158_b : _GEN_5857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5859 = 8'h9f == r_count_27_io_out ? io_r_159_b : _GEN_5858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5860 = 8'ha0 == r_count_27_io_out ? io_r_160_b : _GEN_5859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5861 = 8'ha1 == r_count_27_io_out ? io_r_161_b : _GEN_5860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5862 = 8'ha2 == r_count_27_io_out ? io_r_162_b : _GEN_5861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5863 = 8'ha3 == r_count_27_io_out ? io_r_163_b : _GEN_5862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5864 = 8'ha4 == r_count_27_io_out ? io_r_164_b : _GEN_5863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5865 = 8'ha5 == r_count_27_io_out ? io_r_165_b : _GEN_5864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5866 = 8'ha6 == r_count_27_io_out ? io_r_166_b : _GEN_5865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5867 = 8'ha7 == r_count_27_io_out ? io_r_167_b : _GEN_5866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5868 = 8'ha8 == r_count_27_io_out ? io_r_168_b : _GEN_5867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5869 = 8'ha9 == r_count_27_io_out ? io_r_169_b : _GEN_5868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5870 = 8'haa == r_count_27_io_out ? io_r_170_b : _GEN_5869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5871 = 8'hab == r_count_27_io_out ? io_r_171_b : _GEN_5870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5872 = 8'hac == r_count_27_io_out ? io_r_172_b : _GEN_5871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5873 = 8'had == r_count_27_io_out ? io_r_173_b : _GEN_5872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5874 = 8'hae == r_count_27_io_out ? io_r_174_b : _GEN_5873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5875 = 8'haf == r_count_27_io_out ? io_r_175_b : _GEN_5874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5876 = 8'hb0 == r_count_27_io_out ? io_r_176_b : _GEN_5875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5877 = 8'hb1 == r_count_27_io_out ? io_r_177_b : _GEN_5876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5878 = 8'hb2 == r_count_27_io_out ? io_r_178_b : _GEN_5877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5879 = 8'hb3 == r_count_27_io_out ? io_r_179_b : _GEN_5878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5880 = 8'hb4 == r_count_27_io_out ? io_r_180_b : _GEN_5879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5881 = 8'hb5 == r_count_27_io_out ? io_r_181_b : _GEN_5880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5882 = 8'hb6 == r_count_27_io_out ? io_r_182_b : _GEN_5881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5883 = 8'hb7 == r_count_27_io_out ? io_r_183_b : _GEN_5882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5884 = 8'hb8 == r_count_27_io_out ? io_r_184_b : _GEN_5883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5885 = 8'hb9 == r_count_27_io_out ? io_r_185_b : _GEN_5884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5886 = 8'hba == r_count_27_io_out ? io_r_186_b : _GEN_5885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5887 = 8'hbb == r_count_27_io_out ? io_r_187_b : _GEN_5886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5888 = 8'hbc == r_count_27_io_out ? io_r_188_b : _GEN_5887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5889 = 8'hbd == r_count_27_io_out ? io_r_189_b : _GEN_5888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5890 = 8'hbe == r_count_27_io_out ? io_r_190_b : _GEN_5889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5891 = 8'hbf == r_count_27_io_out ? io_r_191_b : _GEN_5890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5892 = 8'hc0 == r_count_27_io_out ? io_r_192_b : _GEN_5891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5893 = 8'hc1 == r_count_27_io_out ? io_r_193_b : _GEN_5892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5894 = 8'hc2 == r_count_27_io_out ? io_r_194_b : _GEN_5893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5895 = 8'hc3 == r_count_27_io_out ? io_r_195_b : _GEN_5894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5896 = 8'hc4 == r_count_27_io_out ? io_r_196_b : _GEN_5895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5897 = 8'hc5 == r_count_27_io_out ? io_r_197_b : _GEN_5896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5898 = 8'hc6 == r_count_27_io_out ? io_r_198_b : _GEN_5897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5901 = 8'h1 == r_count_28_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5902 = 8'h2 == r_count_28_io_out ? io_r_2_b : _GEN_5901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5903 = 8'h3 == r_count_28_io_out ? io_r_3_b : _GEN_5902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5904 = 8'h4 == r_count_28_io_out ? io_r_4_b : _GEN_5903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5905 = 8'h5 == r_count_28_io_out ? io_r_5_b : _GEN_5904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5906 = 8'h6 == r_count_28_io_out ? io_r_6_b : _GEN_5905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5907 = 8'h7 == r_count_28_io_out ? io_r_7_b : _GEN_5906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5908 = 8'h8 == r_count_28_io_out ? io_r_8_b : _GEN_5907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5909 = 8'h9 == r_count_28_io_out ? io_r_9_b : _GEN_5908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5910 = 8'ha == r_count_28_io_out ? io_r_10_b : _GEN_5909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5911 = 8'hb == r_count_28_io_out ? io_r_11_b : _GEN_5910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5912 = 8'hc == r_count_28_io_out ? io_r_12_b : _GEN_5911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5913 = 8'hd == r_count_28_io_out ? io_r_13_b : _GEN_5912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5914 = 8'he == r_count_28_io_out ? io_r_14_b : _GEN_5913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5915 = 8'hf == r_count_28_io_out ? io_r_15_b : _GEN_5914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5916 = 8'h10 == r_count_28_io_out ? io_r_16_b : _GEN_5915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5917 = 8'h11 == r_count_28_io_out ? io_r_17_b : _GEN_5916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5918 = 8'h12 == r_count_28_io_out ? io_r_18_b : _GEN_5917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5919 = 8'h13 == r_count_28_io_out ? io_r_19_b : _GEN_5918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5920 = 8'h14 == r_count_28_io_out ? io_r_20_b : _GEN_5919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5921 = 8'h15 == r_count_28_io_out ? io_r_21_b : _GEN_5920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5922 = 8'h16 == r_count_28_io_out ? io_r_22_b : _GEN_5921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5923 = 8'h17 == r_count_28_io_out ? io_r_23_b : _GEN_5922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5924 = 8'h18 == r_count_28_io_out ? io_r_24_b : _GEN_5923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5925 = 8'h19 == r_count_28_io_out ? io_r_25_b : _GEN_5924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5926 = 8'h1a == r_count_28_io_out ? io_r_26_b : _GEN_5925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5927 = 8'h1b == r_count_28_io_out ? io_r_27_b : _GEN_5926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5928 = 8'h1c == r_count_28_io_out ? io_r_28_b : _GEN_5927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5929 = 8'h1d == r_count_28_io_out ? io_r_29_b : _GEN_5928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5930 = 8'h1e == r_count_28_io_out ? io_r_30_b : _GEN_5929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5931 = 8'h1f == r_count_28_io_out ? io_r_31_b : _GEN_5930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5932 = 8'h20 == r_count_28_io_out ? io_r_32_b : _GEN_5931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5933 = 8'h21 == r_count_28_io_out ? io_r_33_b : _GEN_5932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5934 = 8'h22 == r_count_28_io_out ? io_r_34_b : _GEN_5933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5935 = 8'h23 == r_count_28_io_out ? io_r_35_b : _GEN_5934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5936 = 8'h24 == r_count_28_io_out ? io_r_36_b : _GEN_5935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5937 = 8'h25 == r_count_28_io_out ? io_r_37_b : _GEN_5936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5938 = 8'h26 == r_count_28_io_out ? io_r_38_b : _GEN_5937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5939 = 8'h27 == r_count_28_io_out ? io_r_39_b : _GEN_5938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5940 = 8'h28 == r_count_28_io_out ? io_r_40_b : _GEN_5939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5941 = 8'h29 == r_count_28_io_out ? io_r_41_b : _GEN_5940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5942 = 8'h2a == r_count_28_io_out ? io_r_42_b : _GEN_5941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5943 = 8'h2b == r_count_28_io_out ? io_r_43_b : _GEN_5942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5944 = 8'h2c == r_count_28_io_out ? io_r_44_b : _GEN_5943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5945 = 8'h2d == r_count_28_io_out ? io_r_45_b : _GEN_5944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5946 = 8'h2e == r_count_28_io_out ? io_r_46_b : _GEN_5945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5947 = 8'h2f == r_count_28_io_out ? io_r_47_b : _GEN_5946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5948 = 8'h30 == r_count_28_io_out ? io_r_48_b : _GEN_5947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5949 = 8'h31 == r_count_28_io_out ? io_r_49_b : _GEN_5948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5950 = 8'h32 == r_count_28_io_out ? io_r_50_b : _GEN_5949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5951 = 8'h33 == r_count_28_io_out ? io_r_51_b : _GEN_5950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5952 = 8'h34 == r_count_28_io_out ? io_r_52_b : _GEN_5951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5953 = 8'h35 == r_count_28_io_out ? io_r_53_b : _GEN_5952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5954 = 8'h36 == r_count_28_io_out ? io_r_54_b : _GEN_5953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5955 = 8'h37 == r_count_28_io_out ? io_r_55_b : _GEN_5954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5956 = 8'h38 == r_count_28_io_out ? io_r_56_b : _GEN_5955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5957 = 8'h39 == r_count_28_io_out ? io_r_57_b : _GEN_5956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5958 = 8'h3a == r_count_28_io_out ? io_r_58_b : _GEN_5957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5959 = 8'h3b == r_count_28_io_out ? io_r_59_b : _GEN_5958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5960 = 8'h3c == r_count_28_io_out ? io_r_60_b : _GEN_5959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5961 = 8'h3d == r_count_28_io_out ? io_r_61_b : _GEN_5960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5962 = 8'h3e == r_count_28_io_out ? io_r_62_b : _GEN_5961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5963 = 8'h3f == r_count_28_io_out ? io_r_63_b : _GEN_5962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5964 = 8'h40 == r_count_28_io_out ? io_r_64_b : _GEN_5963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5965 = 8'h41 == r_count_28_io_out ? io_r_65_b : _GEN_5964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5966 = 8'h42 == r_count_28_io_out ? io_r_66_b : _GEN_5965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5967 = 8'h43 == r_count_28_io_out ? io_r_67_b : _GEN_5966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5968 = 8'h44 == r_count_28_io_out ? io_r_68_b : _GEN_5967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5969 = 8'h45 == r_count_28_io_out ? io_r_69_b : _GEN_5968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5970 = 8'h46 == r_count_28_io_out ? io_r_70_b : _GEN_5969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5971 = 8'h47 == r_count_28_io_out ? io_r_71_b : _GEN_5970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5972 = 8'h48 == r_count_28_io_out ? io_r_72_b : _GEN_5971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5973 = 8'h49 == r_count_28_io_out ? io_r_73_b : _GEN_5972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5974 = 8'h4a == r_count_28_io_out ? io_r_74_b : _GEN_5973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5975 = 8'h4b == r_count_28_io_out ? io_r_75_b : _GEN_5974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5976 = 8'h4c == r_count_28_io_out ? io_r_76_b : _GEN_5975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5977 = 8'h4d == r_count_28_io_out ? io_r_77_b : _GEN_5976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5978 = 8'h4e == r_count_28_io_out ? io_r_78_b : _GEN_5977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5979 = 8'h4f == r_count_28_io_out ? io_r_79_b : _GEN_5978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5980 = 8'h50 == r_count_28_io_out ? io_r_80_b : _GEN_5979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5981 = 8'h51 == r_count_28_io_out ? io_r_81_b : _GEN_5980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5982 = 8'h52 == r_count_28_io_out ? io_r_82_b : _GEN_5981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5983 = 8'h53 == r_count_28_io_out ? io_r_83_b : _GEN_5982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5984 = 8'h54 == r_count_28_io_out ? io_r_84_b : _GEN_5983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5985 = 8'h55 == r_count_28_io_out ? io_r_85_b : _GEN_5984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5986 = 8'h56 == r_count_28_io_out ? io_r_86_b : _GEN_5985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5987 = 8'h57 == r_count_28_io_out ? io_r_87_b : _GEN_5986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5988 = 8'h58 == r_count_28_io_out ? io_r_88_b : _GEN_5987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5989 = 8'h59 == r_count_28_io_out ? io_r_89_b : _GEN_5988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5990 = 8'h5a == r_count_28_io_out ? io_r_90_b : _GEN_5989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5991 = 8'h5b == r_count_28_io_out ? io_r_91_b : _GEN_5990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5992 = 8'h5c == r_count_28_io_out ? io_r_92_b : _GEN_5991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5993 = 8'h5d == r_count_28_io_out ? io_r_93_b : _GEN_5992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5994 = 8'h5e == r_count_28_io_out ? io_r_94_b : _GEN_5993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5995 = 8'h5f == r_count_28_io_out ? io_r_95_b : _GEN_5994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5996 = 8'h60 == r_count_28_io_out ? io_r_96_b : _GEN_5995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5997 = 8'h61 == r_count_28_io_out ? io_r_97_b : _GEN_5996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5998 = 8'h62 == r_count_28_io_out ? io_r_98_b : _GEN_5997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5999 = 8'h63 == r_count_28_io_out ? io_r_99_b : _GEN_5998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6000 = 8'h64 == r_count_28_io_out ? io_r_100_b : _GEN_5999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6001 = 8'h65 == r_count_28_io_out ? io_r_101_b : _GEN_6000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6002 = 8'h66 == r_count_28_io_out ? io_r_102_b : _GEN_6001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6003 = 8'h67 == r_count_28_io_out ? io_r_103_b : _GEN_6002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6004 = 8'h68 == r_count_28_io_out ? io_r_104_b : _GEN_6003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6005 = 8'h69 == r_count_28_io_out ? io_r_105_b : _GEN_6004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6006 = 8'h6a == r_count_28_io_out ? io_r_106_b : _GEN_6005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6007 = 8'h6b == r_count_28_io_out ? io_r_107_b : _GEN_6006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6008 = 8'h6c == r_count_28_io_out ? io_r_108_b : _GEN_6007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6009 = 8'h6d == r_count_28_io_out ? io_r_109_b : _GEN_6008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6010 = 8'h6e == r_count_28_io_out ? io_r_110_b : _GEN_6009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6011 = 8'h6f == r_count_28_io_out ? io_r_111_b : _GEN_6010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6012 = 8'h70 == r_count_28_io_out ? io_r_112_b : _GEN_6011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6013 = 8'h71 == r_count_28_io_out ? io_r_113_b : _GEN_6012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6014 = 8'h72 == r_count_28_io_out ? io_r_114_b : _GEN_6013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6015 = 8'h73 == r_count_28_io_out ? io_r_115_b : _GEN_6014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6016 = 8'h74 == r_count_28_io_out ? io_r_116_b : _GEN_6015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6017 = 8'h75 == r_count_28_io_out ? io_r_117_b : _GEN_6016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6018 = 8'h76 == r_count_28_io_out ? io_r_118_b : _GEN_6017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6019 = 8'h77 == r_count_28_io_out ? io_r_119_b : _GEN_6018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6020 = 8'h78 == r_count_28_io_out ? io_r_120_b : _GEN_6019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6021 = 8'h79 == r_count_28_io_out ? io_r_121_b : _GEN_6020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6022 = 8'h7a == r_count_28_io_out ? io_r_122_b : _GEN_6021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6023 = 8'h7b == r_count_28_io_out ? io_r_123_b : _GEN_6022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6024 = 8'h7c == r_count_28_io_out ? io_r_124_b : _GEN_6023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6025 = 8'h7d == r_count_28_io_out ? io_r_125_b : _GEN_6024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6026 = 8'h7e == r_count_28_io_out ? io_r_126_b : _GEN_6025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6027 = 8'h7f == r_count_28_io_out ? io_r_127_b : _GEN_6026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6028 = 8'h80 == r_count_28_io_out ? io_r_128_b : _GEN_6027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6029 = 8'h81 == r_count_28_io_out ? io_r_129_b : _GEN_6028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6030 = 8'h82 == r_count_28_io_out ? io_r_130_b : _GEN_6029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6031 = 8'h83 == r_count_28_io_out ? io_r_131_b : _GEN_6030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6032 = 8'h84 == r_count_28_io_out ? io_r_132_b : _GEN_6031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6033 = 8'h85 == r_count_28_io_out ? io_r_133_b : _GEN_6032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6034 = 8'h86 == r_count_28_io_out ? io_r_134_b : _GEN_6033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6035 = 8'h87 == r_count_28_io_out ? io_r_135_b : _GEN_6034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6036 = 8'h88 == r_count_28_io_out ? io_r_136_b : _GEN_6035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6037 = 8'h89 == r_count_28_io_out ? io_r_137_b : _GEN_6036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6038 = 8'h8a == r_count_28_io_out ? io_r_138_b : _GEN_6037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6039 = 8'h8b == r_count_28_io_out ? io_r_139_b : _GEN_6038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6040 = 8'h8c == r_count_28_io_out ? io_r_140_b : _GEN_6039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6041 = 8'h8d == r_count_28_io_out ? io_r_141_b : _GEN_6040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6042 = 8'h8e == r_count_28_io_out ? io_r_142_b : _GEN_6041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6043 = 8'h8f == r_count_28_io_out ? io_r_143_b : _GEN_6042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6044 = 8'h90 == r_count_28_io_out ? io_r_144_b : _GEN_6043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6045 = 8'h91 == r_count_28_io_out ? io_r_145_b : _GEN_6044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6046 = 8'h92 == r_count_28_io_out ? io_r_146_b : _GEN_6045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6047 = 8'h93 == r_count_28_io_out ? io_r_147_b : _GEN_6046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6048 = 8'h94 == r_count_28_io_out ? io_r_148_b : _GEN_6047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6049 = 8'h95 == r_count_28_io_out ? io_r_149_b : _GEN_6048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6050 = 8'h96 == r_count_28_io_out ? io_r_150_b : _GEN_6049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6051 = 8'h97 == r_count_28_io_out ? io_r_151_b : _GEN_6050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6052 = 8'h98 == r_count_28_io_out ? io_r_152_b : _GEN_6051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6053 = 8'h99 == r_count_28_io_out ? io_r_153_b : _GEN_6052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6054 = 8'h9a == r_count_28_io_out ? io_r_154_b : _GEN_6053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6055 = 8'h9b == r_count_28_io_out ? io_r_155_b : _GEN_6054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6056 = 8'h9c == r_count_28_io_out ? io_r_156_b : _GEN_6055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6057 = 8'h9d == r_count_28_io_out ? io_r_157_b : _GEN_6056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6058 = 8'h9e == r_count_28_io_out ? io_r_158_b : _GEN_6057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6059 = 8'h9f == r_count_28_io_out ? io_r_159_b : _GEN_6058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6060 = 8'ha0 == r_count_28_io_out ? io_r_160_b : _GEN_6059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6061 = 8'ha1 == r_count_28_io_out ? io_r_161_b : _GEN_6060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6062 = 8'ha2 == r_count_28_io_out ? io_r_162_b : _GEN_6061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6063 = 8'ha3 == r_count_28_io_out ? io_r_163_b : _GEN_6062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6064 = 8'ha4 == r_count_28_io_out ? io_r_164_b : _GEN_6063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6065 = 8'ha5 == r_count_28_io_out ? io_r_165_b : _GEN_6064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6066 = 8'ha6 == r_count_28_io_out ? io_r_166_b : _GEN_6065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6067 = 8'ha7 == r_count_28_io_out ? io_r_167_b : _GEN_6066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6068 = 8'ha8 == r_count_28_io_out ? io_r_168_b : _GEN_6067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6069 = 8'ha9 == r_count_28_io_out ? io_r_169_b : _GEN_6068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6070 = 8'haa == r_count_28_io_out ? io_r_170_b : _GEN_6069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6071 = 8'hab == r_count_28_io_out ? io_r_171_b : _GEN_6070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6072 = 8'hac == r_count_28_io_out ? io_r_172_b : _GEN_6071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6073 = 8'had == r_count_28_io_out ? io_r_173_b : _GEN_6072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6074 = 8'hae == r_count_28_io_out ? io_r_174_b : _GEN_6073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6075 = 8'haf == r_count_28_io_out ? io_r_175_b : _GEN_6074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6076 = 8'hb0 == r_count_28_io_out ? io_r_176_b : _GEN_6075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6077 = 8'hb1 == r_count_28_io_out ? io_r_177_b : _GEN_6076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6078 = 8'hb2 == r_count_28_io_out ? io_r_178_b : _GEN_6077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6079 = 8'hb3 == r_count_28_io_out ? io_r_179_b : _GEN_6078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6080 = 8'hb4 == r_count_28_io_out ? io_r_180_b : _GEN_6079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6081 = 8'hb5 == r_count_28_io_out ? io_r_181_b : _GEN_6080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6082 = 8'hb6 == r_count_28_io_out ? io_r_182_b : _GEN_6081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6083 = 8'hb7 == r_count_28_io_out ? io_r_183_b : _GEN_6082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6084 = 8'hb8 == r_count_28_io_out ? io_r_184_b : _GEN_6083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6085 = 8'hb9 == r_count_28_io_out ? io_r_185_b : _GEN_6084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6086 = 8'hba == r_count_28_io_out ? io_r_186_b : _GEN_6085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6087 = 8'hbb == r_count_28_io_out ? io_r_187_b : _GEN_6086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6088 = 8'hbc == r_count_28_io_out ? io_r_188_b : _GEN_6087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6089 = 8'hbd == r_count_28_io_out ? io_r_189_b : _GEN_6088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6090 = 8'hbe == r_count_28_io_out ? io_r_190_b : _GEN_6089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6091 = 8'hbf == r_count_28_io_out ? io_r_191_b : _GEN_6090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6092 = 8'hc0 == r_count_28_io_out ? io_r_192_b : _GEN_6091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6093 = 8'hc1 == r_count_28_io_out ? io_r_193_b : _GEN_6092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6094 = 8'hc2 == r_count_28_io_out ? io_r_194_b : _GEN_6093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6095 = 8'hc3 == r_count_28_io_out ? io_r_195_b : _GEN_6094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6096 = 8'hc4 == r_count_28_io_out ? io_r_196_b : _GEN_6095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6097 = 8'hc5 == r_count_28_io_out ? io_r_197_b : _GEN_6096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6098 = 8'hc6 == r_count_28_io_out ? io_r_198_b : _GEN_6097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6101 = 8'h1 == r_count_29_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6102 = 8'h2 == r_count_29_io_out ? io_r_2_b : _GEN_6101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6103 = 8'h3 == r_count_29_io_out ? io_r_3_b : _GEN_6102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6104 = 8'h4 == r_count_29_io_out ? io_r_4_b : _GEN_6103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6105 = 8'h5 == r_count_29_io_out ? io_r_5_b : _GEN_6104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6106 = 8'h6 == r_count_29_io_out ? io_r_6_b : _GEN_6105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6107 = 8'h7 == r_count_29_io_out ? io_r_7_b : _GEN_6106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6108 = 8'h8 == r_count_29_io_out ? io_r_8_b : _GEN_6107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6109 = 8'h9 == r_count_29_io_out ? io_r_9_b : _GEN_6108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6110 = 8'ha == r_count_29_io_out ? io_r_10_b : _GEN_6109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6111 = 8'hb == r_count_29_io_out ? io_r_11_b : _GEN_6110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6112 = 8'hc == r_count_29_io_out ? io_r_12_b : _GEN_6111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6113 = 8'hd == r_count_29_io_out ? io_r_13_b : _GEN_6112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6114 = 8'he == r_count_29_io_out ? io_r_14_b : _GEN_6113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6115 = 8'hf == r_count_29_io_out ? io_r_15_b : _GEN_6114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6116 = 8'h10 == r_count_29_io_out ? io_r_16_b : _GEN_6115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6117 = 8'h11 == r_count_29_io_out ? io_r_17_b : _GEN_6116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6118 = 8'h12 == r_count_29_io_out ? io_r_18_b : _GEN_6117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6119 = 8'h13 == r_count_29_io_out ? io_r_19_b : _GEN_6118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6120 = 8'h14 == r_count_29_io_out ? io_r_20_b : _GEN_6119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6121 = 8'h15 == r_count_29_io_out ? io_r_21_b : _GEN_6120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6122 = 8'h16 == r_count_29_io_out ? io_r_22_b : _GEN_6121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6123 = 8'h17 == r_count_29_io_out ? io_r_23_b : _GEN_6122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6124 = 8'h18 == r_count_29_io_out ? io_r_24_b : _GEN_6123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6125 = 8'h19 == r_count_29_io_out ? io_r_25_b : _GEN_6124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6126 = 8'h1a == r_count_29_io_out ? io_r_26_b : _GEN_6125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6127 = 8'h1b == r_count_29_io_out ? io_r_27_b : _GEN_6126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6128 = 8'h1c == r_count_29_io_out ? io_r_28_b : _GEN_6127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6129 = 8'h1d == r_count_29_io_out ? io_r_29_b : _GEN_6128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6130 = 8'h1e == r_count_29_io_out ? io_r_30_b : _GEN_6129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6131 = 8'h1f == r_count_29_io_out ? io_r_31_b : _GEN_6130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6132 = 8'h20 == r_count_29_io_out ? io_r_32_b : _GEN_6131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6133 = 8'h21 == r_count_29_io_out ? io_r_33_b : _GEN_6132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6134 = 8'h22 == r_count_29_io_out ? io_r_34_b : _GEN_6133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6135 = 8'h23 == r_count_29_io_out ? io_r_35_b : _GEN_6134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6136 = 8'h24 == r_count_29_io_out ? io_r_36_b : _GEN_6135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6137 = 8'h25 == r_count_29_io_out ? io_r_37_b : _GEN_6136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6138 = 8'h26 == r_count_29_io_out ? io_r_38_b : _GEN_6137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6139 = 8'h27 == r_count_29_io_out ? io_r_39_b : _GEN_6138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6140 = 8'h28 == r_count_29_io_out ? io_r_40_b : _GEN_6139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6141 = 8'h29 == r_count_29_io_out ? io_r_41_b : _GEN_6140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6142 = 8'h2a == r_count_29_io_out ? io_r_42_b : _GEN_6141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6143 = 8'h2b == r_count_29_io_out ? io_r_43_b : _GEN_6142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6144 = 8'h2c == r_count_29_io_out ? io_r_44_b : _GEN_6143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6145 = 8'h2d == r_count_29_io_out ? io_r_45_b : _GEN_6144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6146 = 8'h2e == r_count_29_io_out ? io_r_46_b : _GEN_6145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6147 = 8'h2f == r_count_29_io_out ? io_r_47_b : _GEN_6146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6148 = 8'h30 == r_count_29_io_out ? io_r_48_b : _GEN_6147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6149 = 8'h31 == r_count_29_io_out ? io_r_49_b : _GEN_6148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6150 = 8'h32 == r_count_29_io_out ? io_r_50_b : _GEN_6149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6151 = 8'h33 == r_count_29_io_out ? io_r_51_b : _GEN_6150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6152 = 8'h34 == r_count_29_io_out ? io_r_52_b : _GEN_6151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6153 = 8'h35 == r_count_29_io_out ? io_r_53_b : _GEN_6152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6154 = 8'h36 == r_count_29_io_out ? io_r_54_b : _GEN_6153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6155 = 8'h37 == r_count_29_io_out ? io_r_55_b : _GEN_6154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6156 = 8'h38 == r_count_29_io_out ? io_r_56_b : _GEN_6155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6157 = 8'h39 == r_count_29_io_out ? io_r_57_b : _GEN_6156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6158 = 8'h3a == r_count_29_io_out ? io_r_58_b : _GEN_6157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6159 = 8'h3b == r_count_29_io_out ? io_r_59_b : _GEN_6158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6160 = 8'h3c == r_count_29_io_out ? io_r_60_b : _GEN_6159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6161 = 8'h3d == r_count_29_io_out ? io_r_61_b : _GEN_6160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6162 = 8'h3e == r_count_29_io_out ? io_r_62_b : _GEN_6161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6163 = 8'h3f == r_count_29_io_out ? io_r_63_b : _GEN_6162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6164 = 8'h40 == r_count_29_io_out ? io_r_64_b : _GEN_6163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6165 = 8'h41 == r_count_29_io_out ? io_r_65_b : _GEN_6164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6166 = 8'h42 == r_count_29_io_out ? io_r_66_b : _GEN_6165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6167 = 8'h43 == r_count_29_io_out ? io_r_67_b : _GEN_6166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6168 = 8'h44 == r_count_29_io_out ? io_r_68_b : _GEN_6167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6169 = 8'h45 == r_count_29_io_out ? io_r_69_b : _GEN_6168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6170 = 8'h46 == r_count_29_io_out ? io_r_70_b : _GEN_6169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6171 = 8'h47 == r_count_29_io_out ? io_r_71_b : _GEN_6170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6172 = 8'h48 == r_count_29_io_out ? io_r_72_b : _GEN_6171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6173 = 8'h49 == r_count_29_io_out ? io_r_73_b : _GEN_6172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6174 = 8'h4a == r_count_29_io_out ? io_r_74_b : _GEN_6173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6175 = 8'h4b == r_count_29_io_out ? io_r_75_b : _GEN_6174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6176 = 8'h4c == r_count_29_io_out ? io_r_76_b : _GEN_6175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6177 = 8'h4d == r_count_29_io_out ? io_r_77_b : _GEN_6176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6178 = 8'h4e == r_count_29_io_out ? io_r_78_b : _GEN_6177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6179 = 8'h4f == r_count_29_io_out ? io_r_79_b : _GEN_6178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6180 = 8'h50 == r_count_29_io_out ? io_r_80_b : _GEN_6179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6181 = 8'h51 == r_count_29_io_out ? io_r_81_b : _GEN_6180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6182 = 8'h52 == r_count_29_io_out ? io_r_82_b : _GEN_6181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6183 = 8'h53 == r_count_29_io_out ? io_r_83_b : _GEN_6182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6184 = 8'h54 == r_count_29_io_out ? io_r_84_b : _GEN_6183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6185 = 8'h55 == r_count_29_io_out ? io_r_85_b : _GEN_6184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6186 = 8'h56 == r_count_29_io_out ? io_r_86_b : _GEN_6185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6187 = 8'h57 == r_count_29_io_out ? io_r_87_b : _GEN_6186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6188 = 8'h58 == r_count_29_io_out ? io_r_88_b : _GEN_6187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6189 = 8'h59 == r_count_29_io_out ? io_r_89_b : _GEN_6188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6190 = 8'h5a == r_count_29_io_out ? io_r_90_b : _GEN_6189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6191 = 8'h5b == r_count_29_io_out ? io_r_91_b : _GEN_6190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6192 = 8'h5c == r_count_29_io_out ? io_r_92_b : _GEN_6191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6193 = 8'h5d == r_count_29_io_out ? io_r_93_b : _GEN_6192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6194 = 8'h5e == r_count_29_io_out ? io_r_94_b : _GEN_6193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6195 = 8'h5f == r_count_29_io_out ? io_r_95_b : _GEN_6194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6196 = 8'h60 == r_count_29_io_out ? io_r_96_b : _GEN_6195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6197 = 8'h61 == r_count_29_io_out ? io_r_97_b : _GEN_6196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6198 = 8'h62 == r_count_29_io_out ? io_r_98_b : _GEN_6197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6199 = 8'h63 == r_count_29_io_out ? io_r_99_b : _GEN_6198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6200 = 8'h64 == r_count_29_io_out ? io_r_100_b : _GEN_6199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6201 = 8'h65 == r_count_29_io_out ? io_r_101_b : _GEN_6200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6202 = 8'h66 == r_count_29_io_out ? io_r_102_b : _GEN_6201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6203 = 8'h67 == r_count_29_io_out ? io_r_103_b : _GEN_6202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6204 = 8'h68 == r_count_29_io_out ? io_r_104_b : _GEN_6203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6205 = 8'h69 == r_count_29_io_out ? io_r_105_b : _GEN_6204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6206 = 8'h6a == r_count_29_io_out ? io_r_106_b : _GEN_6205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6207 = 8'h6b == r_count_29_io_out ? io_r_107_b : _GEN_6206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6208 = 8'h6c == r_count_29_io_out ? io_r_108_b : _GEN_6207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6209 = 8'h6d == r_count_29_io_out ? io_r_109_b : _GEN_6208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6210 = 8'h6e == r_count_29_io_out ? io_r_110_b : _GEN_6209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6211 = 8'h6f == r_count_29_io_out ? io_r_111_b : _GEN_6210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6212 = 8'h70 == r_count_29_io_out ? io_r_112_b : _GEN_6211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6213 = 8'h71 == r_count_29_io_out ? io_r_113_b : _GEN_6212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6214 = 8'h72 == r_count_29_io_out ? io_r_114_b : _GEN_6213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6215 = 8'h73 == r_count_29_io_out ? io_r_115_b : _GEN_6214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6216 = 8'h74 == r_count_29_io_out ? io_r_116_b : _GEN_6215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6217 = 8'h75 == r_count_29_io_out ? io_r_117_b : _GEN_6216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6218 = 8'h76 == r_count_29_io_out ? io_r_118_b : _GEN_6217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6219 = 8'h77 == r_count_29_io_out ? io_r_119_b : _GEN_6218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6220 = 8'h78 == r_count_29_io_out ? io_r_120_b : _GEN_6219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6221 = 8'h79 == r_count_29_io_out ? io_r_121_b : _GEN_6220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6222 = 8'h7a == r_count_29_io_out ? io_r_122_b : _GEN_6221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6223 = 8'h7b == r_count_29_io_out ? io_r_123_b : _GEN_6222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6224 = 8'h7c == r_count_29_io_out ? io_r_124_b : _GEN_6223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6225 = 8'h7d == r_count_29_io_out ? io_r_125_b : _GEN_6224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6226 = 8'h7e == r_count_29_io_out ? io_r_126_b : _GEN_6225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6227 = 8'h7f == r_count_29_io_out ? io_r_127_b : _GEN_6226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6228 = 8'h80 == r_count_29_io_out ? io_r_128_b : _GEN_6227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6229 = 8'h81 == r_count_29_io_out ? io_r_129_b : _GEN_6228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6230 = 8'h82 == r_count_29_io_out ? io_r_130_b : _GEN_6229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6231 = 8'h83 == r_count_29_io_out ? io_r_131_b : _GEN_6230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6232 = 8'h84 == r_count_29_io_out ? io_r_132_b : _GEN_6231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6233 = 8'h85 == r_count_29_io_out ? io_r_133_b : _GEN_6232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6234 = 8'h86 == r_count_29_io_out ? io_r_134_b : _GEN_6233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6235 = 8'h87 == r_count_29_io_out ? io_r_135_b : _GEN_6234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6236 = 8'h88 == r_count_29_io_out ? io_r_136_b : _GEN_6235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6237 = 8'h89 == r_count_29_io_out ? io_r_137_b : _GEN_6236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6238 = 8'h8a == r_count_29_io_out ? io_r_138_b : _GEN_6237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6239 = 8'h8b == r_count_29_io_out ? io_r_139_b : _GEN_6238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6240 = 8'h8c == r_count_29_io_out ? io_r_140_b : _GEN_6239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6241 = 8'h8d == r_count_29_io_out ? io_r_141_b : _GEN_6240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6242 = 8'h8e == r_count_29_io_out ? io_r_142_b : _GEN_6241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6243 = 8'h8f == r_count_29_io_out ? io_r_143_b : _GEN_6242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6244 = 8'h90 == r_count_29_io_out ? io_r_144_b : _GEN_6243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6245 = 8'h91 == r_count_29_io_out ? io_r_145_b : _GEN_6244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6246 = 8'h92 == r_count_29_io_out ? io_r_146_b : _GEN_6245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6247 = 8'h93 == r_count_29_io_out ? io_r_147_b : _GEN_6246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6248 = 8'h94 == r_count_29_io_out ? io_r_148_b : _GEN_6247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6249 = 8'h95 == r_count_29_io_out ? io_r_149_b : _GEN_6248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6250 = 8'h96 == r_count_29_io_out ? io_r_150_b : _GEN_6249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6251 = 8'h97 == r_count_29_io_out ? io_r_151_b : _GEN_6250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6252 = 8'h98 == r_count_29_io_out ? io_r_152_b : _GEN_6251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6253 = 8'h99 == r_count_29_io_out ? io_r_153_b : _GEN_6252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6254 = 8'h9a == r_count_29_io_out ? io_r_154_b : _GEN_6253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6255 = 8'h9b == r_count_29_io_out ? io_r_155_b : _GEN_6254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6256 = 8'h9c == r_count_29_io_out ? io_r_156_b : _GEN_6255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6257 = 8'h9d == r_count_29_io_out ? io_r_157_b : _GEN_6256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6258 = 8'h9e == r_count_29_io_out ? io_r_158_b : _GEN_6257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6259 = 8'h9f == r_count_29_io_out ? io_r_159_b : _GEN_6258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6260 = 8'ha0 == r_count_29_io_out ? io_r_160_b : _GEN_6259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6261 = 8'ha1 == r_count_29_io_out ? io_r_161_b : _GEN_6260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6262 = 8'ha2 == r_count_29_io_out ? io_r_162_b : _GEN_6261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6263 = 8'ha3 == r_count_29_io_out ? io_r_163_b : _GEN_6262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6264 = 8'ha4 == r_count_29_io_out ? io_r_164_b : _GEN_6263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6265 = 8'ha5 == r_count_29_io_out ? io_r_165_b : _GEN_6264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6266 = 8'ha6 == r_count_29_io_out ? io_r_166_b : _GEN_6265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6267 = 8'ha7 == r_count_29_io_out ? io_r_167_b : _GEN_6266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6268 = 8'ha8 == r_count_29_io_out ? io_r_168_b : _GEN_6267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6269 = 8'ha9 == r_count_29_io_out ? io_r_169_b : _GEN_6268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6270 = 8'haa == r_count_29_io_out ? io_r_170_b : _GEN_6269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6271 = 8'hab == r_count_29_io_out ? io_r_171_b : _GEN_6270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6272 = 8'hac == r_count_29_io_out ? io_r_172_b : _GEN_6271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6273 = 8'had == r_count_29_io_out ? io_r_173_b : _GEN_6272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6274 = 8'hae == r_count_29_io_out ? io_r_174_b : _GEN_6273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6275 = 8'haf == r_count_29_io_out ? io_r_175_b : _GEN_6274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6276 = 8'hb0 == r_count_29_io_out ? io_r_176_b : _GEN_6275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6277 = 8'hb1 == r_count_29_io_out ? io_r_177_b : _GEN_6276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6278 = 8'hb2 == r_count_29_io_out ? io_r_178_b : _GEN_6277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6279 = 8'hb3 == r_count_29_io_out ? io_r_179_b : _GEN_6278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6280 = 8'hb4 == r_count_29_io_out ? io_r_180_b : _GEN_6279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6281 = 8'hb5 == r_count_29_io_out ? io_r_181_b : _GEN_6280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6282 = 8'hb6 == r_count_29_io_out ? io_r_182_b : _GEN_6281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6283 = 8'hb7 == r_count_29_io_out ? io_r_183_b : _GEN_6282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6284 = 8'hb8 == r_count_29_io_out ? io_r_184_b : _GEN_6283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6285 = 8'hb9 == r_count_29_io_out ? io_r_185_b : _GEN_6284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6286 = 8'hba == r_count_29_io_out ? io_r_186_b : _GEN_6285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6287 = 8'hbb == r_count_29_io_out ? io_r_187_b : _GEN_6286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6288 = 8'hbc == r_count_29_io_out ? io_r_188_b : _GEN_6287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6289 = 8'hbd == r_count_29_io_out ? io_r_189_b : _GEN_6288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6290 = 8'hbe == r_count_29_io_out ? io_r_190_b : _GEN_6289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6291 = 8'hbf == r_count_29_io_out ? io_r_191_b : _GEN_6290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6292 = 8'hc0 == r_count_29_io_out ? io_r_192_b : _GEN_6291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6293 = 8'hc1 == r_count_29_io_out ? io_r_193_b : _GEN_6292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6294 = 8'hc2 == r_count_29_io_out ? io_r_194_b : _GEN_6293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6295 = 8'hc3 == r_count_29_io_out ? io_r_195_b : _GEN_6294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6296 = 8'hc4 == r_count_29_io_out ? io_r_196_b : _GEN_6295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6297 = 8'hc5 == r_count_29_io_out ? io_r_197_b : _GEN_6296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6298 = 8'hc6 == r_count_29_io_out ? io_r_198_b : _GEN_6297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6301 = 8'h1 == r_count_30_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6302 = 8'h2 == r_count_30_io_out ? io_r_2_b : _GEN_6301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6303 = 8'h3 == r_count_30_io_out ? io_r_3_b : _GEN_6302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6304 = 8'h4 == r_count_30_io_out ? io_r_4_b : _GEN_6303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6305 = 8'h5 == r_count_30_io_out ? io_r_5_b : _GEN_6304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6306 = 8'h6 == r_count_30_io_out ? io_r_6_b : _GEN_6305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6307 = 8'h7 == r_count_30_io_out ? io_r_7_b : _GEN_6306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6308 = 8'h8 == r_count_30_io_out ? io_r_8_b : _GEN_6307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6309 = 8'h9 == r_count_30_io_out ? io_r_9_b : _GEN_6308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6310 = 8'ha == r_count_30_io_out ? io_r_10_b : _GEN_6309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6311 = 8'hb == r_count_30_io_out ? io_r_11_b : _GEN_6310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6312 = 8'hc == r_count_30_io_out ? io_r_12_b : _GEN_6311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6313 = 8'hd == r_count_30_io_out ? io_r_13_b : _GEN_6312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6314 = 8'he == r_count_30_io_out ? io_r_14_b : _GEN_6313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6315 = 8'hf == r_count_30_io_out ? io_r_15_b : _GEN_6314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6316 = 8'h10 == r_count_30_io_out ? io_r_16_b : _GEN_6315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6317 = 8'h11 == r_count_30_io_out ? io_r_17_b : _GEN_6316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6318 = 8'h12 == r_count_30_io_out ? io_r_18_b : _GEN_6317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6319 = 8'h13 == r_count_30_io_out ? io_r_19_b : _GEN_6318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6320 = 8'h14 == r_count_30_io_out ? io_r_20_b : _GEN_6319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6321 = 8'h15 == r_count_30_io_out ? io_r_21_b : _GEN_6320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6322 = 8'h16 == r_count_30_io_out ? io_r_22_b : _GEN_6321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6323 = 8'h17 == r_count_30_io_out ? io_r_23_b : _GEN_6322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6324 = 8'h18 == r_count_30_io_out ? io_r_24_b : _GEN_6323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6325 = 8'h19 == r_count_30_io_out ? io_r_25_b : _GEN_6324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6326 = 8'h1a == r_count_30_io_out ? io_r_26_b : _GEN_6325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6327 = 8'h1b == r_count_30_io_out ? io_r_27_b : _GEN_6326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6328 = 8'h1c == r_count_30_io_out ? io_r_28_b : _GEN_6327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6329 = 8'h1d == r_count_30_io_out ? io_r_29_b : _GEN_6328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6330 = 8'h1e == r_count_30_io_out ? io_r_30_b : _GEN_6329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6331 = 8'h1f == r_count_30_io_out ? io_r_31_b : _GEN_6330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6332 = 8'h20 == r_count_30_io_out ? io_r_32_b : _GEN_6331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6333 = 8'h21 == r_count_30_io_out ? io_r_33_b : _GEN_6332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6334 = 8'h22 == r_count_30_io_out ? io_r_34_b : _GEN_6333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6335 = 8'h23 == r_count_30_io_out ? io_r_35_b : _GEN_6334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6336 = 8'h24 == r_count_30_io_out ? io_r_36_b : _GEN_6335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6337 = 8'h25 == r_count_30_io_out ? io_r_37_b : _GEN_6336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6338 = 8'h26 == r_count_30_io_out ? io_r_38_b : _GEN_6337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6339 = 8'h27 == r_count_30_io_out ? io_r_39_b : _GEN_6338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6340 = 8'h28 == r_count_30_io_out ? io_r_40_b : _GEN_6339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6341 = 8'h29 == r_count_30_io_out ? io_r_41_b : _GEN_6340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6342 = 8'h2a == r_count_30_io_out ? io_r_42_b : _GEN_6341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6343 = 8'h2b == r_count_30_io_out ? io_r_43_b : _GEN_6342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6344 = 8'h2c == r_count_30_io_out ? io_r_44_b : _GEN_6343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6345 = 8'h2d == r_count_30_io_out ? io_r_45_b : _GEN_6344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6346 = 8'h2e == r_count_30_io_out ? io_r_46_b : _GEN_6345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6347 = 8'h2f == r_count_30_io_out ? io_r_47_b : _GEN_6346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6348 = 8'h30 == r_count_30_io_out ? io_r_48_b : _GEN_6347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6349 = 8'h31 == r_count_30_io_out ? io_r_49_b : _GEN_6348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6350 = 8'h32 == r_count_30_io_out ? io_r_50_b : _GEN_6349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6351 = 8'h33 == r_count_30_io_out ? io_r_51_b : _GEN_6350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6352 = 8'h34 == r_count_30_io_out ? io_r_52_b : _GEN_6351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6353 = 8'h35 == r_count_30_io_out ? io_r_53_b : _GEN_6352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6354 = 8'h36 == r_count_30_io_out ? io_r_54_b : _GEN_6353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6355 = 8'h37 == r_count_30_io_out ? io_r_55_b : _GEN_6354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6356 = 8'h38 == r_count_30_io_out ? io_r_56_b : _GEN_6355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6357 = 8'h39 == r_count_30_io_out ? io_r_57_b : _GEN_6356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6358 = 8'h3a == r_count_30_io_out ? io_r_58_b : _GEN_6357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6359 = 8'h3b == r_count_30_io_out ? io_r_59_b : _GEN_6358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6360 = 8'h3c == r_count_30_io_out ? io_r_60_b : _GEN_6359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6361 = 8'h3d == r_count_30_io_out ? io_r_61_b : _GEN_6360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6362 = 8'h3e == r_count_30_io_out ? io_r_62_b : _GEN_6361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6363 = 8'h3f == r_count_30_io_out ? io_r_63_b : _GEN_6362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6364 = 8'h40 == r_count_30_io_out ? io_r_64_b : _GEN_6363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6365 = 8'h41 == r_count_30_io_out ? io_r_65_b : _GEN_6364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6366 = 8'h42 == r_count_30_io_out ? io_r_66_b : _GEN_6365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6367 = 8'h43 == r_count_30_io_out ? io_r_67_b : _GEN_6366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6368 = 8'h44 == r_count_30_io_out ? io_r_68_b : _GEN_6367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6369 = 8'h45 == r_count_30_io_out ? io_r_69_b : _GEN_6368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6370 = 8'h46 == r_count_30_io_out ? io_r_70_b : _GEN_6369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6371 = 8'h47 == r_count_30_io_out ? io_r_71_b : _GEN_6370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6372 = 8'h48 == r_count_30_io_out ? io_r_72_b : _GEN_6371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6373 = 8'h49 == r_count_30_io_out ? io_r_73_b : _GEN_6372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6374 = 8'h4a == r_count_30_io_out ? io_r_74_b : _GEN_6373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6375 = 8'h4b == r_count_30_io_out ? io_r_75_b : _GEN_6374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6376 = 8'h4c == r_count_30_io_out ? io_r_76_b : _GEN_6375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6377 = 8'h4d == r_count_30_io_out ? io_r_77_b : _GEN_6376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6378 = 8'h4e == r_count_30_io_out ? io_r_78_b : _GEN_6377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6379 = 8'h4f == r_count_30_io_out ? io_r_79_b : _GEN_6378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6380 = 8'h50 == r_count_30_io_out ? io_r_80_b : _GEN_6379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6381 = 8'h51 == r_count_30_io_out ? io_r_81_b : _GEN_6380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6382 = 8'h52 == r_count_30_io_out ? io_r_82_b : _GEN_6381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6383 = 8'h53 == r_count_30_io_out ? io_r_83_b : _GEN_6382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6384 = 8'h54 == r_count_30_io_out ? io_r_84_b : _GEN_6383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6385 = 8'h55 == r_count_30_io_out ? io_r_85_b : _GEN_6384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6386 = 8'h56 == r_count_30_io_out ? io_r_86_b : _GEN_6385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6387 = 8'h57 == r_count_30_io_out ? io_r_87_b : _GEN_6386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6388 = 8'h58 == r_count_30_io_out ? io_r_88_b : _GEN_6387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6389 = 8'h59 == r_count_30_io_out ? io_r_89_b : _GEN_6388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6390 = 8'h5a == r_count_30_io_out ? io_r_90_b : _GEN_6389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6391 = 8'h5b == r_count_30_io_out ? io_r_91_b : _GEN_6390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6392 = 8'h5c == r_count_30_io_out ? io_r_92_b : _GEN_6391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6393 = 8'h5d == r_count_30_io_out ? io_r_93_b : _GEN_6392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6394 = 8'h5e == r_count_30_io_out ? io_r_94_b : _GEN_6393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6395 = 8'h5f == r_count_30_io_out ? io_r_95_b : _GEN_6394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6396 = 8'h60 == r_count_30_io_out ? io_r_96_b : _GEN_6395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6397 = 8'h61 == r_count_30_io_out ? io_r_97_b : _GEN_6396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6398 = 8'h62 == r_count_30_io_out ? io_r_98_b : _GEN_6397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6399 = 8'h63 == r_count_30_io_out ? io_r_99_b : _GEN_6398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6400 = 8'h64 == r_count_30_io_out ? io_r_100_b : _GEN_6399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6401 = 8'h65 == r_count_30_io_out ? io_r_101_b : _GEN_6400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6402 = 8'h66 == r_count_30_io_out ? io_r_102_b : _GEN_6401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6403 = 8'h67 == r_count_30_io_out ? io_r_103_b : _GEN_6402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6404 = 8'h68 == r_count_30_io_out ? io_r_104_b : _GEN_6403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6405 = 8'h69 == r_count_30_io_out ? io_r_105_b : _GEN_6404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6406 = 8'h6a == r_count_30_io_out ? io_r_106_b : _GEN_6405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6407 = 8'h6b == r_count_30_io_out ? io_r_107_b : _GEN_6406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6408 = 8'h6c == r_count_30_io_out ? io_r_108_b : _GEN_6407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6409 = 8'h6d == r_count_30_io_out ? io_r_109_b : _GEN_6408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6410 = 8'h6e == r_count_30_io_out ? io_r_110_b : _GEN_6409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6411 = 8'h6f == r_count_30_io_out ? io_r_111_b : _GEN_6410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6412 = 8'h70 == r_count_30_io_out ? io_r_112_b : _GEN_6411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6413 = 8'h71 == r_count_30_io_out ? io_r_113_b : _GEN_6412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6414 = 8'h72 == r_count_30_io_out ? io_r_114_b : _GEN_6413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6415 = 8'h73 == r_count_30_io_out ? io_r_115_b : _GEN_6414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6416 = 8'h74 == r_count_30_io_out ? io_r_116_b : _GEN_6415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6417 = 8'h75 == r_count_30_io_out ? io_r_117_b : _GEN_6416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6418 = 8'h76 == r_count_30_io_out ? io_r_118_b : _GEN_6417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6419 = 8'h77 == r_count_30_io_out ? io_r_119_b : _GEN_6418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6420 = 8'h78 == r_count_30_io_out ? io_r_120_b : _GEN_6419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6421 = 8'h79 == r_count_30_io_out ? io_r_121_b : _GEN_6420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6422 = 8'h7a == r_count_30_io_out ? io_r_122_b : _GEN_6421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6423 = 8'h7b == r_count_30_io_out ? io_r_123_b : _GEN_6422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6424 = 8'h7c == r_count_30_io_out ? io_r_124_b : _GEN_6423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6425 = 8'h7d == r_count_30_io_out ? io_r_125_b : _GEN_6424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6426 = 8'h7e == r_count_30_io_out ? io_r_126_b : _GEN_6425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6427 = 8'h7f == r_count_30_io_out ? io_r_127_b : _GEN_6426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6428 = 8'h80 == r_count_30_io_out ? io_r_128_b : _GEN_6427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6429 = 8'h81 == r_count_30_io_out ? io_r_129_b : _GEN_6428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6430 = 8'h82 == r_count_30_io_out ? io_r_130_b : _GEN_6429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6431 = 8'h83 == r_count_30_io_out ? io_r_131_b : _GEN_6430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6432 = 8'h84 == r_count_30_io_out ? io_r_132_b : _GEN_6431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6433 = 8'h85 == r_count_30_io_out ? io_r_133_b : _GEN_6432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6434 = 8'h86 == r_count_30_io_out ? io_r_134_b : _GEN_6433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6435 = 8'h87 == r_count_30_io_out ? io_r_135_b : _GEN_6434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6436 = 8'h88 == r_count_30_io_out ? io_r_136_b : _GEN_6435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6437 = 8'h89 == r_count_30_io_out ? io_r_137_b : _GEN_6436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6438 = 8'h8a == r_count_30_io_out ? io_r_138_b : _GEN_6437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6439 = 8'h8b == r_count_30_io_out ? io_r_139_b : _GEN_6438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6440 = 8'h8c == r_count_30_io_out ? io_r_140_b : _GEN_6439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6441 = 8'h8d == r_count_30_io_out ? io_r_141_b : _GEN_6440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6442 = 8'h8e == r_count_30_io_out ? io_r_142_b : _GEN_6441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6443 = 8'h8f == r_count_30_io_out ? io_r_143_b : _GEN_6442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6444 = 8'h90 == r_count_30_io_out ? io_r_144_b : _GEN_6443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6445 = 8'h91 == r_count_30_io_out ? io_r_145_b : _GEN_6444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6446 = 8'h92 == r_count_30_io_out ? io_r_146_b : _GEN_6445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6447 = 8'h93 == r_count_30_io_out ? io_r_147_b : _GEN_6446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6448 = 8'h94 == r_count_30_io_out ? io_r_148_b : _GEN_6447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6449 = 8'h95 == r_count_30_io_out ? io_r_149_b : _GEN_6448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6450 = 8'h96 == r_count_30_io_out ? io_r_150_b : _GEN_6449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6451 = 8'h97 == r_count_30_io_out ? io_r_151_b : _GEN_6450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6452 = 8'h98 == r_count_30_io_out ? io_r_152_b : _GEN_6451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6453 = 8'h99 == r_count_30_io_out ? io_r_153_b : _GEN_6452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6454 = 8'h9a == r_count_30_io_out ? io_r_154_b : _GEN_6453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6455 = 8'h9b == r_count_30_io_out ? io_r_155_b : _GEN_6454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6456 = 8'h9c == r_count_30_io_out ? io_r_156_b : _GEN_6455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6457 = 8'h9d == r_count_30_io_out ? io_r_157_b : _GEN_6456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6458 = 8'h9e == r_count_30_io_out ? io_r_158_b : _GEN_6457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6459 = 8'h9f == r_count_30_io_out ? io_r_159_b : _GEN_6458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6460 = 8'ha0 == r_count_30_io_out ? io_r_160_b : _GEN_6459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6461 = 8'ha1 == r_count_30_io_out ? io_r_161_b : _GEN_6460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6462 = 8'ha2 == r_count_30_io_out ? io_r_162_b : _GEN_6461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6463 = 8'ha3 == r_count_30_io_out ? io_r_163_b : _GEN_6462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6464 = 8'ha4 == r_count_30_io_out ? io_r_164_b : _GEN_6463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6465 = 8'ha5 == r_count_30_io_out ? io_r_165_b : _GEN_6464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6466 = 8'ha6 == r_count_30_io_out ? io_r_166_b : _GEN_6465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6467 = 8'ha7 == r_count_30_io_out ? io_r_167_b : _GEN_6466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6468 = 8'ha8 == r_count_30_io_out ? io_r_168_b : _GEN_6467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6469 = 8'ha9 == r_count_30_io_out ? io_r_169_b : _GEN_6468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6470 = 8'haa == r_count_30_io_out ? io_r_170_b : _GEN_6469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6471 = 8'hab == r_count_30_io_out ? io_r_171_b : _GEN_6470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6472 = 8'hac == r_count_30_io_out ? io_r_172_b : _GEN_6471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6473 = 8'had == r_count_30_io_out ? io_r_173_b : _GEN_6472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6474 = 8'hae == r_count_30_io_out ? io_r_174_b : _GEN_6473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6475 = 8'haf == r_count_30_io_out ? io_r_175_b : _GEN_6474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6476 = 8'hb0 == r_count_30_io_out ? io_r_176_b : _GEN_6475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6477 = 8'hb1 == r_count_30_io_out ? io_r_177_b : _GEN_6476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6478 = 8'hb2 == r_count_30_io_out ? io_r_178_b : _GEN_6477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6479 = 8'hb3 == r_count_30_io_out ? io_r_179_b : _GEN_6478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6480 = 8'hb4 == r_count_30_io_out ? io_r_180_b : _GEN_6479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6481 = 8'hb5 == r_count_30_io_out ? io_r_181_b : _GEN_6480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6482 = 8'hb6 == r_count_30_io_out ? io_r_182_b : _GEN_6481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6483 = 8'hb7 == r_count_30_io_out ? io_r_183_b : _GEN_6482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6484 = 8'hb8 == r_count_30_io_out ? io_r_184_b : _GEN_6483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6485 = 8'hb9 == r_count_30_io_out ? io_r_185_b : _GEN_6484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6486 = 8'hba == r_count_30_io_out ? io_r_186_b : _GEN_6485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6487 = 8'hbb == r_count_30_io_out ? io_r_187_b : _GEN_6486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6488 = 8'hbc == r_count_30_io_out ? io_r_188_b : _GEN_6487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6489 = 8'hbd == r_count_30_io_out ? io_r_189_b : _GEN_6488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6490 = 8'hbe == r_count_30_io_out ? io_r_190_b : _GEN_6489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6491 = 8'hbf == r_count_30_io_out ? io_r_191_b : _GEN_6490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6492 = 8'hc0 == r_count_30_io_out ? io_r_192_b : _GEN_6491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6493 = 8'hc1 == r_count_30_io_out ? io_r_193_b : _GEN_6492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6494 = 8'hc2 == r_count_30_io_out ? io_r_194_b : _GEN_6493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6495 = 8'hc3 == r_count_30_io_out ? io_r_195_b : _GEN_6494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6496 = 8'hc4 == r_count_30_io_out ? io_r_196_b : _GEN_6495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6497 = 8'hc5 == r_count_30_io_out ? io_r_197_b : _GEN_6496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6498 = 8'hc6 == r_count_30_io_out ? io_r_198_b : _GEN_6497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6501 = 8'h1 == r_count_31_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6502 = 8'h2 == r_count_31_io_out ? io_r_2_b : _GEN_6501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6503 = 8'h3 == r_count_31_io_out ? io_r_3_b : _GEN_6502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6504 = 8'h4 == r_count_31_io_out ? io_r_4_b : _GEN_6503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6505 = 8'h5 == r_count_31_io_out ? io_r_5_b : _GEN_6504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6506 = 8'h6 == r_count_31_io_out ? io_r_6_b : _GEN_6505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6507 = 8'h7 == r_count_31_io_out ? io_r_7_b : _GEN_6506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6508 = 8'h8 == r_count_31_io_out ? io_r_8_b : _GEN_6507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6509 = 8'h9 == r_count_31_io_out ? io_r_9_b : _GEN_6508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6510 = 8'ha == r_count_31_io_out ? io_r_10_b : _GEN_6509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6511 = 8'hb == r_count_31_io_out ? io_r_11_b : _GEN_6510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6512 = 8'hc == r_count_31_io_out ? io_r_12_b : _GEN_6511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6513 = 8'hd == r_count_31_io_out ? io_r_13_b : _GEN_6512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6514 = 8'he == r_count_31_io_out ? io_r_14_b : _GEN_6513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6515 = 8'hf == r_count_31_io_out ? io_r_15_b : _GEN_6514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6516 = 8'h10 == r_count_31_io_out ? io_r_16_b : _GEN_6515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6517 = 8'h11 == r_count_31_io_out ? io_r_17_b : _GEN_6516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6518 = 8'h12 == r_count_31_io_out ? io_r_18_b : _GEN_6517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6519 = 8'h13 == r_count_31_io_out ? io_r_19_b : _GEN_6518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6520 = 8'h14 == r_count_31_io_out ? io_r_20_b : _GEN_6519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6521 = 8'h15 == r_count_31_io_out ? io_r_21_b : _GEN_6520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6522 = 8'h16 == r_count_31_io_out ? io_r_22_b : _GEN_6521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6523 = 8'h17 == r_count_31_io_out ? io_r_23_b : _GEN_6522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6524 = 8'h18 == r_count_31_io_out ? io_r_24_b : _GEN_6523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6525 = 8'h19 == r_count_31_io_out ? io_r_25_b : _GEN_6524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6526 = 8'h1a == r_count_31_io_out ? io_r_26_b : _GEN_6525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6527 = 8'h1b == r_count_31_io_out ? io_r_27_b : _GEN_6526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6528 = 8'h1c == r_count_31_io_out ? io_r_28_b : _GEN_6527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6529 = 8'h1d == r_count_31_io_out ? io_r_29_b : _GEN_6528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6530 = 8'h1e == r_count_31_io_out ? io_r_30_b : _GEN_6529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6531 = 8'h1f == r_count_31_io_out ? io_r_31_b : _GEN_6530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6532 = 8'h20 == r_count_31_io_out ? io_r_32_b : _GEN_6531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6533 = 8'h21 == r_count_31_io_out ? io_r_33_b : _GEN_6532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6534 = 8'h22 == r_count_31_io_out ? io_r_34_b : _GEN_6533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6535 = 8'h23 == r_count_31_io_out ? io_r_35_b : _GEN_6534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6536 = 8'h24 == r_count_31_io_out ? io_r_36_b : _GEN_6535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6537 = 8'h25 == r_count_31_io_out ? io_r_37_b : _GEN_6536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6538 = 8'h26 == r_count_31_io_out ? io_r_38_b : _GEN_6537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6539 = 8'h27 == r_count_31_io_out ? io_r_39_b : _GEN_6538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6540 = 8'h28 == r_count_31_io_out ? io_r_40_b : _GEN_6539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6541 = 8'h29 == r_count_31_io_out ? io_r_41_b : _GEN_6540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6542 = 8'h2a == r_count_31_io_out ? io_r_42_b : _GEN_6541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6543 = 8'h2b == r_count_31_io_out ? io_r_43_b : _GEN_6542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6544 = 8'h2c == r_count_31_io_out ? io_r_44_b : _GEN_6543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6545 = 8'h2d == r_count_31_io_out ? io_r_45_b : _GEN_6544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6546 = 8'h2e == r_count_31_io_out ? io_r_46_b : _GEN_6545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6547 = 8'h2f == r_count_31_io_out ? io_r_47_b : _GEN_6546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6548 = 8'h30 == r_count_31_io_out ? io_r_48_b : _GEN_6547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6549 = 8'h31 == r_count_31_io_out ? io_r_49_b : _GEN_6548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6550 = 8'h32 == r_count_31_io_out ? io_r_50_b : _GEN_6549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6551 = 8'h33 == r_count_31_io_out ? io_r_51_b : _GEN_6550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6552 = 8'h34 == r_count_31_io_out ? io_r_52_b : _GEN_6551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6553 = 8'h35 == r_count_31_io_out ? io_r_53_b : _GEN_6552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6554 = 8'h36 == r_count_31_io_out ? io_r_54_b : _GEN_6553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6555 = 8'h37 == r_count_31_io_out ? io_r_55_b : _GEN_6554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6556 = 8'h38 == r_count_31_io_out ? io_r_56_b : _GEN_6555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6557 = 8'h39 == r_count_31_io_out ? io_r_57_b : _GEN_6556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6558 = 8'h3a == r_count_31_io_out ? io_r_58_b : _GEN_6557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6559 = 8'h3b == r_count_31_io_out ? io_r_59_b : _GEN_6558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6560 = 8'h3c == r_count_31_io_out ? io_r_60_b : _GEN_6559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6561 = 8'h3d == r_count_31_io_out ? io_r_61_b : _GEN_6560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6562 = 8'h3e == r_count_31_io_out ? io_r_62_b : _GEN_6561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6563 = 8'h3f == r_count_31_io_out ? io_r_63_b : _GEN_6562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6564 = 8'h40 == r_count_31_io_out ? io_r_64_b : _GEN_6563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6565 = 8'h41 == r_count_31_io_out ? io_r_65_b : _GEN_6564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6566 = 8'h42 == r_count_31_io_out ? io_r_66_b : _GEN_6565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6567 = 8'h43 == r_count_31_io_out ? io_r_67_b : _GEN_6566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6568 = 8'h44 == r_count_31_io_out ? io_r_68_b : _GEN_6567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6569 = 8'h45 == r_count_31_io_out ? io_r_69_b : _GEN_6568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6570 = 8'h46 == r_count_31_io_out ? io_r_70_b : _GEN_6569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6571 = 8'h47 == r_count_31_io_out ? io_r_71_b : _GEN_6570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6572 = 8'h48 == r_count_31_io_out ? io_r_72_b : _GEN_6571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6573 = 8'h49 == r_count_31_io_out ? io_r_73_b : _GEN_6572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6574 = 8'h4a == r_count_31_io_out ? io_r_74_b : _GEN_6573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6575 = 8'h4b == r_count_31_io_out ? io_r_75_b : _GEN_6574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6576 = 8'h4c == r_count_31_io_out ? io_r_76_b : _GEN_6575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6577 = 8'h4d == r_count_31_io_out ? io_r_77_b : _GEN_6576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6578 = 8'h4e == r_count_31_io_out ? io_r_78_b : _GEN_6577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6579 = 8'h4f == r_count_31_io_out ? io_r_79_b : _GEN_6578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6580 = 8'h50 == r_count_31_io_out ? io_r_80_b : _GEN_6579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6581 = 8'h51 == r_count_31_io_out ? io_r_81_b : _GEN_6580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6582 = 8'h52 == r_count_31_io_out ? io_r_82_b : _GEN_6581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6583 = 8'h53 == r_count_31_io_out ? io_r_83_b : _GEN_6582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6584 = 8'h54 == r_count_31_io_out ? io_r_84_b : _GEN_6583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6585 = 8'h55 == r_count_31_io_out ? io_r_85_b : _GEN_6584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6586 = 8'h56 == r_count_31_io_out ? io_r_86_b : _GEN_6585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6587 = 8'h57 == r_count_31_io_out ? io_r_87_b : _GEN_6586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6588 = 8'h58 == r_count_31_io_out ? io_r_88_b : _GEN_6587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6589 = 8'h59 == r_count_31_io_out ? io_r_89_b : _GEN_6588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6590 = 8'h5a == r_count_31_io_out ? io_r_90_b : _GEN_6589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6591 = 8'h5b == r_count_31_io_out ? io_r_91_b : _GEN_6590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6592 = 8'h5c == r_count_31_io_out ? io_r_92_b : _GEN_6591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6593 = 8'h5d == r_count_31_io_out ? io_r_93_b : _GEN_6592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6594 = 8'h5e == r_count_31_io_out ? io_r_94_b : _GEN_6593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6595 = 8'h5f == r_count_31_io_out ? io_r_95_b : _GEN_6594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6596 = 8'h60 == r_count_31_io_out ? io_r_96_b : _GEN_6595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6597 = 8'h61 == r_count_31_io_out ? io_r_97_b : _GEN_6596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6598 = 8'h62 == r_count_31_io_out ? io_r_98_b : _GEN_6597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6599 = 8'h63 == r_count_31_io_out ? io_r_99_b : _GEN_6598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6600 = 8'h64 == r_count_31_io_out ? io_r_100_b : _GEN_6599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6601 = 8'h65 == r_count_31_io_out ? io_r_101_b : _GEN_6600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6602 = 8'h66 == r_count_31_io_out ? io_r_102_b : _GEN_6601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6603 = 8'h67 == r_count_31_io_out ? io_r_103_b : _GEN_6602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6604 = 8'h68 == r_count_31_io_out ? io_r_104_b : _GEN_6603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6605 = 8'h69 == r_count_31_io_out ? io_r_105_b : _GEN_6604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6606 = 8'h6a == r_count_31_io_out ? io_r_106_b : _GEN_6605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6607 = 8'h6b == r_count_31_io_out ? io_r_107_b : _GEN_6606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6608 = 8'h6c == r_count_31_io_out ? io_r_108_b : _GEN_6607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6609 = 8'h6d == r_count_31_io_out ? io_r_109_b : _GEN_6608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6610 = 8'h6e == r_count_31_io_out ? io_r_110_b : _GEN_6609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6611 = 8'h6f == r_count_31_io_out ? io_r_111_b : _GEN_6610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6612 = 8'h70 == r_count_31_io_out ? io_r_112_b : _GEN_6611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6613 = 8'h71 == r_count_31_io_out ? io_r_113_b : _GEN_6612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6614 = 8'h72 == r_count_31_io_out ? io_r_114_b : _GEN_6613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6615 = 8'h73 == r_count_31_io_out ? io_r_115_b : _GEN_6614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6616 = 8'h74 == r_count_31_io_out ? io_r_116_b : _GEN_6615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6617 = 8'h75 == r_count_31_io_out ? io_r_117_b : _GEN_6616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6618 = 8'h76 == r_count_31_io_out ? io_r_118_b : _GEN_6617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6619 = 8'h77 == r_count_31_io_out ? io_r_119_b : _GEN_6618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6620 = 8'h78 == r_count_31_io_out ? io_r_120_b : _GEN_6619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6621 = 8'h79 == r_count_31_io_out ? io_r_121_b : _GEN_6620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6622 = 8'h7a == r_count_31_io_out ? io_r_122_b : _GEN_6621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6623 = 8'h7b == r_count_31_io_out ? io_r_123_b : _GEN_6622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6624 = 8'h7c == r_count_31_io_out ? io_r_124_b : _GEN_6623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6625 = 8'h7d == r_count_31_io_out ? io_r_125_b : _GEN_6624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6626 = 8'h7e == r_count_31_io_out ? io_r_126_b : _GEN_6625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6627 = 8'h7f == r_count_31_io_out ? io_r_127_b : _GEN_6626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6628 = 8'h80 == r_count_31_io_out ? io_r_128_b : _GEN_6627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6629 = 8'h81 == r_count_31_io_out ? io_r_129_b : _GEN_6628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6630 = 8'h82 == r_count_31_io_out ? io_r_130_b : _GEN_6629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6631 = 8'h83 == r_count_31_io_out ? io_r_131_b : _GEN_6630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6632 = 8'h84 == r_count_31_io_out ? io_r_132_b : _GEN_6631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6633 = 8'h85 == r_count_31_io_out ? io_r_133_b : _GEN_6632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6634 = 8'h86 == r_count_31_io_out ? io_r_134_b : _GEN_6633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6635 = 8'h87 == r_count_31_io_out ? io_r_135_b : _GEN_6634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6636 = 8'h88 == r_count_31_io_out ? io_r_136_b : _GEN_6635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6637 = 8'h89 == r_count_31_io_out ? io_r_137_b : _GEN_6636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6638 = 8'h8a == r_count_31_io_out ? io_r_138_b : _GEN_6637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6639 = 8'h8b == r_count_31_io_out ? io_r_139_b : _GEN_6638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6640 = 8'h8c == r_count_31_io_out ? io_r_140_b : _GEN_6639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6641 = 8'h8d == r_count_31_io_out ? io_r_141_b : _GEN_6640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6642 = 8'h8e == r_count_31_io_out ? io_r_142_b : _GEN_6641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6643 = 8'h8f == r_count_31_io_out ? io_r_143_b : _GEN_6642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6644 = 8'h90 == r_count_31_io_out ? io_r_144_b : _GEN_6643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6645 = 8'h91 == r_count_31_io_out ? io_r_145_b : _GEN_6644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6646 = 8'h92 == r_count_31_io_out ? io_r_146_b : _GEN_6645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6647 = 8'h93 == r_count_31_io_out ? io_r_147_b : _GEN_6646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6648 = 8'h94 == r_count_31_io_out ? io_r_148_b : _GEN_6647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6649 = 8'h95 == r_count_31_io_out ? io_r_149_b : _GEN_6648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6650 = 8'h96 == r_count_31_io_out ? io_r_150_b : _GEN_6649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6651 = 8'h97 == r_count_31_io_out ? io_r_151_b : _GEN_6650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6652 = 8'h98 == r_count_31_io_out ? io_r_152_b : _GEN_6651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6653 = 8'h99 == r_count_31_io_out ? io_r_153_b : _GEN_6652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6654 = 8'h9a == r_count_31_io_out ? io_r_154_b : _GEN_6653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6655 = 8'h9b == r_count_31_io_out ? io_r_155_b : _GEN_6654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6656 = 8'h9c == r_count_31_io_out ? io_r_156_b : _GEN_6655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6657 = 8'h9d == r_count_31_io_out ? io_r_157_b : _GEN_6656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6658 = 8'h9e == r_count_31_io_out ? io_r_158_b : _GEN_6657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6659 = 8'h9f == r_count_31_io_out ? io_r_159_b : _GEN_6658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6660 = 8'ha0 == r_count_31_io_out ? io_r_160_b : _GEN_6659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6661 = 8'ha1 == r_count_31_io_out ? io_r_161_b : _GEN_6660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6662 = 8'ha2 == r_count_31_io_out ? io_r_162_b : _GEN_6661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6663 = 8'ha3 == r_count_31_io_out ? io_r_163_b : _GEN_6662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6664 = 8'ha4 == r_count_31_io_out ? io_r_164_b : _GEN_6663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6665 = 8'ha5 == r_count_31_io_out ? io_r_165_b : _GEN_6664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6666 = 8'ha6 == r_count_31_io_out ? io_r_166_b : _GEN_6665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6667 = 8'ha7 == r_count_31_io_out ? io_r_167_b : _GEN_6666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6668 = 8'ha8 == r_count_31_io_out ? io_r_168_b : _GEN_6667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6669 = 8'ha9 == r_count_31_io_out ? io_r_169_b : _GEN_6668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6670 = 8'haa == r_count_31_io_out ? io_r_170_b : _GEN_6669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6671 = 8'hab == r_count_31_io_out ? io_r_171_b : _GEN_6670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6672 = 8'hac == r_count_31_io_out ? io_r_172_b : _GEN_6671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6673 = 8'had == r_count_31_io_out ? io_r_173_b : _GEN_6672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6674 = 8'hae == r_count_31_io_out ? io_r_174_b : _GEN_6673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6675 = 8'haf == r_count_31_io_out ? io_r_175_b : _GEN_6674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6676 = 8'hb0 == r_count_31_io_out ? io_r_176_b : _GEN_6675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6677 = 8'hb1 == r_count_31_io_out ? io_r_177_b : _GEN_6676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6678 = 8'hb2 == r_count_31_io_out ? io_r_178_b : _GEN_6677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6679 = 8'hb3 == r_count_31_io_out ? io_r_179_b : _GEN_6678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6680 = 8'hb4 == r_count_31_io_out ? io_r_180_b : _GEN_6679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6681 = 8'hb5 == r_count_31_io_out ? io_r_181_b : _GEN_6680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6682 = 8'hb6 == r_count_31_io_out ? io_r_182_b : _GEN_6681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6683 = 8'hb7 == r_count_31_io_out ? io_r_183_b : _GEN_6682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6684 = 8'hb8 == r_count_31_io_out ? io_r_184_b : _GEN_6683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6685 = 8'hb9 == r_count_31_io_out ? io_r_185_b : _GEN_6684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6686 = 8'hba == r_count_31_io_out ? io_r_186_b : _GEN_6685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6687 = 8'hbb == r_count_31_io_out ? io_r_187_b : _GEN_6686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6688 = 8'hbc == r_count_31_io_out ? io_r_188_b : _GEN_6687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6689 = 8'hbd == r_count_31_io_out ? io_r_189_b : _GEN_6688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6690 = 8'hbe == r_count_31_io_out ? io_r_190_b : _GEN_6689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6691 = 8'hbf == r_count_31_io_out ? io_r_191_b : _GEN_6690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6692 = 8'hc0 == r_count_31_io_out ? io_r_192_b : _GEN_6691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6693 = 8'hc1 == r_count_31_io_out ? io_r_193_b : _GEN_6692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6694 = 8'hc2 == r_count_31_io_out ? io_r_194_b : _GEN_6693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6695 = 8'hc3 == r_count_31_io_out ? io_r_195_b : _GEN_6694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6696 = 8'hc4 == r_count_31_io_out ? io_r_196_b : _GEN_6695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6697 = 8'hc5 == r_count_31_io_out ? io_r_197_b : _GEN_6696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6698 = 8'hc6 == r_count_31_io_out ? io_r_198_b : _GEN_6697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6701 = 8'h1 == r_count_32_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6702 = 8'h2 == r_count_32_io_out ? io_r_2_b : _GEN_6701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6703 = 8'h3 == r_count_32_io_out ? io_r_3_b : _GEN_6702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6704 = 8'h4 == r_count_32_io_out ? io_r_4_b : _GEN_6703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6705 = 8'h5 == r_count_32_io_out ? io_r_5_b : _GEN_6704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6706 = 8'h6 == r_count_32_io_out ? io_r_6_b : _GEN_6705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6707 = 8'h7 == r_count_32_io_out ? io_r_7_b : _GEN_6706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6708 = 8'h8 == r_count_32_io_out ? io_r_8_b : _GEN_6707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6709 = 8'h9 == r_count_32_io_out ? io_r_9_b : _GEN_6708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6710 = 8'ha == r_count_32_io_out ? io_r_10_b : _GEN_6709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6711 = 8'hb == r_count_32_io_out ? io_r_11_b : _GEN_6710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6712 = 8'hc == r_count_32_io_out ? io_r_12_b : _GEN_6711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6713 = 8'hd == r_count_32_io_out ? io_r_13_b : _GEN_6712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6714 = 8'he == r_count_32_io_out ? io_r_14_b : _GEN_6713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6715 = 8'hf == r_count_32_io_out ? io_r_15_b : _GEN_6714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6716 = 8'h10 == r_count_32_io_out ? io_r_16_b : _GEN_6715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6717 = 8'h11 == r_count_32_io_out ? io_r_17_b : _GEN_6716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6718 = 8'h12 == r_count_32_io_out ? io_r_18_b : _GEN_6717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6719 = 8'h13 == r_count_32_io_out ? io_r_19_b : _GEN_6718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6720 = 8'h14 == r_count_32_io_out ? io_r_20_b : _GEN_6719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6721 = 8'h15 == r_count_32_io_out ? io_r_21_b : _GEN_6720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6722 = 8'h16 == r_count_32_io_out ? io_r_22_b : _GEN_6721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6723 = 8'h17 == r_count_32_io_out ? io_r_23_b : _GEN_6722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6724 = 8'h18 == r_count_32_io_out ? io_r_24_b : _GEN_6723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6725 = 8'h19 == r_count_32_io_out ? io_r_25_b : _GEN_6724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6726 = 8'h1a == r_count_32_io_out ? io_r_26_b : _GEN_6725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6727 = 8'h1b == r_count_32_io_out ? io_r_27_b : _GEN_6726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6728 = 8'h1c == r_count_32_io_out ? io_r_28_b : _GEN_6727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6729 = 8'h1d == r_count_32_io_out ? io_r_29_b : _GEN_6728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6730 = 8'h1e == r_count_32_io_out ? io_r_30_b : _GEN_6729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6731 = 8'h1f == r_count_32_io_out ? io_r_31_b : _GEN_6730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6732 = 8'h20 == r_count_32_io_out ? io_r_32_b : _GEN_6731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6733 = 8'h21 == r_count_32_io_out ? io_r_33_b : _GEN_6732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6734 = 8'h22 == r_count_32_io_out ? io_r_34_b : _GEN_6733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6735 = 8'h23 == r_count_32_io_out ? io_r_35_b : _GEN_6734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6736 = 8'h24 == r_count_32_io_out ? io_r_36_b : _GEN_6735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6737 = 8'h25 == r_count_32_io_out ? io_r_37_b : _GEN_6736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6738 = 8'h26 == r_count_32_io_out ? io_r_38_b : _GEN_6737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6739 = 8'h27 == r_count_32_io_out ? io_r_39_b : _GEN_6738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6740 = 8'h28 == r_count_32_io_out ? io_r_40_b : _GEN_6739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6741 = 8'h29 == r_count_32_io_out ? io_r_41_b : _GEN_6740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6742 = 8'h2a == r_count_32_io_out ? io_r_42_b : _GEN_6741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6743 = 8'h2b == r_count_32_io_out ? io_r_43_b : _GEN_6742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6744 = 8'h2c == r_count_32_io_out ? io_r_44_b : _GEN_6743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6745 = 8'h2d == r_count_32_io_out ? io_r_45_b : _GEN_6744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6746 = 8'h2e == r_count_32_io_out ? io_r_46_b : _GEN_6745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6747 = 8'h2f == r_count_32_io_out ? io_r_47_b : _GEN_6746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6748 = 8'h30 == r_count_32_io_out ? io_r_48_b : _GEN_6747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6749 = 8'h31 == r_count_32_io_out ? io_r_49_b : _GEN_6748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6750 = 8'h32 == r_count_32_io_out ? io_r_50_b : _GEN_6749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6751 = 8'h33 == r_count_32_io_out ? io_r_51_b : _GEN_6750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6752 = 8'h34 == r_count_32_io_out ? io_r_52_b : _GEN_6751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6753 = 8'h35 == r_count_32_io_out ? io_r_53_b : _GEN_6752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6754 = 8'h36 == r_count_32_io_out ? io_r_54_b : _GEN_6753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6755 = 8'h37 == r_count_32_io_out ? io_r_55_b : _GEN_6754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6756 = 8'h38 == r_count_32_io_out ? io_r_56_b : _GEN_6755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6757 = 8'h39 == r_count_32_io_out ? io_r_57_b : _GEN_6756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6758 = 8'h3a == r_count_32_io_out ? io_r_58_b : _GEN_6757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6759 = 8'h3b == r_count_32_io_out ? io_r_59_b : _GEN_6758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6760 = 8'h3c == r_count_32_io_out ? io_r_60_b : _GEN_6759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6761 = 8'h3d == r_count_32_io_out ? io_r_61_b : _GEN_6760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6762 = 8'h3e == r_count_32_io_out ? io_r_62_b : _GEN_6761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6763 = 8'h3f == r_count_32_io_out ? io_r_63_b : _GEN_6762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6764 = 8'h40 == r_count_32_io_out ? io_r_64_b : _GEN_6763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6765 = 8'h41 == r_count_32_io_out ? io_r_65_b : _GEN_6764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6766 = 8'h42 == r_count_32_io_out ? io_r_66_b : _GEN_6765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6767 = 8'h43 == r_count_32_io_out ? io_r_67_b : _GEN_6766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6768 = 8'h44 == r_count_32_io_out ? io_r_68_b : _GEN_6767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6769 = 8'h45 == r_count_32_io_out ? io_r_69_b : _GEN_6768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6770 = 8'h46 == r_count_32_io_out ? io_r_70_b : _GEN_6769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6771 = 8'h47 == r_count_32_io_out ? io_r_71_b : _GEN_6770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6772 = 8'h48 == r_count_32_io_out ? io_r_72_b : _GEN_6771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6773 = 8'h49 == r_count_32_io_out ? io_r_73_b : _GEN_6772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6774 = 8'h4a == r_count_32_io_out ? io_r_74_b : _GEN_6773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6775 = 8'h4b == r_count_32_io_out ? io_r_75_b : _GEN_6774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6776 = 8'h4c == r_count_32_io_out ? io_r_76_b : _GEN_6775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6777 = 8'h4d == r_count_32_io_out ? io_r_77_b : _GEN_6776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6778 = 8'h4e == r_count_32_io_out ? io_r_78_b : _GEN_6777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6779 = 8'h4f == r_count_32_io_out ? io_r_79_b : _GEN_6778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6780 = 8'h50 == r_count_32_io_out ? io_r_80_b : _GEN_6779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6781 = 8'h51 == r_count_32_io_out ? io_r_81_b : _GEN_6780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6782 = 8'h52 == r_count_32_io_out ? io_r_82_b : _GEN_6781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6783 = 8'h53 == r_count_32_io_out ? io_r_83_b : _GEN_6782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6784 = 8'h54 == r_count_32_io_out ? io_r_84_b : _GEN_6783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6785 = 8'h55 == r_count_32_io_out ? io_r_85_b : _GEN_6784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6786 = 8'h56 == r_count_32_io_out ? io_r_86_b : _GEN_6785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6787 = 8'h57 == r_count_32_io_out ? io_r_87_b : _GEN_6786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6788 = 8'h58 == r_count_32_io_out ? io_r_88_b : _GEN_6787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6789 = 8'h59 == r_count_32_io_out ? io_r_89_b : _GEN_6788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6790 = 8'h5a == r_count_32_io_out ? io_r_90_b : _GEN_6789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6791 = 8'h5b == r_count_32_io_out ? io_r_91_b : _GEN_6790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6792 = 8'h5c == r_count_32_io_out ? io_r_92_b : _GEN_6791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6793 = 8'h5d == r_count_32_io_out ? io_r_93_b : _GEN_6792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6794 = 8'h5e == r_count_32_io_out ? io_r_94_b : _GEN_6793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6795 = 8'h5f == r_count_32_io_out ? io_r_95_b : _GEN_6794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6796 = 8'h60 == r_count_32_io_out ? io_r_96_b : _GEN_6795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6797 = 8'h61 == r_count_32_io_out ? io_r_97_b : _GEN_6796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6798 = 8'h62 == r_count_32_io_out ? io_r_98_b : _GEN_6797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6799 = 8'h63 == r_count_32_io_out ? io_r_99_b : _GEN_6798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6800 = 8'h64 == r_count_32_io_out ? io_r_100_b : _GEN_6799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6801 = 8'h65 == r_count_32_io_out ? io_r_101_b : _GEN_6800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6802 = 8'h66 == r_count_32_io_out ? io_r_102_b : _GEN_6801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6803 = 8'h67 == r_count_32_io_out ? io_r_103_b : _GEN_6802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6804 = 8'h68 == r_count_32_io_out ? io_r_104_b : _GEN_6803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6805 = 8'h69 == r_count_32_io_out ? io_r_105_b : _GEN_6804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6806 = 8'h6a == r_count_32_io_out ? io_r_106_b : _GEN_6805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6807 = 8'h6b == r_count_32_io_out ? io_r_107_b : _GEN_6806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6808 = 8'h6c == r_count_32_io_out ? io_r_108_b : _GEN_6807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6809 = 8'h6d == r_count_32_io_out ? io_r_109_b : _GEN_6808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6810 = 8'h6e == r_count_32_io_out ? io_r_110_b : _GEN_6809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6811 = 8'h6f == r_count_32_io_out ? io_r_111_b : _GEN_6810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6812 = 8'h70 == r_count_32_io_out ? io_r_112_b : _GEN_6811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6813 = 8'h71 == r_count_32_io_out ? io_r_113_b : _GEN_6812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6814 = 8'h72 == r_count_32_io_out ? io_r_114_b : _GEN_6813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6815 = 8'h73 == r_count_32_io_out ? io_r_115_b : _GEN_6814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6816 = 8'h74 == r_count_32_io_out ? io_r_116_b : _GEN_6815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6817 = 8'h75 == r_count_32_io_out ? io_r_117_b : _GEN_6816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6818 = 8'h76 == r_count_32_io_out ? io_r_118_b : _GEN_6817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6819 = 8'h77 == r_count_32_io_out ? io_r_119_b : _GEN_6818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6820 = 8'h78 == r_count_32_io_out ? io_r_120_b : _GEN_6819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6821 = 8'h79 == r_count_32_io_out ? io_r_121_b : _GEN_6820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6822 = 8'h7a == r_count_32_io_out ? io_r_122_b : _GEN_6821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6823 = 8'h7b == r_count_32_io_out ? io_r_123_b : _GEN_6822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6824 = 8'h7c == r_count_32_io_out ? io_r_124_b : _GEN_6823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6825 = 8'h7d == r_count_32_io_out ? io_r_125_b : _GEN_6824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6826 = 8'h7e == r_count_32_io_out ? io_r_126_b : _GEN_6825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6827 = 8'h7f == r_count_32_io_out ? io_r_127_b : _GEN_6826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6828 = 8'h80 == r_count_32_io_out ? io_r_128_b : _GEN_6827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6829 = 8'h81 == r_count_32_io_out ? io_r_129_b : _GEN_6828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6830 = 8'h82 == r_count_32_io_out ? io_r_130_b : _GEN_6829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6831 = 8'h83 == r_count_32_io_out ? io_r_131_b : _GEN_6830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6832 = 8'h84 == r_count_32_io_out ? io_r_132_b : _GEN_6831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6833 = 8'h85 == r_count_32_io_out ? io_r_133_b : _GEN_6832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6834 = 8'h86 == r_count_32_io_out ? io_r_134_b : _GEN_6833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6835 = 8'h87 == r_count_32_io_out ? io_r_135_b : _GEN_6834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6836 = 8'h88 == r_count_32_io_out ? io_r_136_b : _GEN_6835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6837 = 8'h89 == r_count_32_io_out ? io_r_137_b : _GEN_6836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6838 = 8'h8a == r_count_32_io_out ? io_r_138_b : _GEN_6837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6839 = 8'h8b == r_count_32_io_out ? io_r_139_b : _GEN_6838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6840 = 8'h8c == r_count_32_io_out ? io_r_140_b : _GEN_6839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6841 = 8'h8d == r_count_32_io_out ? io_r_141_b : _GEN_6840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6842 = 8'h8e == r_count_32_io_out ? io_r_142_b : _GEN_6841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6843 = 8'h8f == r_count_32_io_out ? io_r_143_b : _GEN_6842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6844 = 8'h90 == r_count_32_io_out ? io_r_144_b : _GEN_6843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6845 = 8'h91 == r_count_32_io_out ? io_r_145_b : _GEN_6844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6846 = 8'h92 == r_count_32_io_out ? io_r_146_b : _GEN_6845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6847 = 8'h93 == r_count_32_io_out ? io_r_147_b : _GEN_6846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6848 = 8'h94 == r_count_32_io_out ? io_r_148_b : _GEN_6847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6849 = 8'h95 == r_count_32_io_out ? io_r_149_b : _GEN_6848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6850 = 8'h96 == r_count_32_io_out ? io_r_150_b : _GEN_6849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6851 = 8'h97 == r_count_32_io_out ? io_r_151_b : _GEN_6850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6852 = 8'h98 == r_count_32_io_out ? io_r_152_b : _GEN_6851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6853 = 8'h99 == r_count_32_io_out ? io_r_153_b : _GEN_6852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6854 = 8'h9a == r_count_32_io_out ? io_r_154_b : _GEN_6853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6855 = 8'h9b == r_count_32_io_out ? io_r_155_b : _GEN_6854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6856 = 8'h9c == r_count_32_io_out ? io_r_156_b : _GEN_6855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6857 = 8'h9d == r_count_32_io_out ? io_r_157_b : _GEN_6856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6858 = 8'h9e == r_count_32_io_out ? io_r_158_b : _GEN_6857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6859 = 8'h9f == r_count_32_io_out ? io_r_159_b : _GEN_6858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6860 = 8'ha0 == r_count_32_io_out ? io_r_160_b : _GEN_6859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6861 = 8'ha1 == r_count_32_io_out ? io_r_161_b : _GEN_6860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6862 = 8'ha2 == r_count_32_io_out ? io_r_162_b : _GEN_6861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6863 = 8'ha3 == r_count_32_io_out ? io_r_163_b : _GEN_6862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6864 = 8'ha4 == r_count_32_io_out ? io_r_164_b : _GEN_6863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6865 = 8'ha5 == r_count_32_io_out ? io_r_165_b : _GEN_6864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6866 = 8'ha6 == r_count_32_io_out ? io_r_166_b : _GEN_6865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6867 = 8'ha7 == r_count_32_io_out ? io_r_167_b : _GEN_6866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6868 = 8'ha8 == r_count_32_io_out ? io_r_168_b : _GEN_6867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6869 = 8'ha9 == r_count_32_io_out ? io_r_169_b : _GEN_6868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6870 = 8'haa == r_count_32_io_out ? io_r_170_b : _GEN_6869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6871 = 8'hab == r_count_32_io_out ? io_r_171_b : _GEN_6870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6872 = 8'hac == r_count_32_io_out ? io_r_172_b : _GEN_6871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6873 = 8'had == r_count_32_io_out ? io_r_173_b : _GEN_6872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6874 = 8'hae == r_count_32_io_out ? io_r_174_b : _GEN_6873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6875 = 8'haf == r_count_32_io_out ? io_r_175_b : _GEN_6874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6876 = 8'hb0 == r_count_32_io_out ? io_r_176_b : _GEN_6875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6877 = 8'hb1 == r_count_32_io_out ? io_r_177_b : _GEN_6876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6878 = 8'hb2 == r_count_32_io_out ? io_r_178_b : _GEN_6877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6879 = 8'hb3 == r_count_32_io_out ? io_r_179_b : _GEN_6878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6880 = 8'hb4 == r_count_32_io_out ? io_r_180_b : _GEN_6879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6881 = 8'hb5 == r_count_32_io_out ? io_r_181_b : _GEN_6880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6882 = 8'hb6 == r_count_32_io_out ? io_r_182_b : _GEN_6881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6883 = 8'hb7 == r_count_32_io_out ? io_r_183_b : _GEN_6882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6884 = 8'hb8 == r_count_32_io_out ? io_r_184_b : _GEN_6883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6885 = 8'hb9 == r_count_32_io_out ? io_r_185_b : _GEN_6884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6886 = 8'hba == r_count_32_io_out ? io_r_186_b : _GEN_6885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6887 = 8'hbb == r_count_32_io_out ? io_r_187_b : _GEN_6886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6888 = 8'hbc == r_count_32_io_out ? io_r_188_b : _GEN_6887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6889 = 8'hbd == r_count_32_io_out ? io_r_189_b : _GEN_6888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6890 = 8'hbe == r_count_32_io_out ? io_r_190_b : _GEN_6889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6891 = 8'hbf == r_count_32_io_out ? io_r_191_b : _GEN_6890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6892 = 8'hc0 == r_count_32_io_out ? io_r_192_b : _GEN_6891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6893 = 8'hc1 == r_count_32_io_out ? io_r_193_b : _GEN_6892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6894 = 8'hc2 == r_count_32_io_out ? io_r_194_b : _GEN_6893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6895 = 8'hc3 == r_count_32_io_out ? io_r_195_b : _GEN_6894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6896 = 8'hc4 == r_count_32_io_out ? io_r_196_b : _GEN_6895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6897 = 8'hc5 == r_count_32_io_out ? io_r_197_b : _GEN_6896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6898 = 8'hc6 == r_count_32_io_out ? io_r_198_b : _GEN_6897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6901 = 8'h1 == r_count_33_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6902 = 8'h2 == r_count_33_io_out ? io_r_2_b : _GEN_6901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6903 = 8'h3 == r_count_33_io_out ? io_r_3_b : _GEN_6902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6904 = 8'h4 == r_count_33_io_out ? io_r_4_b : _GEN_6903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6905 = 8'h5 == r_count_33_io_out ? io_r_5_b : _GEN_6904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6906 = 8'h6 == r_count_33_io_out ? io_r_6_b : _GEN_6905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6907 = 8'h7 == r_count_33_io_out ? io_r_7_b : _GEN_6906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6908 = 8'h8 == r_count_33_io_out ? io_r_8_b : _GEN_6907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6909 = 8'h9 == r_count_33_io_out ? io_r_9_b : _GEN_6908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6910 = 8'ha == r_count_33_io_out ? io_r_10_b : _GEN_6909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6911 = 8'hb == r_count_33_io_out ? io_r_11_b : _GEN_6910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6912 = 8'hc == r_count_33_io_out ? io_r_12_b : _GEN_6911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6913 = 8'hd == r_count_33_io_out ? io_r_13_b : _GEN_6912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6914 = 8'he == r_count_33_io_out ? io_r_14_b : _GEN_6913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6915 = 8'hf == r_count_33_io_out ? io_r_15_b : _GEN_6914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6916 = 8'h10 == r_count_33_io_out ? io_r_16_b : _GEN_6915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6917 = 8'h11 == r_count_33_io_out ? io_r_17_b : _GEN_6916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6918 = 8'h12 == r_count_33_io_out ? io_r_18_b : _GEN_6917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6919 = 8'h13 == r_count_33_io_out ? io_r_19_b : _GEN_6918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6920 = 8'h14 == r_count_33_io_out ? io_r_20_b : _GEN_6919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6921 = 8'h15 == r_count_33_io_out ? io_r_21_b : _GEN_6920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6922 = 8'h16 == r_count_33_io_out ? io_r_22_b : _GEN_6921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6923 = 8'h17 == r_count_33_io_out ? io_r_23_b : _GEN_6922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6924 = 8'h18 == r_count_33_io_out ? io_r_24_b : _GEN_6923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6925 = 8'h19 == r_count_33_io_out ? io_r_25_b : _GEN_6924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6926 = 8'h1a == r_count_33_io_out ? io_r_26_b : _GEN_6925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6927 = 8'h1b == r_count_33_io_out ? io_r_27_b : _GEN_6926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6928 = 8'h1c == r_count_33_io_out ? io_r_28_b : _GEN_6927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6929 = 8'h1d == r_count_33_io_out ? io_r_29_b : _GEN_6928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6930 = 8'h1e == r_count_33_io_out ? io_r_30_b : _GEN_6929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6931 = 8'h1f == r_count_33_io_out ? io_r_31_b : _GEN_6930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6932 = 8'h20 == r_count_33_io_out ? io_r_32_b : _GEN_6931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6933 = 8'h21 == r_count_33_io_out ? io_r_33_b : _GEN_6932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6934 = 8'h22 == r_count_33_io_out ? io_r_34_b : _GEN_6933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6935 = 8'h23 == r_count_33_io_out ? io_r_35_b : _GEN_6934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6936 = 8'h24 == r_count_33_io_out ? io_r_36_b : _GEN_6935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6937 = 8'h25 == r_count_33_io_out ? io_r_37_b : _GEN_6936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6938 = 8'h26 == r_count_33_io_out ? io_r_38_b : _GEN_6937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6939 = 8'h27 == r_count_33_io_out ? io_r_39_b : _GEN_6938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6940 = 8'h28 == r_count_33_io_out ? io_r_40_b : _GEN_6939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6941 = 8'h29 == r_count_33_io_out ? io_r_41_b : _GEN_6940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6942 = 8'h2a == r_count_33_io_out ? io_r_42_b : _GEN_6941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6943 = 8'h2b == r_count_33_io_out ? io_r_43_b : _GEN_6942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6944 = 8'h2c == r_count_33_io_out ? io_r_44_b : _GEN_6943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6945 = 8'h2d == r_count_33_io_out ? io_r_45_b : _GEN_6944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6946 = 8'h2e == r_count_33_io_out ? io_r_46_b : _GEN_6945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6947 = 8'h2f == r_count_33_io_out ? io_r_47_b : _GEN_6946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6948 = 8'h30 == r_count_33_io_out ? io_r_48_b : _GEN_6947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6949 = 8'h31 == r_count_33_io_out ? io_r_49_b : _GEN_6948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6950 = 8'h32 == r_count_33_io_out ? io_r_50_b : _GEN_6949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6951 = 8'h33 == r_count_33_io_out ? io_r_51_b : _GEN_6950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6952 = 8'h34 == r_count_33_io_out ? io_r_52_b : _GEN_6951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6953 = 8'h35 == r_count_33_io_out ? io_r_53_b : _GEN_6952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6954 = 8'h36 == r_count_33_io_out ? io_r_54_b : _GEN_6953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6955 = 8'h37 == r_count_33_io_out ? io_r_55_b : _GEN_6954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6956 = 8'h38 == r_count_33_io_out ? io_r_56_b : _GEN_6955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6957 = 8'h39 == r_count_33_io_out ? io_r_57_b : _GEN_6956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6958 = 8'h3a == r_count_33_io_out ? io_r_58_b : _GEN_6957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6959 = 8'h3b == r_count_33_io_out ? io_r_59_b : _GEN_6958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6960 = 8'h3c == r_count_33_io_out ? io_r_60_b : _GEN_6959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6961 = 8'h3d == r_count_33_io_out ? io_r_61_b : _GEN_6960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6962 = 8'h3e == r_count_33_io_out ? io_r_62_b : _GEN_6961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6963 = 8'h3f == r_count_33_io_out ? io_r_63_b : _GEN_6962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6964 = 8'h40 == r_count_33_io_out ? io_r_64_b : _GEN_6963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6965 = 8'h41 == r_count_33_io_out ? io_r_65_b : _GEN_6964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6966 = 8'h42 == r_count_33_io_out ? io_r_66_b : _GEN_6965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6967 = 8'h43 == r_count_33_io_out ? io_r_67_b : _GEN_6966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6968 = 8'h44 == r_count_33_io_out ? io_r_68_b : _GEN_6967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6969 = 8'h45 == r_count_33_io_out ? io_r_69_b : _GEN_6968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6970 = 8'h46 == r_count_33_io_out ? io_r_70_b : _GEN_6969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6971 = 8'h47 == r_count_33_io_out ? io_r_71_b : _GEN_6970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6972 = 8'h48 == r_count_33_io_out ? io_r_72_b : _GEN_6971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6973 = 8'h49 == r_count_33_io_out ? io_r_73_b : _GEN_6972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6974 = 8'h4a == r_count_33_io_out ? io_r_74_b : _GEN_6973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6975 = 8'h4b == r_count_33_io_out ? io_r_75_b : _GEN_6974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6976 = 8'h4c == r_count_33_io_out ? io_r_76_b : _GEN_6975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6977 = 8'h4d == r_count_33_io_out ? io_r_77_b : _GEN_6976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6978 = 8'h4e == r_count_33_io_out ? io_r_78_b : _GEN_6977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6979 = 8'h4f == r_count_33_io_out ? io_r_79_b : _GEN_6978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6980 = 8'h50 == r_count_33_io_out ? io_r_80_b : _GEN_6979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6981 = 8'h51 == r_count_33_io_out ? io_r_81_b : _GEN_6980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6982 = 8'h52 == r_count_33_io_out ? io_r_82_b : _GEN_6981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6983 = 8'h53 == r_count_33_io_out ? io_r_83_b : _GEN_6982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6984 = 8'h54 == r_count_33_io_out ? io_r_84_b : _GEN_6983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6985 = 8'h55 == r_count_33_io_out ? io_r_85_b : _GEN_6984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6986 = 8'h56 == r_count_33_io_out ? io_r_86_b : _GEN_6985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6987 = 8'h57 == r_count_33_io_out ? io_r_87_b : _GEN_6986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6988 = 8'h58 == r_count_33_io_out ? io_r_88_b : _GEN_6987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6989 = 8'h59 == r_count_33_io_out ? io_r_89_b : _GEN_6988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6990 = 8'h5a == r_count_33_io_out ? io_r_90_b : _GEN_6989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6991 = 8'h5b == r_count_33_io_out ? io_r_91_b : _GEN_6990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6992 = 8'h5c == r_count_33_io_out ? io_r_92_b : _GEN_6991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6993 = 8'h5d == r_count_33_io_out ? io_r_93_b : _GEN_6992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6994 = 8'h5e == r_count_33_io_out ? io_r_94_b : _GEN_6993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6995 = 8'h5f == r_count_33_io_out ? io_r_95_b : _GEN_6994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6996 = 8'h60 == r_count_33_io_out ? io_r_96_b : _GEN_6995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6997 = 8'h61 == r_count_33_io_out ? io_r_97_b : _GEN_6996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6998 = 8'h62 == r_count_33_io_out ? io_r_98_b : _GEN_6997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6999 = 8'h63 == r_count_33_io_out ? io_r_99_b : _GEN_6998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7000 = 8'h64 == r_count_33_io_out ? io_r_100_b : _GEN_6999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7001 = 8'h65 == r_count_33_io_out ? io_r_101_b : _GEN_7000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7002 = 8'h66 == r_count_33_io_out ? io_r_102_b : _GEN_7001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7003 = 8'h67 == r_count_33_io_out ? io_r_103_b : _GEN_7002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7004 = 8'h68 == r_count_33_io_out ? io_r_104_b : _GEN_7003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7005 = 8'h69 == r_count_33_io_out ? io_r_105_b : _GEN_7004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7006 = 8'h6a == r_count_33_io_out ? io_r_106_b : _GEN_7005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7007 = 8'h6b == r_count_33_io_out ? io_r_107_b : _GEN_7006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7008 = 8'h6c == r_count_33_io_out ? io_r_108_b : _GEN_7007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7009 = 8'h6d == r_count_33_io_out ? io_r_109_b : _GEN_7008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7010 = 8'h6e == r_count_33_io_out ? io_r_110_b : _GEN_7009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7011 = 8'h6f == r_count_33_io_out ? io_r_111_b : _GEN_7010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7012 = 8'h70 == r_count_33_io_out ? io_r_112_b : _GEN_7011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7013 = 8'h71 == r_count_33_io_out ? io_r_113_b : _GEN_7012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7014 = 8'h72 == r_count_33_io_out ? io_r_114_b : _GEN_7013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7015 = 8'h73 == r_count_33_io_out ? io_r_115_b : _GEN_7014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7016 = 8'h74 == r_count_33_io_out ? io_r_116_b : _GEN_7015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7017 = 8'h75 == r_count_33_io_out ? io_r_117_b : _GEN_7016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7018 = 8'h76 == r_count_33_io_out ? io_r_118_b : _GEN_7017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7019 = 8'h77 == r_count_33_io_out ? io_r_119_b : _GEN_7018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7020 = 8'h78 == r_count_33_io_out ? io_r_120_b : _GEN_7019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7021 = 8'h79 == r_count_33_io_out ? io_r_121_b : _GEN_7020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7022 = 8'h7a == r_count_33_io_out ? io_r_122_b : _GEN_7021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7023 = 8'h7b == r_count_33_io_out ? io_r_123_b : _GEN_7022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7024 = 8'h7c == r_count_33_io_out ? io_r_124_b : _GEN_7023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7025 = 8'h7d == r_count_33_io_out ? io_r_125_b : _GEN_7024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7026 = 8'h7e == r_count_33_io_out ? io_r_126_b : _GEN_7025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7027 = 8'h7f == r_count_33_io_out ? io_r_127_b : _GEN_7026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7028 = 8'h80 == r_count_33_io_out ? io_r_128_b : _GEN_7027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7029 = 8'h81 == r_count_33_io_out ? io_r_129_b : _GEN_7028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7030 = 8'h82 == r_count_33_io_out ? io_r_130_b : _GEN_7029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7031 = 8'h83 == r_count_33_io_out ? io_r_131_b : _GEN_7030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7032 = 8'h84 == r_count_33_io_out ? io_r_132_b : _GEN_7031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7033 = 8'h85 == r_count_33_io_out ? io_r_133_b : _GEN_7032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7034 = 8'h86 == r_count_33_io_out ? io_r_134_b : _GEN_7033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7035 = 8'h87 == r_count_33_io_out ? io_r_135_b : _GEN_7034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7036 = 8'h88 == r_count_33_io_out ? io_r_136_b : _GEN_7035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7037 = 8'h89 == r_count_33_io_out ? io_r_137_b : _GEN_7036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7038 = 8'h8a == r_count_33_io_out ? io_r_138_b : _GEN_7037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7039 = 8'h8b == r_count_33_io_out ? io_r_139_b : _GEN_7038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7040 = 8'h8c == r_count_33_io_out ? io_r_140_b : _GEN_7039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7041 = 8'h8d == r_count_33_io_out ? io_r_141_b : _GEN_7040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7042 = 8'h8e == r_count_33_io_out ? io_r_142_b : _GEN_7041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7043 = 8'h8f == r_count_33_io_out ? io_r_143_b : _GEN_7042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7044 = 8'h90 == r_count_33_io_out ? io_r_144_b : _GEN_7043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7045 = 8'h91 == r_count_33_io_out ? io_r_145_b : _GEN_7044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7046 = 8'h92 == r_count_33_io_out ? io_r_146_b : _GEN_7045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7047 = 8'h93 == r_count_33_io_out ? io_r_147_b : _GEN_7046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7048 = 8'h94 == r_count_33_io_out ? io_r_148_b : _GEN_7047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7049 = 8'h95 == r_count_33_io_out ? io_r_149_b : _GEN_7048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7050 = 8'h96 == r_count_33_io_out ? io_r_150_b : _GEN_7049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7051 = 8'h97 == r_count_33_io_out ? io_r_151_b : _GEN_7050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7052 = 8'h98 == r_count_33_io_out ? io_r_152_b : _GEN_7051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7053 = 8'h99 == r_count_33_io_out ? io_r_153_b : _GEN_7052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7054 = 8'h9a == r_count_33_io_out ? io_r_154_b : _GEN_7053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7055 = 8'h9b == r_count_33_io_out ? io_r_155_b : _GEN_7054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7056 = 8'h9c == r_count_33_io_out ? io_r_156_b : _GEN_7055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7057 = 8'h9d == r_count_33_io_out ? io_r_157_b : _GEN_7056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7058 = 8'h9e == r_count_33_io_out ? io_r_158_b : _GEN_7057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7059 = 8'h9f == r_count_33_io_out ? io_r_159_b : _GEN_7058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7060 = 8'ha0 == r_count_33_io_out ? io_r_160_b : _GEN_7059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7061 = 8'ha1 == r_count_33_io_out ? io_r_161_b : _GEN_7060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7062 = 8'ha2 == r_count_33_io_out ? io_r_162_b : _GEN_7061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7063 = 8'ha3 == r_count_33_io_out ? io_r_163_b : _GEN_7062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7064 = 8'ha4 == r_count_33_io_out ? io_r_164_b : _GEN_7063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7065 = 8'ha5 == r_count_33_io_out ? io_r_165_b : _GEN_7064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7066 = 8'ha6 == r_count_33_io_out ? io_r_166_b : _GEN_7065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7067 = 8'ha7 == r_count_33_io_out ? io_r_167_b : _GEN_7066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7068 = 8'ha8 == r_count_33_io_out ? io_r_168_b : _GEN_7067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7069 = 8'ha9 == r_count_33_io_out ? io_r_169_b : _GEN_7068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7070 = 8'haa == r_count_33_io_out ? io_r_170_b : _GEN_7069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7071 = 8'hab == r_count_33_io_out ? io_r_171_b : _GEN_7070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7072 = 8'hac == r_count_33_io_out ? io_r_172_b : _GEN_7071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7073 = 8'had == r_count_33_io_out ? io_r_173_b : _GEN_7072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7074 = 8'hae == r_count_33_io_out ? io_r_174_b : _GEN_7073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7075 = 8'haf == r_count_33_io_out ? io_r_175_b : _GEN_7074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7076 = 8'hb0 == r_count_33_io_out ? io_r_176_b : _GEN_7075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7077 = 8'hb1 == r_count_33_io_out ? io_r_177_b : _GEN_7076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7078 = 8'hb2 == r_count_33_io_out ? io_r_178_b : _GEN_7077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7079 = 8'hb3 == r_count_33_io_out ? io_r_179_b : _GEN_7078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7080 = 8'hb4 == r_count_33_io_out ? io_r_180_b : _GEN_7079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7081 = 8'hb5 == r_count_33_io_out ? io_r_181_b : _GEN_7080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7082 = 8'hb6 == r_count_33_io_out ? io_r_182_b : _GEN_7081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7083 = 8'hb7 == r_count_33_io_out ? io_r_183_b : _GEN_7082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7084 = 8'hb8 == r_count_33_io_out ? io_r_184_b : _GEN_7083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7085 = 8'hb9 == r_count_33_io_out ? io_r_185_b : _GEN_7084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7086 = 8'hba == r_count_33_io_out ? io_r_186_b : _GEN_7085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7087 = 8'hbb == r_count_33_io_out ? io_r_187_b : _GEN_7086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7088 = 8'hbc == r_count_33_io_out ? io_r_188_b : _GEN_7087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7089 = 8'hbd == r_count_33_io_out ? io_r_189_b : _GEN_7088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7090 = 8'hbe == r_count_33_io_out ? io_r_190_b : _GEN_7089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7091 = 8'hbf == r_count_33_io_out ? io_r_191_b : _GEN_7090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7092 = 8'hc0 == r_count_33_io_out ? io_r_192_b : _GEN_7091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7093 = 8'hc1 == r_count_33_io_out ? io_r_193_b : _GEN_7092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7094 = 8'hc2 == r_count_33_io_out ? io_r_194_b : _GEN_7093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7095 = 8'hc3 == r_count_33_io_out ? io_r_195_b : _GEN_7094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7096 = 8'hc4 == r_count_33_io_out ? io_r_196_b : _GEN_7095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7097 = 8'hc5 == r_count_33_io_out ? io_r_197_b : _GEN_7096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7098 = 8'hc6 == r_count_33_io_out ? io_r_198_b : _GEN_7097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7101 = 8'h1 == r_count_34_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7102 = 8'h2 == r_count_34_io_out ? io_r_2_b : _GEN_7101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7103 = 8'h3 == r_count_34_io_out ? io_r_3_b : _GEN_7102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7104 = 8'h4 == r_count_34_io_out ? io_r_4_b : _GEN_7103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7105 = 8'h5 == r_count_34_io_out ? io_r_5_b : _GEN_7104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7106 = 8'h6 == r_count_34_io_out ? io_r_6_b : _GEN_7105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7107 = 8'h7 == r_count_34_io_out ? io_r_7_b : _GEN_7106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7108 = 8'h8 == r_count_34_io_out ? io_r_8_b : _GEN_7107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7109 = 8'h9 == r_count_34_io_out ? io_r_9_b : _GEN_7108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7110 = 8'ha == r_count_34_io_out ? io_r_10_b : _GEN_7109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7111 = 8'hb == r_count_34_io_out ? io_r_11_b : _GEN_7110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7112 = 8'hc == r_count_34_io_out ? io_r_12_b : _GEN_7111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7113 = 8'hd == r_count_34_io_out ? io_r_13_b : _GEN_7112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7114 = 8'he == r_count_34_io_out ? io_r_14_b : _GEN_7113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7115 = 8'hf == r_count_34_io_out ? io_r_15_b : _GEN_7114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7116 = 8'h10 == r_count_34_io_out ? io_r_16_b : _GEN_7115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7117 = 8'h11 == r_count_34_io_out ? io_r_17_b : _GEN_7116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7118 = 8'h12 == r_count_34_io_out ? io_r_18_b : _GEN_7117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7119 = 8'h13 == r_count_34_io_out ? io_r_19_b : _GEN_7118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7120 = 8'h14 == r_count_34_io_out ? io_r_20_b : _GEN_7119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7121 = 8'h15 == r_count_34_io_out ? io_r_21_b : _GEN_7120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7122 = 8'h16 == r_count_34_io_out ? io_r_22_b : _GEN_7121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7123 = 8'h17 == r_count_34_io_out ? io_r_23_b : _GEN_7122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7124 = 8'h18 == r_count_34_io_out ? io_r_24_b : _GEN_7123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7125 = 8'h19 == r_count_34_io_out ? io_r_25_b : _GEN_7124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7126 = 8'h1a == r_count_34_io_out ? io_r_26_b : _GEN_7125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7127 = 8'h1b == r_count_34_io_out ? io_r_27_b : _GEN_7126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7128 = 8'h1c == r_count_34_io_out ? io_r_28_b : _GEN_7127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7129 = 8'h1d == r_count_34_io_out ? io_r_29_b : _GEN_7128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7130 = 8'h1e == r_count_34_io_out ? io_r_30_b : _GEN_7129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7131 = 8'h1f == r_count_34_io_out ? io_r_31_b : _GEN_7130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7132 = 8'h20 == r_count_34_io_out ? io_r_32_b : _GEN_7131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7133 = 8'h21 == r_count_34_io_out ? io_r_33_b : _GEN_7132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7134 = 8'h22 == r_count_34_io_out ? io_r_34_b : _GEN_7133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7135 = 8'h23 == r_count_34_io_out ? io_r_35_b : _GEN_7134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7136 = 8'h24 == r_count_34_io_out ? io_r_36_b : _GEN_7135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7137 = 8'h25 == r_count_34_io_out ? io_r_37_b : _GEN_7136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7138 = 8'h26 == r_count_34_io_out ? io_r_38_b : _GEN_7137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7139 = 8'h27 == r_count_34_io_out ? io_r_39_b : _GEN_7138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7140 = 8'h28 == r_count_34_io_out ? io_r_40_b : _GEN_7139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7141 = 8'h29 == r_count_34_io_out ? io_r_41_b : _GEN_7140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7142 = 8'h2a == r_count_34_io_out ? io_r_42_b : _GEN_7141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7143 = 8'h2b == r_count_34_io_out ? io_r_43_b : _GEN_7142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7144 = 8'h2c == r_count_34_io_out ? io_r_44_b : _GEN_7143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7145 = 8'h2d == r_count_34_io_out ? io_r_45_b : _GEN_7144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7146 = 8'h2e == r_count_34_io_out ? io_r_46_b : _GEN_7145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7147 = 8'h2f == r_count_34_io_out ? io_r_47_b : _GEN_7146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7148 = 8'h30 == r_count_34_io_out ? io_r_48_b : _GEN_7147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7149 = 8'h31 == r_count_34_io_out ? io_r_49_b : _GEN_7148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7150 = 8'h32 == r_count_34_io_out ? io_r_50_b : _GEN_7149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7151 = 8'h33 == r_count_34_io_out ? io_r_51_b : _GEN_7150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7152 = 8'h34 == r_count_34_io_out ? io_r_52_b : _GEN_7151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7153 = 8'h35 == r_count_34_io_out ? io_r_53_b : _GEN_7152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7154 = 8'h36 == r_count_34_io_out ? io_r_54_b : _GEN_7153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7155 = 8'h37 == r_count_34_io_out ? io_r_55_b : _GEN_7154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7156 = 8'h38 == r_count_34_io_out ? io_r_56_b : _GEN_7155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7157 = 8'h39 == r_count_34_io_out ? io_r_57_b : _GEN_7156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7158 = 8'h3a == r_count_34_io_out ? io_r_58_b : _GEN_7157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7159 = 8'h3b == r_count_34_io_out ? io_r_59_b : _GEN_7158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7160 = 8'h3c == r_count_34_io_out ? io_r_60_b : _GEN_7159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7161 = 8'h3d == r_count_34_io_out ? io_r_61_b : _GEN_7160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7162 = 8'h3e == r_count_34_io_out ? io_r_62_b : _GEN_7161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7163 = 8'h3f == r_count_34_io_out ? io_r_63_b : _GEN_7162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7164 = 8'h40 == r_count_34_io_out ? io_r_64_b : _GEN_7163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7165 = 8'h41 == r_count_34_io_out ? io_r_65_b : _GEN_7164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7166 = 8'h42 == r_count_34_io_out ? io_r_66_b : _GEN_7165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7167 = 8'h43 == r_count_34_io_out ? io_r_67_b : _GEN_7166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7168 = 8'h44 == r_count_34_io_out ? io_r_68_b : _GEN_7167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7169 = 8'h45 == r_count_34_io_out ? io_r_69_b : _GEN_7168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7170 = 8'h46 == r_count_34_io_out ? io_r_70_b : _GEN_7169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7171 = 8'h47 == r_count_34_io_out ? io_r_71_b : _GEN_7170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7172 = 8'h48 == r_count_34_io_out ? io_r_72_b : _GEN_7171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7173 = 8'h49 == r_count_34_io_out ? io_r_73_b : _GEN_7172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7174 = 8'h4a == r_count_34_io_out ? io_r_74_b : _GEN_7173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7175 = 8'h4b == r_count_34_io_out ? io_r_75_b : _GEN_7174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7176 = 8'h4c == r_count_34_io_out ? io_r_76_b : _GEN_7175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7177 = 8'h4d == r_count_34_io_out ? io_r_77_b : _GEN_7176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7178 = 8'h4e == r_count_34_io_out ? io_r_78_b : _GEN_7177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7179 = 8'h4f == r_count_34_io_out ? io_r_79_b : _GEN_7178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7180 = 8'h50 == r_count_34_io_out ? io_r_80_b : _GEN_7179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7181 = 8'h51 == r_count_34_io_out ? io_r_81_b : _GEN_7180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7182 = 8'h52 == r_count_34_io_out ? io_r_82_b : _GEN_7181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7183 = 8'h53 == r_count_34_io_out ? io_r_83_b : _GEN_7182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7184 = 8'h54 == r_count_34_io_out ? io_r_84_b : _GEN_7183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7185 = 8'h55 == r_count_34_io_out ? io_r_85_b : _GEN_7184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7186 = 8'h56 == r_count_34_io_out ? io_r_86_b : _GEN_7185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7187 = 8'h57 == r_count_34_io_out ? io_r_87_b : _GEN_7186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7188 = 8'h58 == r_count_34_io_out ? io_r_88_b : _GEN_7187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7189 = 8'h59 == r_count_34_io_out ? io_r_89_b : _GEN_7188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7190 = 8'h5a == r_count_34_io_out ? io_r_90_b : _GEN_7189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7191 = 8'h5b == r_count_34_io_out ? io_r_91_b : _GEN_7190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7192 = 8'h5c == r_count_34_io_out ? io_r_92_b : _GEN_7191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7193 = 8'h5d == r_count_34_io_out ? io_r_93_b : _GEN_7192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7194 = 8'h5e == r_count_34_io_out ? io_r_94_b : _GEN_7193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7195 = 8'h5f == r_count_34_io_out ? io_r_95_b : _GEN_7194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7196 = 8'h60 == r_count_34_io_out ? io_r_96_b : _GEN_7195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7197 = 8'h61 == r_count_34_io_out ? io_r_97_b : _GEN_7196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7198 = 8'h62 == r_count_34_io_out ? io_r_98_b : _GEN_7197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7199 = 8'h63 == r_count_34_io_out ? io_r_99_b : _GEN_7198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7200 = 8'h64 == r_count_34_io_out ? io_r_100_b : _GEN_7199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7201 = 8'h65 == r_count_34_io_out ? io_r_101_b : _GEN_7200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7202 = 8'h66 == r_count_34_io_out ? io_r_102_b : _GEN_7201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7203 = 8'h67 == r_count_34_io_out ? io_r_103_b : _GEN_7202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7204 = 8'h68 == r_count_34_io_out ? io_r_104_b : _GEN_7203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7205 = 8'h69 == r_count_34_io_out ? io_r_105_b : _GEN_7204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7206 = 8'h6a == r_count_34_io_out ? io_r_106_b : _GEN_7205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7207 = 8'h6b == r_count_34_io_out ? io_r_107_b : _GEN_7206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7208 = 8'h6c == r_count_34_io_out ? io_r_108_b : _GEN_7207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7209 = 8'h6d == r_count_34_io_out ? io_r_109_b : _GEN_7208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7210 = 8'h6e == r_count_34_io_out ? io_r_110_b : _GEN_7209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7211 = 8'h6f == r_count_34_io_out ? io_r_111_b : _GEN_7210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7212 = 8'h70 == r_count_34_io_out ? io_r_112_b : _GEN_7211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7213 = 8'h71 == r_count_34_io_out ? io_r_113_b : _GEN_7212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7214 = 8'h72 == r_count_34_io_out ? io_r_114_b : _GEN_7213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7215 = 8'h73 == r_count_34_io_out ? io_r_115_b : _GEN_7214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7216 = 8'h74 == r_count_34_io_out ? io_r_116_b : _GEN_7215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7217 = 8'h75 == r_count_34_io_out ? io_r_117_b : _GEN_7216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7218 = 8'h76 == r_count_34_io_out ? io_r_118_b : _GEN_7217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7219 = 8'h77 == r_count_34_io_out ? io_r_119_b : _GEN_7218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7220 = 8'h78 == r_count_34_io_out ? io_r_120_b : _GEN_7219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7221 = 8'h79 == r_count_34_io_out ? io_r_121_b : _GEN_7220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7222 = 8'h7a == r_count_34_io_out ? io_r_122_b : _GEN_7221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7223 = 8'h7b == r_count_34_io_out ? io_r_123_b : _GEN_7222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7224 = 8'h7c == r_count_34_io_out ? io_r_124_b : _GEN_7223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7225 = 8'h7d == r_count_34_io_out ? io_r_125_b : _GEN_7224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7226 = 8'h7e == r_count_34_io_out ? io_r_126_b : _GEN_7225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7227 = 8'h7f == r_count_34_io_out ? io_r_127_b : _GEN_7226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7228 = 8'h80 == r_count_34_io_out ? io_r_128_b : _GEN_7227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7229 = 8'h81 == r_count_34_io_out ? io_r_129_b : _GEN_7228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7230 = 8'h82 == r_count_34_io_out ? io_r_130_b : _GEN_7229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7231 = 8'h83 == r_count_34_io_out ? io_r_131_b : _GEN_7230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7232 = 8'h84 == r_count_34_io_out ? io_r_132_b : _GEN_7231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7233 = 8'h85 == r_count_34_io_out ? io_r_133_b : _GEN_7232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7234 = 8'h86 == r_count_34_io_out ? io_r_134_b : _GEN_7233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7235 = 8'h87 == r_count_34_io_out ? io_r_135_b : _GEN_7234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7236 = 8'h88 == r_count_34_io_out ? io_r_136_b : _GEN_7235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7237 = 8'h89 == r_count_34_io_out ? io_r_137_b : _GEN_7236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7238 = 8'h8a == r_count_34_io_out ? io_r_138_b : _GEN_7237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7239 = 8'h8b == r_count_34_io_out ? io_r_139_b : _GEN_7238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7240 = 8'h8c == r_count_34_io_out ? io_r_140_b : _GEN_7239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7241 = 8'h8d == r_count_34_io_out ? io_r_141_b : _GEN_7240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7242 = 8'h8e == r_count_34_io_out ? io_r_142_b : _GEN_7241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7243 = 8'h8f == r_count_34_io_out ? io_r_143_b : _GEN_7242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7244 = 8'h90 == r_count_34_io_out ? io_r_144_b : _GEN_7243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7245 = 8'h91 == r_count_34_io_out ? io_r_145_b : _GEN_7244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7246 = 8'h92 == r_count_34_io_out ? io_r_146_b : _GEN_7245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7247 = 8'h93 == r_count_34_io_out ? io_r_147_b : _GEN_7246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7248 = 8'h94 == r_count_34_io_out ? io_r_148_b : _GEN_7247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7249 = 8'h95 == r_count_34_io_out ? io_r_149_b : _GEN_7248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7250 = 8'h96 == r_count_34_io_out ? io_r_150_b : _GEN_7249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7251 = 8'h97 == r_count_34_io_out ? io_r_151_b : _GEN_7250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7252 = 8'h98 == r_count_34_io_out ? io_r_152_b : _GEN_7251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7253 = 8'h99 == r_count_34_io_out ? io_r_153_b : _GEN_7252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7254 = 8'h9a == r_count_34_io_out ? io_r_154_b : _GEN_7253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7255 = 8'h9b == r_count_34_io_out ? io_r_155_b : _GEN_7254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7256 = 8'h9c == r_count_34_io_out ? io_r_156_b : _GEN_7255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7257 = 8'h9d == r_count_34_io_out ? io_r_157_b : _GEN_7256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7258 = 8'h9e == r_count_34_io_out ? io_r_158_b : _GEN_7257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7259 = 8'h9f == r_count_34_io_out ? io_r_159_b : _GEN_7258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7260 = 8'ha0 == r_count_34_io_out ? io_r_160_b : _GEN_7259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7261 = 8'ha1 == r_count_34_io_out ? io_r_161_b : _GEN_7260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7262 = 8'ha2 == r_count_34_io_out ? io_r_162_b : _GEN_7261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7263 = 8'ha3 == r_count_34_io_out ? io_r_163_b : _GEN_7262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7264 = 8'ha4 == r_count_34_io_out ? io_r_164_b : _GEN_7263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7265 = 8'ha5 == r_count_34_io_out ? io_r_165_b : _GEN_7264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7266 = 8'ha6 == r_count_34_io_out ? io_r_166_b : _GEN_7265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7267 = 8'ha7 == r_count_34_io_out ? io_r_167_b : _GEN_7266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7268 = 8'ha8 == r_count_34_io_out ? io_r_168_b : _GEN_7267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7269 = 8'ha9 == r_count_34_io_out ? io_r_169_b : _GEN_7268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7270 = 8'haa == r_count_34_io_out ? io_r_170_b : _GEN_7269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7271 = 8'hab == r_count_34_io_out ? io_r_171_b : _GEN_7270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7272 = 8'hac == r_count_34_io_out ? io_r_172_b : _GEN_7271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7273 = 8'had == r_count_34_io_out ? io_r_173_b : _GEN_7272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7274 = 8'hae == r_count_34_io_out ? io_r_174_b : _GEN_7273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7275 = 8'haf == r_count_34_io_out ? io_r_175_b : _GEN_7274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7276 = 8'hb0 == r_count_34_io_out ? io_r_176_b : _GEN_7275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7277 = 8'hb1 == r_count_34_io_out ? io_r_177_b : _GEN_7276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7278 = 8'hb2 == r_count_34_io_out ? io_r_178_b : _GEN_7277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7279 = 8'hb3 == r_count_34_io_out ? io_r_179_b : _GEN_7278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7280 = 8'hb4 == r_count_34_io_out ? io_r_180_b : _GEN_7279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7281 = 8'hb5 == r_count_34_io_out ? io_r_181_b : _GEN_7280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7282 = 8'hb6 == r_count_34_io_out ? io_r_182_b : _GEN_7281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7283 = 8'hb7 == r_count_34_io_out ? io_r_183_b : _GEN_7282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7284 = 8'hb8 == r_count_34_io_out ? io_r_184_b : _GEN_7283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7285 = 8'hb9 == r_count_34_io_out ? io_r_185_b : _GEN_7284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7286 = 8'hba == r_count_34_io_out ? io_r_186_b : _GEN_7285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7287 = 8'hbb == r_count_34_io_out ? io_r_187_b : _GEN_7286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7288 = 8'hbc == r_count_34_io_out ? io_r_188_b : _GEN_7287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7289 = 8'hbd == r_count_34_io_out ? io_r_189_b : _GEN_7288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7290 = 8'hbe == r_count_34_io_out ? io_r_190_b : _GEN_7289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7291 = 8'hbf == r_count_34_io_out ? io_r_191_b : _GEN_7290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7292 = 8'hc0 == r_count_34_io_out ? io_r_192_b : _GEN_7291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7293 = 8'hc1 == r_count_34_io_out ? io_r_193_b : _GEN_7292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7294 = 8'hc2 == r_count_34_io_out ? io_r_194_b : _GEN_7293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7295 = 8'hc3 == r_count_34_io_out ? io_r_195_b : _GEN_7294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7296 = 8'hc4 == r_count_34_io_out ? io_r_196_b : _GEN_7295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7297 = 8'hc5 == r_count_34_io_out ? io_r_197_b : _GEN_7296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7298 = 8'hc6 == r_count_34_io_out ? io_r_198_b : _GEN_7297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7301 = 8'h1 == r_count_35_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7302 = 8'h2 == r_count_35_io_out ? io_r_2_b : _GEN_7301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7303 = 8'h3 == r_count_35_io_out ? io_r_3_b : _GEN_7302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7304 = 8'h4 == r_count_35_io_out ? io_r_4_b : _GEN_7303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7305 = 8'h5 == r_count_35_io_out ? io_r_5_b : _GEN_7304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7306 = 8'h6 == r_count_35_io_out ? io_r_6_b : _GEN_7305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7307 = 8'h7 == r_count_35_io_out ? io_r_7_b : _GEN_7306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7308 = 8'h8 == r_count_35_io_out ? io_r_8_b : _GEN_7307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7309 = 8'h9 == r_count_35_io_out ? io_r_9_b : _GEN_7308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7310 = 8'ha == r_count_35_io_out ? io_r_10_b : _GEN_7309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7311 = 8'hb == r_count_35_io_out ? io_r_11_b : _GEN_7310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7312 = 8'hc == r_count_35_io_out ? io_r_12_b : _GEN_7311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7313 = 8'hd == r_count_35_io_out ? io_r_13_b : _GEN_7312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7314 = 8'he == r_count_35_io_out ? io_r_14_b : _GEN_7313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7315 = 8'hf == r_count_35_io_out ? io_r_15_b : _GEN_7314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7316 = 8'h10 == r_count_35_io_out ? io_r_16_b : _GEN_7315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7317 = 8'h11 == r_count_35_io_out ? io_r_17_b : _GEN_7316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7318 = 8'h12 == r_count_35_io_out ? io_r_18_b : _GEN_7317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7319 = 8'h13 == r_count_35_io_out ? io_r_19_b : _GEN_7318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7320 = 8'h14 == r_count_35_io_out ? io_r_20_b : _GEN_7319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7321 = 8'h15 == r_count_35_io_out ? io_r_21_b : _GEN_7320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7322 = 8'h16 == r_count_35_io_out ? io_r_22_b : _GEN_7321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7323 = 8'h17 == r_count_35_io_out ? io_r_23_b : _GEN_7322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7324 = 8'h18 == r_count_35_io_out ? io_r_24_b : _GEN_7323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7325 = 8'h19 == r_count_35_io_out ? io_r_25_b : _GEN_7324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7326 = 8'h1a == r_count_35_io_out ? io_r_26_b : _GEN_7325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7327 = 8'h1b == r_count_35_io_out ? io_r_27_b : _GEN_7326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7328 = 8'h1c == r_count_35_io_out ? io_r_28_b : _GEN_7327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7329 = 8'h1d == r_count_35_io_out ? io_r_29_b : _GEN_7328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7330 = 8'h1e == r_count_35_io_out ? io_r_30_b : _GEN_7329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7331 = 8'h1f == r_count_35_io_out ? io_r_31_b : _GEN_7330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7332 = 8'h20 == r_count_35_io_out ? io_r_32_b : _GEN_7331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7333 = 8'h21 == r_count_35_io_out ? io_r_33_b : _GEN_7332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7334 = 8'h22 == r_count_35_io_out ? io_r_34_b : _GEN_7333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7335 = 8'h23 == r_count_35_io_out ? io_r_35_b : _GEN_7334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7336 = 8'h24 == r_count_35_io_out ? io_r_36_b : _GEN_7335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7337 = 8'h25 == r_count_35_io_out ? io_r_37_b : _GEN_7336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7338 = 8'h26 == r_count_35_io_out ? io_r_38_b : _GEN_7337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7339 = 8'h27 == r_count_35_io_out ? io_r_39_b : _GEN_7338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7340 = 8'h28 == r_count_35_io_out ? io_r_40_b : _GEN_7339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7341 = 8'h29 == r_count_35_io_out ? io_r_41_b : _GEN_7340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7342 = 8'h2a == r_count_35_io_out ? io_r_42_b : _GEN_7341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7343 = 8'h2b == r_count_35_io_out ? io_r_43_b : _GEN_7342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7344 = 8'h2c == r_count_35_io_out ? io_r_44_b : _GEN_7343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7345 = 8'h2d == r_count_35_io_out ? io_r_45_b : _GEN_7344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7346 = 8'h2e == r_count_35_io_out ? io_r_46_b : _GEN_7345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7347 = 8'h2f == r_count_35_io_out ? io_r_47_b : _GEN_7346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7348 = 8'h30 == r_count_35_io_out ? io_r_48_b : _GEN_7347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7349 = 8'h31 == r_count_35_io_out ? io_r_49_b : _GEN_7348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7350 = 8'h32 == r_count_35_io_out ? io_r_50_b : _GEN_7349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7351 = 8'h33 == r_count_35_io_out ? io_r_51_b : _GEN_7350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7352 = 8'h34 == r_count_35_io_out ? io_r_52_b : _GEN_7351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7353 = 8'h35 == r_count_35_io_out ? io_r_53_b : _GEN_7352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7354 = 8'h36 == r_count_35_io_out ? io_r_54_b : _GEN_7353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7355 = 8'h37 == r_count_35_io_out ? io_r_55_b : _GEN_7354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7356 = 8'h38 == r_count_35_io_out ? io_r_56_b : _GEN_7355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7357 = 8'h39 == r_count_35_io_out ? io_r_57_b : _GEN_7356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7358 = 8'h3a == r_count_35_io_out ? io_r_58_b : _GEN_7357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7359 = 8'h3b == r_count_35_io_out ? io_r_59_b : _GEN_7358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7360 = 8'h3c == r_count_35_io_out ? io_r_60_b : _GEN_7359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7361 = 8'h3d == r_count_35_io_out ? io_r_61_b : _GEN_7360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7362 = 8'h3e == r_count_35_io_out ? io_r_62_b : _GEN_7361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7363 = 8'h3f == r_count_35_io_out ? io_r_63_b : _GEN_7362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7364 = 8'h40 == r_count_35_io_out ? io_r_64_b : _GEN_7363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7365 = 8'h41 == r_count_35_io_out ? io_r_65_b : _GEN_7364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7366 = 8'h42 == r_count_35_io_out ? io_r_66_b : _GEN_7365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7367 = 8'h43 == r_count_35_io_out ? io_r_67_b : _GEN_7366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7368 = 8'h44 == r_count_35_io_out ? io_r_68_b : _GEN_7367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7369 = 8'h45 == r_count_35_io_out ? io_r_69_b : _GEN_7368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7370 = 8'h46 == r_count_35_io_out ? io_r_70_b : _GEN_7369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7371 = 8'h47 == r_count_35_io_out ? io_r_71_b : _GEN_7370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7372 = 8'h48 == r_count_35_io_out ? io_r_72_b : _GEN_7371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7373 = 8'h49 == r_count_35_io_out ? io_r_73_b : _GEN_7372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7374 = 8'h4a == r_count_35_io_out ? io_r_74_b : _GEN_7373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7375 = 8'h4b == r_count_35_io_out ? io_r_75_b : _GEN_7374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7376 = 8'h4c == r_count_35_io_out ? io_r_76_b : _GEN_7375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7377 = 8'h4d == r_count_35_io_out ? io_r_77_b : _GEN_7376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7378 = 8'h4e == r_count_35_io_out ? io_r_78_b : _GEN_7377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7379 = 8'h4f == r_count_35_io_out ? io_r_79_b : _GEN_7378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7380 = 8'h50 == r_count_35_io_out ? io_r_80_b : _GEN_7379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7381 = 8'h51 == r_count_35_io_out ? io_r_81_b : _GEN_7380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7382 = 8'h52 == r_count_35_io_out ? io_r_82_b : _GEN_7381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7383 = 8'h53 == r_count_35_io_out ? io_r_83_b : _GEN_7382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7384 = 8'h54 == r_count_35_io_out ? io_r_84_b : _GEN_7383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7385 = 8'h55 == r_count_35_io_out ? io_r_85_b : _GEN_7384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7386 = 8'h56 == r_count_35_io_out ? io_r_86_b : _GEN_7385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7387 = 8'h57 == r_count_35_io_out ? io_r_87_b : _GEN_7386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7388 = 8'h58 == r_count_35_io_out ? io_r_88_b : _GEN_7387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7389 = 8'h59 == r_count_35_io_out ? io_r_89_b : _GEN_7388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7390 = 8'h5a == r_count_35_io_out ? io_r_90_b : _GEN_7389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7391 = 8'h5b == r_count_35_io_out ? io_r_91_b : _GEN_7390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7392 = 8'h5c == r_count_35_io_out ? io_r_92_b : _GEN_7391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7393 = 8'h5d == r_count_35_io_out ? io_r_93_b : _GEN_7392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7394 = 8'h5e == r_count_35_io_out ? io_r_94_b : _GEN_7393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7395 = 8'h5f == r_count_35_io_out ? io_r_95_b : _GEN_7394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7396 = 8'h60 == r_count_35_io_out ? io_r_96_b : _GEN_7395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7397 = 8'h61 == r_count_35_io_out ? io_r_97_b : _GEN_7396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7398 = 8'h62 == r_count_35_io_out ? io_r_98_b : _GEN_7397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7399 = 8'h63 == r_count_35_io_out ? io_r_99_b : _GEN_7398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7400 = 8'h64 == r_count_35_io_out ? io_r_100_b : _GEN_7399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7401 = 8'h65 == r_count_35_io_out ? io_r_101_b : _GEN_7400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7402 = 8'h66 == r_count_35_io_out ? io_r_102_b : _GEN_7401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7403 = 8'h67 == r_count_35_io_out ? io_r_103_b : _GEN_7402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7404 = 8'h68 == r_count_35_io_out ? io_r_104_b : _GEN_7403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7405 = 8'h69 == r_count_35_io_out ? io_r_105_b : _GEN_7404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7406 = 8'h6a == r_count_35_io_out ? io_r_106_b : _GEN_7405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7407 = 8'h6b == r_count_35_io_out ? io_r_107_b : _GEN_7406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7408 = 8'h6c == r_count_35_io_out ? io_r_108_b : _GEN_7407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7409 = 8'h6d == r_count_35_io_out ? io_r_109_b : _GEN_7408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7410 = 8'h6e == r_count_35_io_out ? io_r_110_b : _GEN_7409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7411 = 8'h6f == r_count_35_io_out ? io_r_111_b : _GEN_7410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7412 = 8'h70 == r_count_35_io_out ? io_r_112_b : _GEN_7411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7413 = 8'h71 == r_count_35_io_out ? io_r_113_b : _GEN_7412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7414 = 8'h72 == r_count_35_io_out ? io_r_114_b : _GEN_7413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7415 = 8'h73 == r_count_35_io_out ? io_r_115_b : _GEN_7414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7416 = 8'h74 == r_count_35_io_out ? io_r_116_b : _GEN_7415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7417 = 8'h75 == r_count_35_io_out ? io_r_117_b : _GEN_7416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7418 = 8'h76 == r_count_35_io_out ? io_r_118_b : _GEN_7417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7419 = 8'h77 == r_count_35_io_out ? io_r_119_b : _GEN_7418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7420 = 8'h78 == r_count_35_io_out ? io_r_120_b : _GEN_7419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7421 = 8'h79 == r_count_35_io_out ? io_r_121_b : _GEN_7420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7422 = 8'h7a == r_count_35_io_out ? io_r_122_b : _GEN_7421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7423 = 8'h7b == r_count_35_io_out ? io_r_123_b : _GEN_7422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7424 = 8'h7c == r_count_35_io_out ? io_r_124_b : _GEN_7423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7425 = 8'h7d == r_count_35_io_out ? io_r_125_b : _GEN_7424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7426 = 8'h7e == r_count_35_io_out ? io_r_126_b : _GEN_7425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7427 = 8'h7f == r_count_35_io_out ? io_r_127_b : _GEN_7426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7428 = 8'h80 == r_count_35_io_out ? io_r_128_b : _GEN_7427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7429 = 8'h81 == r_count_35_io_out ? io_r_129_b : _GEN_7428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7430 = 8'h82 == r_count_35_io_out ? io_r_130_b : _GEN_7429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7431 = 8'h83 == r_count_35_io_out ? io_r_131_b : _GEN_7430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7432 = 8'h84 == r_count_35_io_out ? io_r_132_b : _GEN_7431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7433 = 8'h85 == r_count_35_io_out ? io_r_133_b : _GEN_7432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7434 = 8'h86 == r_count_35_io_out ? io_r_134_b : _GEN_7433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7435 = 8'h87 == r_count_35_io_out ? io_r_135_b : _GEN_7434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7436 = 8'h88 == r_count_35_io_out ? io_r_136_b : _GEN_7435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7437 = 8'h89 == r_count_35_io_out ? io_r_137_b : _GEN_7436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7438 = 8'h8a == r_count_35_io_out ? io_r_138_b : _GEN_7437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7439 = 8'h8b == r_count_35_io_out ? io_r_139_b : _GEN_7438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7440 = 8'h8c == r_count_35_io_out ? io_r_140_b : _GEN_7439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7441 = 8'h8d == r_count_35_io_out ? io_r_141_b : _GEN_7440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7442 = 8'h8e == r_count_35_io_out ? io_r_142_b : _GEN_7441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7443 = 8'h8f == r_count_35_io_out ? io_r_143_b : _GEN_7442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7444 = 8'h90 == r_count_35_io_out ? io_r_144_b : _GEN_7443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7445 = 8'h91 == r_count_35_io_out ? io_r_145_b : _GEN_7444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7446 = 8'h92 == r_count_35_io_out ? io_r_146_b : _GEN_7445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7447 = 8'h93 == r_count_35_io_out ? io_r_147_b : _GEN_7446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7448 = 8'h94 == r_count_35_io_out ? io_r_148_b : _GEN_7447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7449 = 8'h95 == r_count_35_io_out ? io_r_149_b : _GEN_7448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7450 = 8'h96 == r_count_35_io_out ? io_r_150_b : _GEN_7449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7451 = 8'h97 == r_count_35_io_out ? io_r_151_b : _GEN_7450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7452 = 8'h98 == r_count_35_io_out ? io_r_152_b : _GEN_7451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7453 = 8'h99 == r_count_35_io_out ? io_r_153_b : _GEN_7452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7454 = 8'h9a == r_count_35_io_out ? io_r_154_b : _GEN_7453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7455 = 8'h9b == r_count_35_io_out ? io_r_155_b : _GEN_7454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7456 = 8'h9c == r_count_35_io_out ? io_r_156_b : _GEN_7455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7457 = 8'h9d == r_count_35_io_out ? io_r_157_b : _GEN_7456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7458 = 8'h9e == r_count_35_io_out ? io_r_158_b : _GEN_7457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7459 = 8'h9f == r_count_35_io_out ? io_r_159_b : _GEN_7458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7460 = 8'ha0 == r_count_35_io_out ? io_r_160_b : _GEN_7459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7461 = 8'ha1 == r_count_35_io_out ? io_r_161_b : _GEN_7460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7462 = 8'ha2 == r_count_35_io_out ? io_r_162_b : _GEN_7461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7463 = 8'ha3 == r_count_35_io_out ? io_r_163_b : _GEN_7462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7464 = 8'ha4 == r_count_35_io_out ? io_r_164_b : _GEN_7463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7465 = 8'ha5 == r_count_35_io_out ? io_r_165_b : _GEN_7464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7466 = 8'ha6 == r_count_35_io_out ? io_r_166_b : _GEN_7465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7467 = 8'ha7 == r_count_35_io_out ? io_r_167_b : _GEN_7466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7468 = 8'ha8 == r_count_35_io_out ? io_r_168_b : _GEN_7467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7469 = 8'ha9 == r_count_35_io_out ? io_r_169_b : _GEN_7468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7470 = 8'haa == r_count_35_io_out ? io_r_170_b : _GEN_7469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7471 = 8'hab == r_count_35_io_out ? io_r_171_b : _GEN_7470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7472 = 8'hac == r_count_35_io_out ? io_r_172_b : _GEN_7471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7473 = 8'had == r_count_35_io_out ? io_r_173_b : _GEN_7472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7474 = 8'hae == r_count_35_io_out ? io_r_174_b : _GEN_7473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7475 = 8'haf == r_count_35_io_out ? io_r_175_b : _GEN_7474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7476 = 8'hb0 == r_count_35_io_out ? io_r_176_b : _GEN_7475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7477 = 8'hb1 == r_count_35_io_out ? io_r_177_b : _GEN_7476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7478 = 8'hb2 == r_count_35_io_out ? io_r_178_b : _GEN_7477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7479 = 8'hb3 == r_count_35_io_out ? io_r_179_b : _GEN_7478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7480 = 8'hb4 == r_count_35_io_out ? io_r_180_b : _GEN_7479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7481 = 8'hb5 == r_count_35_io_out ? io_r_181_b : _GEN_7480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7482 = 8'hb6 == r_count_35_io_out ? io_r_182_b : _GEN_7481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7483 = 8'hb7 == r_count_35_io_out ? io_r_183_b : _GEN_7482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7484 = 8'hb8 == r_count_35_io_out ? io_r_184_b : _GEN_7483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7485 = 8'hb9 == r_count_35_io_out ? io_r_185_b : _GEN_7484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7486 = 8'hba == r_count_35_io_out ? io_r_186_b : _GEN_7485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7487 = 8'hbb == r_count_35_io_out ? io_r_187_b : _GEN_7486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7488 = 8'hbc == r_count_35_io_out ? io_r_188_b : _GEN_7487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7489 = 8'hbd == r_count_35_io_out ? io_r_189_b : _GEN_7488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7490 = 8'hbe == r_count_35_io_out ? io_r_190_b : _GEN_7489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7491 = 8'hbf == r_count_35_io_out ? io_r_191_b : _GEN_7490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7492 = 8'hc0 == r_count_35_io_out ? io_r_192_b : _GEN_7491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7493 = 8'hc1 == r_count_35_io_out ? io_r_193_b : _GEN_7492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7494 = 8'hc2 == r_count_35_io_out ? io_r_194_b : _GEN_7493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7495 = 8'hc3 == r_count_35_io_out ? io_r_195_b : _GEN_7494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7496 = 8'hc4 == r_count_35_io_out ? io_r_196_b : _GEN_7495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7497 = 8'hc5 == r_count_35_io_out ? io_r_197_b : _GEN_7496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7498 = 8'hc6 == r_count_35_io_out ? io_r_198_b : _GEN_7497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7501 = 8'h1 == r_count_36_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7502 = 8'h2 == r_count_36_io_out ? io_r_2_b : _GEN_7501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7503 = 8'h3 == r_count_36_io_out ? io_r_3_b : _GEN_7502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7504 = 8'h4 == r_count_36_io_out ? io_r_4_b : _GEN_7503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7505 = 8'h5 == r_count_36_io_out ? io_r_5_b : _GEN_7504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7506 = 8'h6 == r_count_36_io_out ? io_r_6_b : _GEN_7505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7507 = 8'h7 == r_count_36_io_out ? io_r_7_b : _GEN_7506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7508 = 8'h8 == r_count_36_io_out ? io_r_8_b : _GEN_7507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7509 = 8'h9 == r_count_36_io_out ? io_r_9_b : _GEN_7508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7510 = 8'ha == r_count_36_io_out ? io_r_10_b : _GEN_7509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7511 = 8'hb == r_count_36_io_out ? io_r_11_b : _GEN_7510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7512 = 8'hc == r_count_36_io_out ? io_r_12_b : _GEN_7511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7513 = 8'hd == r_count_36_io_out ? io_r_13_b : _GEN_7512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7514 = 8'he == r_count_36_io_out ? io_r_14_b : _GEN_7513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7515 = 8'hf == r_count_36_io_out ? io_r_15_b : _GEN_7514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7516 = 8'h10 == r_count_36_io_out ? io_r_16_b : _GEN_7515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7517 = 8'h11 == r_count_36_io_out ? io_r_17_b : _GEN_7516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7518 = 8'h12 == r_count_36_io_out ? io_r_18_b : _GEN_7517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7519 = 8'h13 == r_count_36_io_out ? io_r_19_b : _GEN_7518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7520 = 8'h14 == r_count_36_io_out ? io_r_20_b : _GEN_7519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7521 = 8'h15 == r_count_36_io_out ? io_r_21_b : _GEN_7520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7522 = 8'h16 == r_count_36_io_out ? io_r_22_b : _GEN_7521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7523 = 8'h17 == r_count_36_io_out ? io_r_23_b : _GEN_7522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7524 = 8'h18 == r_count_36_io_out ? io_r_24_b : _GEN_7523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7525 = 8'h19 == r_count_36_io_out ? io_r_25_b : _GEN_7524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7526 = 8'h1a == r_count_36_io_out ? io_r_26_b : _GEN_7525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7527 = 8'h1b == r_count_36_io_out ? io_r_27_b : _GEN_7526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7528 = 8'h1c == r_count_36_io_out ? io_r_28_b : _GEN_7527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7529 = 8'h1d == r_count_36_io_out ? io_r_29_b : _GEN_7528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7530 = 8'h1e == r_count_36_io_out ? io_r_30_b : _GEN_7529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7531 = 8'h1f == r_count_36_io_out ? io_r_31_b : _GEN_7530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7532 = 8'h20 == r_count_36_io_out ? io_r_32_b : _GEN_7531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7533 = 8'h21 == r_count_36_io_out ? io_r_33_b : _GEN_7532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7534 = 8'h22 == r_count_36_io_out ? io_r_34_b : _GEN_7533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7535 = 8'h23 == r_count_36_io_out ? io_r_35_b : _GEN_7534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7536 = 8'h24 == r_count_36_io_out ? io_r_36_b : _GEN_7535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7537 = 8'h25 == r_count_36_io_out ? io_r_37_b : _GEN_7536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7538 = 8'h26 == r_count_36_io_out ? io_r_38_b : _GEN_7537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7539 = 8'h27 == r_count_36_io_out ? io_r_39_b : _GEN_7538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7540 = 8'h28 == r_count_36_io_out ? io_r_40_b : _GEN_7539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7541 = 8'h29 == r_count_36_io_out ? io_r_41_b : _GEN_7540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7542 = 8'h2a == r_count_36_io_out ? io_r_42_b : _GEN_7541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7543 = 8'h2b == r_count_36_io_out ? io_r_43_b : _GEN_7542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7544 = 8'h2c == r_count_36_io_out ? io_r_44_b : _GEN_7543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7545 = 8'h2d == r_count_36_io_out ? io_r_45_b : _GEN_7544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7546 = 8'h2e == r_count_36_io_out ? io_r_46_b : _GEN_7545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7547 = 8'h2f == r_count_36_io_out ? io_r_47_b : _GEN_7546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7548 = 8'h30 == r_count_36_io_out ? io_r_48_b : _GEN_7547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7549 = 8'h31 == r_count_36_io_out ? io_r_49_b : _GEN_7548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7550 = 8'h32 == r_count_36_io_out ? io_r_50_b : _GEN_7549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7551 = 8'h33 == r_count_36_io_out ? io_r_51_b : _GEN_7550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7552 = 8'h34 == r_count_36_io_out ? io_r_52_b : _GEN_7551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7553 = 8'h35 == r_count_36_io_out ? io_r_53_b : _GEN_7552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7554 = 8'h36 == r_count_36_io_out ? io_r_54_b : _GEN_7553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7555 = 8'h37 == r_count_36_io_out ? io_r_55_b : _GEN_7554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7556 = 8'h38 == r_count_36_io_out ? io_r_56_b : _GEN_7555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7557 = 8'h39 == r_count_36_io_out ? io_r_57_b : _GEN_7556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7558 = 8'h3a == r_count_36_io_out ? io_r_58_b : _GEN_7557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7559 = 8'h3b == r_count_36_io_out ? io_r_59_b : _GEN_7558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7560 = 8'h3c == r_count_36_io_out ? io_r_60_b : _GEN_7559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7561 = 8'h3d == r_count_36_io_out ? io_r_61_b : _GEN_7560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7562 = 8'h3e == r_count_36_io_out ? io_r_62_b : _GEN_7561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7563 = 8'h3f == r_count_36_io_out ? io_r_63_b : _GEN_7562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7564 = 8'h40 == r_count_36_io_out ? io_r_64_b : _GEN_7563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7565 = 8'h41 == r_count_36_io_out ? io_r_65_b : _GEN_7564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7566 = 8'h42 == r_count_36_io_out ? io_r_66_b : _GEN_7565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7567 = 8'h43 == r_count_36_io_out ? io_r_67_b : _GEN_7566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7568 = 8'h44 == r_count_36_io_out ? io_r_68_b : _GEN_7567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7569 = 8'h45 == r_count_36_io_out ? io_r_69_b : _GEN_7568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7570 = 8'h46 == r_count_36_io_out ? io_r_70_b : _GEN_7569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7571 = 8'h47 == r_count_36_io_out ? io_r_71_b : _GEN_7570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7572 = 8'h48 == r_count_36_io_out ? io_r_72_b : _GEN_7571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7573 = 8'h49 == r_count_36_io_out ? io_r_73_b : _GEN_7572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7574 = 8'h4a == r_count_36_io_out ? io_r_74_b : _GEN_7573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7575 = 8'h4b == r_count_36_io_out ? io_r_75_b : _GEN_7574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7576 = 8'h4c == r_count_36_io_out ? io_r_76_b : _GEN_7575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7577 = 8'h4d == r_count_36_io_out ? io_r_77_b : _GEN_7576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7578 = 8'h4e == r_count_36_io_out ? io_r_78_b : _GEN_7577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7579 = 8'h4f == r_count_36_io_out ? io_r_79_b : _GEN_7578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7580 = 8'h50 == r_count_36_io_out ? io_r_80_b : _GEN_7579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7581 = 8'h51 == r_count_36_io_out ? io_r_81_b : _GEN_7580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7582 = 8'h52 == r_count_36_io_out ? io_r_82_b : _GEN_7581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7583 = 8'h53 == r_count_36_io_out ? io_r_83_b : _GEN_7582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7584 = 8'h54 == r_count_36_io_out ? io_r_84_b : _GEN_7583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7585 = 8'h55 == r_count_36_io_out ? io_r_85_b : _GEN_7584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7586 = 8'h56 == r_count_36_io_out ? io_r_86_b : _GEN_7585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7587 = 8'h57 == r_count_36_io_out ? io_r_87_b : _GEN_7586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7588 = 8'h58 == r_count_36_io_out ? io_r_88_b : _GEN_7587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7589 = 8'h59 == r_count_36_io_out ? io_r_89_b : _GEN_7588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7590 = 8'h5a == r_count_36_io_out ? io_r_90_b : _GEN_7589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7591 = 8'h5b == r_count_36_io_out ? io_r_91_b : _GEN_7590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7592 = 8'h5c == r_count_36_io_out ? io_r_92_b : _GEN_7591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7593 = 8'h5d == r_count_36_io_out ? io_r_93_b : _GEN_7592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7594 = 8'h5e == r_count_36_io_out ? io_r_94_b : _GEN_7593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7595 = 8'h5f == r_count_36_io_out ? io_r_95_b : _GEN_7594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7596 = 8'h60 == r_count_36_io_out ? io_r_96_b : _GEN_7595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7597 = 8'h61 == r_count_36_io_out ? io_r_97_b : _GEN_7596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7598 = 8'h62 == r_count_36_io_out ? io_r_98_b : _GEN_7597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7599 = 8'h63 == r_count_36_io_out ? io_r_99_b : _GEN_7598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7600 = 8'h64 == r_count_36_io_out ? io_r_100_b : _GEN_7599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7601 = 8'h65 == r_count_36_io_out ? io_r_101_b : _GEN_7600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7602 = 8'h66 == r_count_36_io_out ? io_r_102_b : _GEN_7601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7603 = 8'h67 == r_count_36_io_out ? io_r_103_b : _GEN_7602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7604 = 8'h68 == r_count_36_io_out ? io_r_104_b : _GEN_7603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7605 = 8'h69 == r_count_36_io_out ? io_r_105_b : _GEN_7604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7606 = 8'h6a == r_count_36_io_out ? io_r_106_b : _GEN_7605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7607 = 8'h6b == r_count_36_io_out ? io_r_107_b : _GEN_7606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7608 = 8'h6c == r_count_36_io_out ? io_r_108_b : _GEN_7607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7609 = 8'h6d == r_count_36_io_out ? io_r_109_b : _GEN_7608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7610 = 8'h6e == r_count_36_io_out ? io_r_110_b : _GEN_7609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7611 = 8'h6f == r_count_36_io_out ? io_r_111_b : _GEN_7610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7612 = 8'h70 == r_count_36_io_out ? io_r_112_b : _GEN_7611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7613 = 8'h71 == r_count_36_io_out ? io_r_113_b : _GEN_7612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7614 = 8'h72 == r_count_36_io_out ? io_r_114_b : _GEN_7613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7615 = 8'h73 == r_count_36_io_out ? io_r_115_b : _GEN_7614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7616 = 8'h74 == r_count_36_io_out ? io_r_116_b : _GEN_7615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7617 = 8'h75 == r_count_36_io_out ? io_r_117_b : _GEN_7616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7618 = 8'h76 == r_count_36_io_out ? io_r_118_b : _GEN_7617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7619 = 8'h77 == r_count_36_io_out ? io_r_119_b : _GEN_7618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7620 = 8'h78 == r_count_36_io_out ? io_r_120_b : _GEN_7619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7621 = 8'h79 == r_count_36_io_out ? io_r_121_b : _GEN_7620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7622 = 8'h7a == r_count_36_io_out ? io_r_122_b : _GEN_7621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7623 = 8'h7b == r_count_36_io_out ? io_r_123_b : _GEN_7622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7624 = 8'h7c == r_count_36_io_out ? io_r_124_b : _GEN_7623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7625 = 8'h7d == r_count_36_io_out ? io_r_125_b : _GEN_7624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7626 = 8'h7e == r_count_36_io_out ? io_r_126_b : _GEN_7625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7627 = 8'h7f == r_count_36_io_out ? io_r_127_b : _GEN_7626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7628 = 8'h80 == r_count_36_io_out ? io_r_128_b : _GEN_7627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7629 = 8'h81 == r_count_36_io_out ? io_r_129_b : _GEN_7628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7630 = 8'h82 == r_count_36_io_out ? io_r_130_b : _GEN_7629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7631 = 8'h83 == r_count_36_io_out ? io_r_131_b : _GEN_7630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7632 = 8'h84 == r_count_36_io_out ? io_r_132_b : _GEN_7631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7633 = 8'h85 == r_count_36_io_out ? io_r_133_b : _GEN_7632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7634 = 8'h86 == r_count_36_io_out ? io_r_134_b : _GEN_7633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7635 = 8'h87 == r_count_36_io_out ? io_r_135_b : _GEN_7634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7636 = 8'h88 == r_count_36_io_out ? io_r_136_b : _GEN_7635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7637 = 8'h89 == r_count_36_io_out ? io_r_137_b : _GEN_7636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7638 = 8'h8a == r_count_36_io_out ? io_r_138_b : _GEN_7637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7639 = 8'h8b == r_count_36_io_out ? io_r_139_b : _GEN_7638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7640 = 8'h8c == r_count_36_io_out ? io_r_140_b : _GEN_7639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7641 = 8'h8d == r_count_36_io_out ? io_r_141_b : _GEN_7640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7642 = 8'h8e == r_count_36_io_out ? io_r_142_b : _GEN_7641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7643 = 8'h8f == r_count_36_io_out ? io_r_143_b : _GEN_7642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7644 = 8'h90 == r_count_36_io_out ? io_r_144_b : _GEN_7643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7645 = 8'h91 == r_count_36_io_out ? io_r_145_b : _GEN_7644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7646 = 8'h92 == r_count_36_io_out ? io_r_146_b : _GEN_7645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7647 = 8'h93 == r_count_36_io_out ? io_r_147_b : _GEN_7646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7648 = 8'h94 == r_count_36_io_out ? io_r_148_b : _GEN_7647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7649 = 8'h95 == r_count_36_io_out ? io_r_149_b : _GEN_7648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7650 = 8'h96 == r_count_36_io_out ? io_r_150_b : _GEN_7649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7651 = 8'h97 == r_count_36_io_out ? io_r_151_b : _GEN_7650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7652 = 8'h98 == r_count_36_io_out ? io_r_152_b : _GEN_7651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7653 = 8'h99 == r_count_36_io_out ? io_r_153_b : _GEN_7652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7654 = 8'h9a == r_count_36_io_out ? io_r_154_b : _GEN_7653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7655 = 8'h9b == r_count_36_io_out ? io_r_155_b : _GEN_7654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7656 = 8'h9c == r_count_36_io_out ? io_r_156_b : _GEN_7655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7657 = 8'h9d == r_count_36_io_out ? io_r_157_b : _GEN_7656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7658 = 8'h9e == r_count_36_io_out ? io_r_158_b : _GEN_7657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7659 = 8'h9f == r_count_36_io_out ? io_r_159_b : _GEN_7658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7660 = 8'ha0 == r_count_36_io_out ? io_r_160_b : _GEN_7659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7661 = 8'ha1 == r_count_36_io_out ? io_r_161_b : _GEN_7660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7662 = 8'ha2 == r_count_36_io_out ? io_r_162_b : _GEN_7661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7663 = 8'ha3 == r_count_36_io_out ? io_r_163_b : _GEN_7662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7664 = 8'ha4 == r_count_36_io_out ? io_r_164_b : _GEN_7663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7665 = 8'ha5 == r_count_36_io_out ? io_r_165_b : _GEN_7664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7666 = 8'ha6 == r_count_36_io_out ? io_r_166_b : _GEN_7665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7667 = 8'ha7 == r_count_36_io_out ? io_r_167_b : _GEN_7666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7668 = 8'ha8 == r_count_36_io_out ? io_r_168_b : _GEN_7667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7669 = 8'ha9 == r_count_36_io_out ? io_r_169_b : _GEN_7668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7670 = 8'haa == r_count_36_io_out ? io_r_170_b : _GEN_7669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7671 = 8'hab == r_count_36_io_out ? io_r_171_b : _GEN_7670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7672 = 8'hac == r_count_36_io_out ? io_r_172_b : _GEN_7671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7673 = 8'had == r_count_36_io_out ? io_r_173_b : _GEN_7672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7674 = 8'hae == r_count_36_io_out ? io_r_174_b : _GEN_7673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7675 = 8'haf == r_count_36_io_out ? io_r_175_b : _GEN_7674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7676 = 8'hb0 == r_count_36_io_out ? io_r_176_b : _GEN_7675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7677 = 8'hb1 == r_count_36_io_out ? io_r_177_b : _GEN_7676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7678 = 8'hb2 == r_count_36_io_out ? io_r_178_b : _GEN_7677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7679 = 8'hb3 == r_count_36_io_out ? io_r_179_b : _GEN_7678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7680 = 8'hb4 == r_count_36_io_out ? io_r_180_b : _GEN_7679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7681 = 8'hb5 == r_count_36_io_out ? io_r_181_b : _GEN_7680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7682 = 8'hb6 == r_count_36_io_out ? io_r_182_b : _GEN_7681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7683 = 8'hb7 == r_count_36_io_out ? io_r_183_b : _GEN_7682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7684 = 8'hb8 == r_count_36_io_out ? io_r_184_b : _GEN_7683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7685 = 8'hb9 == r_count_36_io_out ? io_r_185_b : _GEN_7684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7686 = 8'hba == r_count_36_io_out ? io_r_186_b : _GEN_7685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7687 = 8'hbb == r_count_36_io_out ? io_r_187_b : _GEN_7686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7688 = 8'hbc == r_count_36_io_out ? io_r_188_b : _GEN_7687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7689 = 8'hbd == r_count_36_io_out ? io_r_189_b : _GEN_7688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7690 = 8'hbe == r_count_36_io_out ? io_r_190_b : _GEN_7689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7691 = 8'hbf == r_count_36_io_out ? io_r_191_b : _GEN_7690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7692 = 8'hc0 == r_count_36_io_out ? io_r_192_b : _GEN_7691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7693 = 8'hc1 == r_count_36_io_out ? io_r_193_b : _GEN_7692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7694 = 8'hc2 == r_count_36_io_out ? io_r_194_b : _GEN_7693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7695 = 8'hc3 == r_count_36_io_out ? io_r_195_b : _GEN_7694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7696 = 8'hc4 == r_count_36_io_out ? io_r_196_b : _GEN_7695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7697 = 8'hc5 == r_count_36_io_out ? io_r_197_b : _GEN_7696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7698 = 8'hc6 == r_count_36_io_out ? io_r_198_b : _GEN_7697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7701 = 8'h1 == r_count_37_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7702 = 8'h2 == r_count_37_io_out ? io_r_2_b : _GEN_7701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7703 = 8'h3 == r_count_37_io_out ? io_r_3_b : _GEN_7702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7704 = 8'h4 == r_count_37_io_out ? io_r_4_b : _GEN_7703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7705 = 8'h5 == r_count_37_io_out ? io_r_5_b : _GEN_7704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7706 = 8'h6 == r_count_37_io_out ? io_r_6_b : _GEN_7705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7707 = 8'h7 == r_count_37_io_out ? io_r_7_b : _GEN_7706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7708 = 8'h8 == r_count_37_io_out ? io_r_8_b : _GEN_7707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7709 = 8'h9 == r_count_37_io_out ? io_r_9_b : _GEN_7708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7710 = 8'ha == r_count_37_io_out ? io_r_10_b : _GEN_7709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7711 = 8'hb == r_count_37_io_out ? io_r_11_b : _GEN_7710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7712 = 8'hc == r_count_37_io_out ? io_r_12_b : _GEN_7711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7713 = 8'hd == r_count_37_io_out ? io_r_13_b : _GEN_7712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7714 = 8'he == r_count_37_io_out ? io_r_14_b : _GEN_7713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7715 = 8'hf == r_count_37_io_out ? io_r_15_b : _GEN_7714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7716 = 8'h10 == r_count_37_io_out ? io_r_16_b : _GEN_7715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7717 = 8'h11 == r_count_37_io_out ? io_r_17_b : _GEN_7716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7718 = 8'h12 == r_count_37_io_out ? io_r_18_b : _GEN_7717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7719 = 8'h13 == r_count_37_io_out ? io_r_19_b : _GEN_7718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7720 = 8'h14 == r_count_37_io_out ? io_r_20_b : _GEN_7719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7721 = 8'h15 == r_count_37_io_out ? io_r_21_b : _GEN_7720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7722 = 8'h16 == r_count_37_io_out ? io_r_22_b : _GEN_7721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7723 = 8'h17 == r_count_37_io_out ? io_r_23_b : _GEN_7722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7724 = 8'h18 == r_count_37_io_out ? io_r_24_b : _GEN_7723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7725 = 8'h19 == r_count_37_io_out ? io_r_25_b : _GEN_7724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7726 = 8'h1a == r_count_37_io_out ? io_r_26_b : _GEN_7725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7727 = 8'h1b == r_count_37_io_out ? io_r_27_b : _GEN_7726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7728 = 8'h1c == r_count_37_io_out ? io_r_28_b : _GEN_7727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7729 = 8'h1d == r_count_37_io_out ? io_r_29_b : _GEN_7728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7730 = 8'h1e == r_count_37_io_out ? io_r_30_b : _GEN_7729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7731 = 8'h1f == r_count_37_io_out ? io_r_31_b : _GEN_7730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7732 = 8'h20 == r_count_37_io_out ? io_r_32_b : _GEN_7731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7733 = 8'h21 == r_count_37_io_out ? io_r_33_b : _GEN_7732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7734 = 8'h22 == r_count_37_io_out ? io_r_34_b : _GEN_7733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7735 = 8'h23 == r_count_37_io_out ? io_r_35_b : _GEN_7734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7736 = 8'h24 == r_count_37_io_out ? io_r_36_b : _GEN_7735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7737 = 8'h25 == r_count_37_io_out ? io_r_37_b : _GEN_7736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7738 = 8'h26 == r_count_37_io_out ? io_r_38_b : _GEN_7737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7739 = 8'h27 == r_count_37_io_out ? io_r_39_b : _GEN_7738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7740 = 8'h28 == r_count_37_io_out ? io_r_40_b : _GEN_7739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7741 = 8'h29 == r_count_37_io_out ? io_r_41_b : _GEN_7740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7742 = 8'h2a == r_count_37_io_out ? io_r_42_b : _GEN_7741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7743 = 8'h2b == r_count_37_io_out ? io_r_43_b : _GEN_7742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7744 = 8'h2c == r_count_37_io_out ? io_r_44_b : _GEN_7743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7745 = 8'h2d == r_count_37_io_out ? io_r_45_b : _GEN_7744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7746 = 8'h2e == r_count_37_io_out ? io_r_46_b : _GEN_7745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7747 = 8'h2f == r_count_37_io_out ? io_r_47_b : _GEN_7746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7748 = 8'h30 == r_count_37_io_out ? io_r_48_b : _GEN_7747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7749 = 8'h31 == r_count_37_io_out ? io_r_49_b : _GEN_7748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7750 = 8'h32 == r_count_37_io_out ? io_r_50_b : _GEN_7749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7751 = 8'h33 == r_count_37_io_out ? io_r_51_b : _GEN_7750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7752 = 8'h34 == r_count_37_io_out ? io_r_52_b : _GEN_7751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7753 = 8'h35 == r_count_37_io_out ? io_r_53_b : _GEN_7752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7754 = 8'h36 == r_count_37_io_out ? io_r_54_b : _GEN_7753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7755 = 8'h37 == r_count_37_io_out ? io_r_55_b : _GEN_7754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7756 = 8'h38 == r_count_37_io_out ? io_r_56_b : _GEN_7755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7757 = 8'h39 == r_count_37_io_out ? io_r_57_b : _GEN_7756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7758 = 8'h3a == r_count_37_io_out ? io_r_58_b : _GEN_7757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7759 = 8'h3b == r_count_37_io_out ? io_r_59_b : _GEN_7758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7760 = 8'h3c == r_count_37_io_out ? io_r_60_b : _GEN_7759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7761 = 8'h3d == r_count_37_io_out ? io_r_61_b : _GEN_7760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7762 = 8'h3e == r_count_37_io_out ? io_r_62_b : _GEN_7761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7763 = 8'h3f == r_count_37_io_out ? io_r_63_b : _GEN_7762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7764 = 8'h40 == r_count_37_io_out ? io_r_64_b : _GEN_7763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7765 = 8'h41 == r_count_37_io_out ? io_r_65_b : _GEN_7764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7766 = 8'h42 == r_count_37_io_out ? io_r_66_b : _GEN_7765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7767 = 8'h43 == r_count_37_io_out ? io_r_67_b : _GEN_7766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7768 = 8'h44 == r_count_37_io_out ? io_r_68_b : _GEN_7767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7769 = 8'h45 == r_count_37_io_out ? io_r_69_b : _GEN_7768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7770 = 8'h46 == r_count_37_io_out ? io_r_70_b : _GEN_7769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7771 = 8'h47 == r_count_37_io_out ? io_r_71_b : _GEN_7770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7772 = 8'h48 == r_count_37_io_out ? io_r_72_b : _GEN_7771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7773 = 8'h49 == r_count_37_io_out ? io_r_73_b : _GEN_7772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7774 = 8'h4a == r_count_37_io_out ? io_r_74_b : _GEN_7773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7775 = 8'h4b == r_count_37_io_out ? io_r_75_b : _GEN_7774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7776 = 8'h4c == r_count_37_io_out ? io_r_76_b : _GEN_7775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7777 = 8'h4d == r_count_37_io_out ? io_r_77_b : _GEN_7776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7778 = 8'h4e == r_count_37_io_out ? io_r_78_b : _GEN_7777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7779 = 8'h4f == r_count_37_io_out ? io_r_79_b : _GEN_7778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7780 = 8'h50 == r_count_37_io_out ? io_r_80_b : _GEN_7779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7781 = 8'h51 == r_count_37_io_out ? io_r_81_b : _GEN_7780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7782 = 8'h52 == r_count_37_io_out ? io_r_82_b : _GEN_7781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7783 = 8'h53 == r_count_37_io_out ? io_r_83_b : _GEN_7782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7784 = 8'h54 == r_count_37_io_out ? io_r_84_b : _GEN_7783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7785 = 8'h55 == r_count_37_io_out ? io_r_85_b : _GEN_7784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7786 = 8'h56 == r_count_37_io_out ? io_r_86_b : _GEN_7785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7787 = 8'h57 == r_count_37_io_out ? io_r_87_b : _GEN_7786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7788 = 8'h58 == r_count_37_io_out ? io_r_88_b : _GEN_7787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7789 = 8'h59 == r_count_37_io_out ? io_r_89_b : _GEN_7788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7790 = 8'h5a == r_count_37_io_out ? io_r_90_b : _GEN_7789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7791 = 8'h5b == r_count_37_io_out ? io_r_91_b : _GEN_7790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7792 = 8'h5c == r_count_37_io_out ? io_r_92_b : _GEN_7791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7793 = 8'h5d == r_count_37_io_out ? io_r_93_b : _GEN_7792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7794 = 8'h5e == r_count_37_io_out ? io_r_94_b : _GEN_7793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7795 = 8'h5f == r_count_37_io_out ? io_r_95_b : _GEN_7794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7796 = 8'h60 == r_count_37_io_out ? io_r_96_b : _GEN_7795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7797 = 8'h61 == r_count_37_io_out ? io_r_97_b : _GEN_7796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7798 = 8'h62 == r_count_37_io_out ? io_r_98_b : _GEN_7797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7799 = 8'h63 == r_count_37_io_out ? io_r_99_b : _GEN_7798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7800 = 8'h64 == r_count_37_io_out ? io_r_100_b : _GEN_7799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7801 = 8'h65 == r_count_37_io_out ? io_r_101_b : _GEN_7800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7802 = 8'h66 == r_count_37_io_out ? io_r_102_b : _GEN_7801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7803 = 8'h67 == r_count_37_io_out ? io_r_103_b : _GEN_7802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7804 = 8'h68 == r_count_37_io_out ? io_r_104_b : _GEN_7803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7805 = 8'h69 == r_count_37_io_out ? io_r_105_b : _GEN_7804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7806 = 8'h6a == r_count_37_io_out ? io_r_106_b : _GEN_7805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7807 = 8'h6b == r_count_37_io_out ? io_r_107_b : _GEN_7806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7808 = 8'h6c == r_count_37_io_out ? io_r_108_b : _GEN_7807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7809 = 8'h6d == r_count_37_io_out ? io_r_109_b : _GEN_7808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7810 = 8'h6e == r_count_37_io_out ? io_r_110_b : _GEN_7809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7811 = 8'h6f == r_count_37_io_out ? io_r_111_b : _GEN_7810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7812 = 8'h70 == r_count_37_io_out ? io_r_112_b : _GEN_7811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7813 = 8'h71 == r_count_37_io_out ? io_r_113_b : _GEN_7812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7814 = 8'h72 == r_count_37_io_out ? io_r_114_b : _GEN_7813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7815 = 8'h73 == r_count_37_io_out ? io_r_115_b : _GEN_7814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7816 = 8'h74 == r_count_37_io_out ? io_r_116_b : _GEN_7815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7817 = 8'h75 == r_count_37_io_out ? io_r_117_b : _GEN_7816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7818 = 8'h76 == r_count_37_io_out ? io_r_118_b : _GEN_7817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7819 = 8'h77 == r_count_37_io_out ? io_r_119_b : _GEN_7818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7820 = 8'h78 == r_count_37_io_out ? io_r_120_b : _GEN_7819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7821 = 8'h79 == r_count_37_io_out ? io_r_121_b : _GEN_7820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7822 = 8'h7a == r_count_37_io_out ? io_r_122_b : _GEN_7821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7823 = 8'h7b == r_count_37_io_out ? io_r_123_b : _GEN_7822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7824 = 8'h7c == r_count_37_io_out ? io_r_124_b : _GEN_7823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7825 = 8'h7d == r_count_37_io_out ? io_r_125_b : _GEN_7824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7826 = 8'h7e == r_count_37_io_out ? io_r_126_b : _GEN_7825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7827 = 8'h7f == r_count_37_io_out ? io_r_127_b : _GEN_7826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7828 = 8'h80 == r_count_37_io_out ? io_r_128_b : _GEN_7827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7829 = 8'h81 == r_count_37_io_out ? io_r_129_b : _GEN_7828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7830 = 8'h82 == r_count_37_io_out ? io_r_130_b : _GEN_7829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7831 = 8'h83 == r_count_37_io_out ? io_r_131_b : _GEN_7830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7832 = 8'h84 == r_count_37_io_out ? io_r_132_b : _GEN_7831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7833 = 8'h85 == r_count_37_io_out ? io_r_133_b : _GEN_7832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7834 = 8'h86 == r_count_37_io_out ? io_r_134_b : _GEN_7833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7835 = 8'h87 == r_count_37_io_out ? io_r_135_b : _GEN_7834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7836 = 8'h88 == r_count_37_io_out ? io_r_136_b : _GEN_7835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7837 = 8'h89 == r_count_37_io_out ? io_r_137_b : _GEN_7836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7838 = 8'h8a == r_count_37_io_out ? io_r_138_b : _GEN_7837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7839 = 8'h8b == r_count_37_io_out ? io_r_139_b : _GEN_7838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7840 = 8'h8c == r_count_37_io_out ? io_r_140_b : _GEN_7839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7841 = 8'h8d == r_count_37_io_out ? io_r_141_b : _GEN_7840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7842 = 8'h8e == r_count_37_io_out ? io_r_142_b : _GEN_7841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7843 = 8'h8f == r_count_37_io_out ? io_r_143_b : _GEN_7842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7844 = 8'h90 == r_count_37_io_out ? io_r_144_b : _GEN_7843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7845 = 8'h91 == r_count_37_io_out ? io_r_145_b : _GEN_7844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7846 = 8'h92 == r_count_37_io_out ? io_r_146_b : _GEN_7845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7847 = 8'h93 == r_count_37_io_out ? io_r_147_b : _GEN_7846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7848 = 8'h94 == r_count_37_io_out ? io_r_148_b : _GEN_7847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7849 = 8'h95 == r_count_37_io_out ? io_r_149_b : _GEN_7848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7850 = 8'h96 == r_count_37_io_out ? io_r_150_b : _GEN_7849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7851 = 8'h97 == r_count_37_io_out ? io_r_151_b : _GEN_7850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7852 = 8'h98 == r_count_37_io_out ? io_r_152_b : _GEN_7851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7853 = 8'h99 == r_count_37_io_out ? io_r_153_b : _GEN_7852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7854 = 8'h9a == r_count_37_io_out ? io_r_154_b : _GEN_7853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7855 = 8'h9b == r_count_37_io_out ? io_r_155_b : _GEN_7854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7856 = 8'h9c == r_count_37_io_out ? io_r_156_b : _GEN_7855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7857 = 8'h9d == r_count_37_io_out ? io_r_157_b : _GEN_7856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7858 = 8'h9e == r_count_37_io_out ? io_r_158_b : _GEN_7857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7859 = 8'h9f == r_count_37_io_out ? io_r_159_b : _GEN_7858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7860 = 8'ha0 == r_count_37_io_out ? io_r_160_b : _GEN_7859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7861 = 8'ha1 == r_count_37_io_out ? io_r_161_b : _GEN_7860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7862 = 8'ha2 == r_count_37_io_out ? io_r_162_b : _GEN_7861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7863 = 8'ha3 == r_count_37_io_out ? io_r_163_b : _GEN_7862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7864 = 8'ha4 == r_count_37_io_out ? io_r_164_b : _GEN_7863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7865 = 8'ha5 == r_count_37_io_out ? io_r_165_b : _GEN_7864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7866 = 8'ha6 == r_count_37_io_out ? io_r_166_b : _GEN_7865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7867 = 8'ha7 == r_count_37_io_out ? io_r_167_b : _GEN_7866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7868 = 8'ha8 == r_count_37_io_out ? io_r_168_b : _GEN_7867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7869 = 8'ha9 == r_count_37_io_out ? io_r_169_b : _GEN_7868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7870 = 8'haa == r_count_37_io_out ? io_r_170_b : _GEN_7869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7871 = 8'hab == r_count_37_io_out ? io_r_171_b : _GEN_7870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7872 = 8'hac == r_count_37_io_out ? io_r_172_b : _GEN_7871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7873 = 8'had == r_count_37_io_out ? io_r_173_b : _GEN_7872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7874 = 8'hae == r_count_37_io_out ? io_r_174_b : _GEN_7873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7875 = 8'haf == r_count_37_io_out ? io_r_175_b : _GEN_7874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7876 = 8'hb0 == r_count_37_io_out ? io_r_176_b : _GEN_7875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7877 = 8'hb1 == r_count_37_io_out ? io_r_177_b : _GEN_7876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7878 = 8'hb2 == r_count_37_io_out ? io_r_178_b : _GEN_7877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7879 = 8'hb3 == r_count_37_io_out ? io_r_179_b : _GEN_7878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7880 = 8'hb4 == r_count_37_io_out ? io_r_180_b : _GEN_7879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7881 = 8'hb5 == r_count_37_io_out ? io_r_181_b : _GEN_7880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7882 = 8'hb6 == r_count_37_io_out ? io_r_182_b : _GEN_7881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7883 = 8'hb7 == r_count_37_io_out ? io_r_183_b : _GEN_7882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7884 = 8'hb8 == r_count_37_io_out ? io_r_184_b : _GEN_7883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7885 = 8'hb9 == r_count_37_io_out ? io_r_185_b : _GEN_7884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7886 = 8'hba == r_count_37_io_out ? io_r_186_b : _GEN_7885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7887 = 8'hbb == r_count_37_io_out ? io_r_187_b : _GEN_7886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7888 = 8'hbc == r_count_37_io_out ? io_r_188_b : _GEN_7887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7889 = 8'hbd == r_count_37_io_out ? io_r_189_b : _GEN_7888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7890 = 8'hbe == r_count_37_io_out ? io_r_190_b : _GEN_7889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7891 = 8'hbf == r_count_37_io_out ? io_r_191_b : _GEN_7890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7892 = 8'hc0 == r_count_37_io_out ? io_r_192_b : _GEN_7891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7893 = 8'hc1 == r_count_37_io_out ? io_r_193_b : _GEN_7892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7894 = 8'hc2 == r_count_37_io_out ? io_r_194_b : _GEN_7893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7895 = 8'hc3 == r_count_37_io_out ? io_r_195_b : _GEN_7894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7896 = 8'hc4 == r_count_37_io_out ? io_r_196_b : _GEN_7895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7897 = 8'hc5 == r_count_37_io_out ? io_r_197_b : _GEN_7896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7898 = 8'hc6 == r_count_37_io_out ? io_r_198_b : _GEN_7897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7901 = 8'h1 == r_count_38_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7902 = 8'h2 == r_count_38_io_out ? io_r_2_b : _GEN_7901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7903 = 8'h3 == r_count_38_io_out ? io_r_3_b : _GEN_7902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7904 = 8'h4 == r_count_38_io_out ? io_r_4_b : _GEN_7903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7905 = 8'h5 == r_count_38_io_out ? io_r_5_b : _GEN_7904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7906 = 8'h6 == r_count_38_io_out ? io_r_6_b : _GEN_7905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7907 = 8'h7 == r_count_38_io_out ? io_r_7_b : _GEN_7906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7908 = 8'h8 == r_count_38_io_out ? io_r_8_b : _GEN_7907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7909 = 8'h9 == r_count_38_io_out ? io_r_9_b : _GEN_7908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7910 = 8'ha == r_count_38_io_out ? io_r_10_b : _GEN_7909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7911 = 8'hb == r_count_38_io_out ? io_r_11_b : _GEN_7910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7912 = 8'hc == r_count_38_io_out ? io_r_12_b : _GEN_7911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7913 = 8'hd == r_count_38_io_out ? io_r_13_b : _GEN_7912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7914 = 8'he == r_count_38_io_out ? io_r_14_b : _GEN_7913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7915 = 8'hf == r_count_38_io_out ? io_r_15_b : _GEN_7914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7916 = 8'h10 == r_count_38_io_out ? io_r_16_b : _GEN_7915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7917 = 8'h11 == r_count_38_io_out ? io_r_17_b : _GEN_7916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7918 = 8'h12 == r_count_38_io_out ? io_r_18_b : _GEN_7917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7919 = 8'h13 == r_count_38_io_out ? io_r_19_b : _GEN_7918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7920 = 8'h14 == r_count_38_io_out ? io_r_20_b : _GEN_7919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7921 = 8'h15 == r_count_38_io_out ? io_r_21_b : _GEN_7920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7922 = 8'h16 == r_count_38_io_out ? io_r_22_b : _GEN_7921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7923 = 8'h17 == r_count_38_io_out ? io_r_23_b : _GEN_7922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7924 = 8'h18 == r_count_38_io_out ? io_r_24_b : _GEN_7923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7925 = 8'h19 == r_count_38_io_out ? io_r_25_b : _GEN_7924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7926 = 8'h1a == r_count_38_io_out ? io_r_26_b : _GEN_7925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7927 = 8'h1b == r_count_38_io_out ? io_r_27_b : _GEN_7926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7928 = 8'h1c == r_count_38_io_out ? io_r_28_b : _GEN_7927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7929 = 8'h1d == r_count_38_io_out ? io_r_29_b : _GEN_7928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7930 = 8'h1e == r_count_38_io_out ? io_r_30_b : _GEN_7929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7931 = 8'h1f == r_count_38_io_out ? io_r_31_b : _GEN_7930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7932 = 8'h20 == r_count_38_io_out ? io_r_32_b : _GEN_7931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7933 = 8'h21 == r_count_38_io_out ? io_r_33_b : _GEN_7932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7934 = 8'h22 == r_count_38_io_out ? io_r_34_b : _GEN_7933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7935 = 8'h23 == r_count_38_io_out ? io_r_35_b : _GEN_7934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7936 = 8'h24 == r_count_38_io_out ? io_r_36_b : _GEN_7935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7937 = 8'h25 == r_count_38_io_out ? io_r_37_b : _GEN_7936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7938 = 8'h26 == r_count_38_io_out ? io_r_38_b : _GEN_7937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7939 = 8'h27 == r_count_38_io_out ? io_r_39_b : _GEN_7938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7940 = 8'h28 == r_count_38_io_out ? io_r_40_b : _GEN_7939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7941 = 8'h29 == r_count_38_io_out ? io_r_41_b : _GEN_7940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7942 = 8'h2a == r_count_38_io_out ? io_r_42_b : _GEN_7941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7943 = 8'h2b == r_count_38_io_out ? io_r_43_b : _GEN_7942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7944 = 8'h2c == r_count_38_io_out ? io_r_44_b : _GEN_7943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7945 = 8'h2d == r_count_38_io_out ? io_r_45_b : _GEN_7944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7946 = 8'h2e == r_count_38_io_out ? io_r_46_b : _GEN_7945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7947 = 8'h2f == r_count_38_io_out ? io_r_47_b : _GEN_7946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7948 = 8'h30 == r_count_38_io_out ? io_r_48_b : _GEN_7947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7949 = 8'h31 == r_count_38_io_out ? io_r_49_b : _GEN_7948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7950 = 8'h32 == r_count_38_io_out ? io_r_50_b : _GEN_7949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7951 = 8'h33 == r_count_38_io_out ? io_r_51_b : _GEN_7950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7952 = 8'h34 == r_count_38_io_out ? io_r_52_b : _GEN_7951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7953 = 8'h35 == r_count_38_io_out ? io_r_53_b : _GEN_7952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7954 = 8'h36 == r_count_38_io_out ? io_r_54_b : _GEN_7953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7955 = 8'h37 == r_count_38_io_out ? io_r_55_b : _GEN_7954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7956 = 8'h38 == r_count_38_io_out ? io_r_56_b : _GEN_7955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7957 = 8'h39 == r_count_38_io_out ? io_r_57_b : _GEN_7956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7958 = 8'h3a == r_count_38_io_out ? io_r_58_b : _GEN_7957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7959 = 8'h3b == r_count_38_io_out ? io_r_59_b : _GEN_7958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7960 = 8'h3c == r_count_38_io_out ? io_r_60_b : _GEN_7959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7961 = 8'h3d == r_count_38_io_out ? io_r_61_b : _GEN_7960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7962 = 8'h3e == r_count_38_io_out ? io_r_62_b : _GEN_7961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7963 = 8'h3f == r_count_38_io_out ? io_r_63_b : _GEN_7962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7964 = 8'h40 == r_count_38_io_out ? io_r_64_b : _GEN_7963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7965 = 8'h41 == r_count_38_io_out ? io_r_65_b : _GEN_7964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7966 = 8'h42 == r_count_38_io_out ? io_r_66_b : _GEN_7965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7967 = 8'h43 == r_count_38_io_out ? io_r_67_b : _GEN_7966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7968 = 8'h44 == r_count_38_io_out ? io_r_68_b : _GEN_7967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7969 = 8'h45 == r_count_38_io_out ? io_r_69_b : _GEN_7968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7970 = 8'h46 == r_count_38_io_out ? io_r_70_b : _GEN_7969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7971 = 8'h47 == r_count_38_io_out ? io_r_71_b : _GEN_7970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7972 = 8'h48 == r_count_38_io_out ? io_r_72_b : _GEN_7971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7973 = 8'h49 == r_count_38_io_out ? io_r_73_b : _GEN_7972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7974 = 8'h4a == r_count_38_io_out ? io_r_74_b : _GEN_7973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7975 = 8'h4b == r_count_38_io_out ? io_r_75_b : _GEN_7974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7976 = 8'h4c == r_count_38_io_out ? io_r_76_b : _GEN_7975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7977 = 8'h4d == r_count_38_io_out ? io_r_77_b : _GEN_7976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7978 = 8'h4e == r_count_38_io_out ? io_r_78_b : _GEN_7977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7979 = 8'h4f == r_count_38_io_out ? io_r_79_b : _GEN_7978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7980 = 8'h50 == r_count_38_io_out ? io_r_80_b : _GEN_7979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7981 = 8'h51 == r_count_38_io_out ? io_r_81_b : _GEN_7980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7982 = 8'h52 == r_count_38_io_out ? io_r_82_b : _GEN_7981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7983 = 8'h53 == r_count_38_io_out ? io_r_83_b : _GEN_7982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7984 = 8'h54 == r_count_38_io_out ? io_r_84_b : _GEN_7983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7985 = 8'h55 == r_count_38_io_out ? io_r_85_b : _GEN_7984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7986 = 8'h56 == r_count_38_io_out ? io_r_86_b : _GEN_7985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7987 = 8'h57 == r_count_38_io_out ? io_r_87_b : _GEN_7986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7988 = 8'h58 == r_count_38_io_out ? io_r_88_b : _GEN_7987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7989 = 8'h59 == r_count_38_io_out ? io_r_89_b : _GEN_7988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7990 = 8'h5a == r_count_38_io_out ? io_r_90_b : _GEN_7989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7991 = 8'h5b == r_count_38_io_out ? io_r_91_b : _GEN_7990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7992 = 8'h5c == r_count_38_io_out ? io_r_92_b : _GEN_7991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7993 = 8'h5d == r_count_38_io_out ? io_r_93_b : _GEN_7992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7994 = 8'h5e == r_count_38_io_out ? io_r_94_b : _GEN_7993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7995 = 8'h5f == r_count_38_io_out ? io_r_95_b : _GEN_7994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7996 = 8'h60 == r_count_38_io_out ? io_r_96_b : _GEN_7995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7997 = 8'h61 == r_count_38_io_out ? io_r_97_b : _GEN_7996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7998 = 8'h62 == r_count_38_io_out ? io_r_98_b : _GEN_7997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7999 = 8'h63 == r_count_38_io_out ? io_r_99_b : _GEN_7998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8000 = 8'h64 == r_count_38_io_out ? io_r_100_b : _GEN_7999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8001 = 8'h65 == r_count_38_io_out ? io_r_101_b : _GEN_8000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8002 = 8'h66 == r_count_38_io_out ? io_r_102_b : _GEN_8001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8003 = 8'h67 == r_count_38_io_out ? io_r_103_b : _GEN_8002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8004 = 8'h68 == r_count_38_io_out ? io_r_104_b : _GEN_8003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8005 = 8'h69 == r_count_38_io_out ? io_r_105_b : _GEN_8004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8006 = 8'h6a == r_count_38_io_out ? io_r_106_b : _GEN_8005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8007 = 8'h6b == r_count_38_io_out ? io_r_107_b : _GEN_8006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8008 = 8'h6c == r_count_38_io_out ? io_r_108_b : _GEN_8007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8009 = 8'h6d == r_count_38_io_out ? io_r_109_b : _GEN_8008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8010 = 8'h6e == r_count_38_io_out ? io_r_110_b : _GEN_8009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8011 = 8'h6f == r_count_38_io_out ? io_r_111_b : _GEN_8010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8012 = 8'h70 == r_count_38_io_out ? io_r_112_b : _GEN_8011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8013 = 8'h71 == r_count_38_io_out ? io_r_113_b : _GEN_8012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8014 = 8'h72 == r_count_38_io_out ? io_r_114_b : _GEN_8013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8015 = 8'h73 == r_count_38_io_out ? io_r_115_b : _GEN_8014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8016 = 8'h74 == r_count_38_io_out ? io_r_116_b : _GEN_8015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8017 = 8'h75 == r_count_38_io_out ? io_r_117_b : _GEN_8016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8018 = 8'h76 == r_count_38_io_out ? io_r_118_b : _GEN_8017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8019 = 8'h77 == r_count_38_io_out ? io_r_119_b : _GEN_8018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8020 = 8'h78 == r_count_38_io_out ? io_r_120_b : _GEN_8019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8021 = 8'h79 == r_count_38_io_out ? io_r_121_b : _GEN_8020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8022 = 8'h7a == r_count_38_io_out ? io_r_122_b : _GEN_8021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8023 = 8'h7b == r_count_38_io_out ? io_r_123_b : _GEN_8022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8024 = 8'h7c == r_count_38_io_out ? io_r_124_b : _GEN_8023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8025 = 8'h7d == r_count_38_io_out ? io_r_125_b : _GEN_8024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8026 = 8'h7e == r_count_38_io_out ? io_r_126_b : _GEN_8025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8027 = 8'h7f == r_count_38_io_out ? io_r_127_b : _GEN_8026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8028 = 8'h80 == r_count_38_io_out ? io_r_128_b : _GEN_8027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8029 = 8'h81 == r_count_38_io_out ? io_r_129_b : _GEN_8028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8030 = 8'h82 == r_count_38_io_out ? io_r_130_b : _GEN_8029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8031 = 8'h83 == r_count_38_io_out ? io_r_131_b : _GEN_8030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8032 = 8'h84 == r_count_38_io_out ? io_r_132_b : _GEN_8031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8033 = 8'h85 == r_count_38_io_out ? io_r_133_b : _GEN_8032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8034 = 8'h86 == r_count_38_io_out ? io_r_134_b : _GEN_8033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8035 = 8'h87 == r_count_38_io_out ? io_r_135_b : _GEN_8034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8036 = 8'h88 == r_count_38_io_out ? io_r_136_b : _GEN_8035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8037 = 8'h89 == r_count_38_io_out ? io_r_137_b : _GEN_8036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8038 = 8'h8a == r_count_38_io_out ? io_r_138_b : _GEN_8037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8039 = 8'h8b == r_count_38_io_out ? io_r_139_b : _GEN_8038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8040 = 8'h8c == r_count_38_io_out ? io_r_140_b : _GEN_8039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8041 = 8'h8d == r_count_38_io_out ? io_r_141_b : _GEN_8040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8042 = 8'h8e == r_count_38_io_out ? io_r_142_b : _GEN_8041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8043 = 8'h8f == r_count_38_io_out ? io_r_143_b : _GEN_8042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8044 = 8'h90 == r_count_38_io_out ? io_r_144_b : _GEN_8043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8045 = 8'h91 == r_count_38_io_out ? io_r_145_b : _GEN_8044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8046 = 8'h92 == r_count_38_io_out ? io_r_146_b : _GEN_8045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8047 = 8'h93 == r_count_38_io_out ? io_r_147_b : _GEN_8046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8048 = 8'h94 == r_count_38_io_out ? io_r_148_b : _GEN_8047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8049 = 8'h95 == r_count_38_io_out ? io_r_149_b : _GEN_8048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8050 = 8'h96 == r_count_38_io_out ? io_r_150_b : _GEN_8049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8051 = 8'h97 == r_count_38_io_out ? io_r_151_b : _GEN_8050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8052 = 8'h98 == r_count_38_io_out ? io_r_152_b : _GEN_8051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8053 = 8'h99 == r_count_38_io_out ? io_r_153_b : _GEN_8052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8054 = 8'h9a == r_count_38_io_out ? io_r_154_b : _GEN_8053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8055 = 8'h9b == r_count_38_io_out ? io_r_155_b : _GEN_8054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8056 = 8'h9c == r_count_38_io_out ? io_r_156_b : _GEN_8055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8057 = 8'h9d == r_count_38_io_out ? io_r_157_b : _GEN_8056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8058 = 8'h9e == r_count_38_io_out ? io_r_158_b : _GEN_8057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8059 = 8'h9f == r_count_38_io_out ? io_r_159_b : _GEN_8058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8060 = 8'ha0 == r_count_38_io_out ? io_r_160_b : _GEN_8059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8061 = 8'ha1 == r_count_38_io_out ? io_r_161_b : _GEN_8060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8062 = 8'ha2 == r_count_38_io_out ? io_r_162_b : _GEN_8061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8063 = 8'ha3 == r_count_38_io_out ? io_r_163_b : _GEN_8062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8064 = 8'ha4 == r_count_38_io_out ? io_r_164_b : _GEN_8063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8065 = 8'ha5 == r_count_38_io_out ? io_r_165_b : _GEN_8064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8066 = 8'ha6 == r_count_38_io_out ? io_r_166_b : _GEN_8065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8067 = 8'ha7 == r_count_38_io_out ? io_r_167_b : _GEN_8066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8068 = 8'ha8 == r_count_38_io_out ? io_r_168_b : _GEN_8067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8069 = 8'ha9 == r_count_38_io_out ? io_r_169_b : _GEN_8068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8070 = 8'haa == r_count_38_io_out ? io_r_170_b : _GEN_8069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8071 = 8'hab == r_count_38_io_out ? io_r_171_b : _GEN_8070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8072 = 8'hac == r_count_38_io_out ? io_r_172_b : _GEN_8071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8073 = 8'had == r_count_38_io_out ? io_r_173_b : _GEN_8072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8074 = 8'hae == r_count_38_io_out ? io_r_174_b : _GEN_8073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8075 = 8'haf == r_count_38_io_out ? io_r_175_b : _GEN_8074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8076 = 8'hb0 == r_count_38_io_out ? io_r_176_b : _GEN_8075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8077 = 8'hb1 == r_count_38_io_out ? io_r_177_b : _GEN_8076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8078 = 8'hb2 == r_count_38_io_out ? io_r_178_b : _GEN_8077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8079 = 8'hb3 == r_count_38_io_out ? io_r_179_b : _GEN_8078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8080 = 8'hb4 == r_count_38_io_out ? io_r_180_b : _GEN_8079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8081 = 8'hb5 == r_count_38_io_out ? io_r_181_b : _GEN_8080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8082 = 8'hb6 == r_count_38_io_out ? io_r_182_b : _GEN_8081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8083 = 8'hb7 == r_count_38_io_out ? io_r_183_b : _GEN_8082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8084 = 8'hb8 == r_count_38_io_out ? io_r_184_b : _GEN_8083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8085 = 8'hb9 == r_count_38_io_out ? io_r_185_b : _GEN_8084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8086 = 8'hba == r_count_38_io_out ? io_r_186_b : _GEN_8085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8087 = 8'hbb == r_count_38_io_out ? io_r_187_b : _GEN_8086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8088 = 8'hbc == r_count_38_io_out ? io_r_188_b : _GEN_8087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8089 = 8'hbd == r_count_38_io_out ? io_r_189_b : _GEN_8088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8090 = 8'hbe == r_count_38_io_out ? io_r_190_b : _GEN_8089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8091 = 8'hbf == r_count_38_io_out ? io_r_191_b : _GEN_8090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8092 = 8'hc0 == r_count_38_io_out ? io_r_192_b : _GEN_8091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8093 = 8'hc1 == r_count_38_io_out ? io_r_193_b : _GEN_8092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8094 = 8'hc2 == r_count_38_io_out ? io_r_194_b : _GEN_8093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8095 = 8'hc3 == r_count_38_io_out ? io_r_195_b : _GEN_8094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8096 = 8'hc4 == r_count_38_io_out ? io_r_196_b : _GEN_8095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8097 = 8'hc5 == r_count_38_io_out ? io_r_197_b : _GEN_8096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8098 = 8'hc6 == r_count_38_io_out ? io_r_198_b : _GEN_8097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8101 = 8'h1 == r_count_39_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8102 = 8'h2 == r_count_39_io_out ? io_r_2_b : _GEN_8101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8103 = 8'h3 == r_count_39_io_out ? io_r_3_b : _GEN_8102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8104 = 8'h4 == r_count_39_io_out ? io_r_4_b : _GEN_8103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8105 = 8'h5 == r_count_39_io_out ? io_r_5_b : _GEN_8104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8106 = 8'h6 == r_count_39_io_out ? io_r_6_b : _GEN_8105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8107 = 8'h7 == r_count_39_io_out ? io_r_7_b : _GEN_8106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8108 = 8'h8 == r_count_39_io_out ? io_r_8_b : _GEN_8107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8109 = 8'h9 == r_count_39_io_out ? io_r_9_b : _GEN_8108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8110 = 8'ha == r_count_39_io_out ? io_r_10_b : _GEN_8109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8111 = 8'hb == r_count_39_io_out ? io_r_11_b : _GEN_8110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8112 = 8'hc == r_count_39_io_out ? io_r_12_b : _GEN_8111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8113 = 8'hd == r_count_39_io_out ? io_r_13_b : _GEN_8112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8114 = 8'he == r_count_39_io_out ? io_r_14_b : _GEN_8113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8115 = 8'hf == r_count_39_io_out ? io_r_15_b : _GEN_8114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8116 = 8'h10 == r_count_39_io_out ? io_r_16_b : _GEN_8115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8117 = 8'h11 == r_count_39_io_out ? io_r_17_b : _GEN_8116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8118 = 8'h12 == r_count_39_io_out ? io_r_18_b : _GEN_8117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8119 = 8'h13 == r_count_39_io_out ? io_r_19_b : _GEN_8118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8120 = 8'h14 == r_count_39_io_out ? io_r_20_b : _GEN_8119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8121 = 8'h15 == r_count_39_io_out ? io_r_21_b : _GEN_8120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8122 = 8'h16 == r_count_39_io_out ? io_r_22_b : _GEN_8121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8123 = 8'h17 == r_count_39_io_out ? io_r_23_b : _GEN_8122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8124 = 8'h18 == r_count_39_io_out ? io_r_24_b : _GEN_8123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8125 = 8'h19 == r_count_39_io_out ? io_r_25_b : _GEN_8124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8126 = 8'h1a == r_count_39_io_out ? io_r_26_b : _GEN_8125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8127 = 8'h1b == r_count_39_io_out ? io_r_27_b : _GEN_8126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8128 = 8'h1c == r_count_39_io_out ? io_r_28_b : _GEN_8127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8129 = 8'h1d == r_count_39_io_out ? io_r_29_b : _GEN_8128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8130 = 8'h1e == r_count_39_io_out ? io_r_30_b : _GEN_8129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8131 = 8'h1f == r_count_39_io_out ? io_r_31_b : _GEN_8130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8132 = 8'h20 == r_count_39_io_out ? io_r_32_b : _GEN_8131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8133 = 8'h21 == r_count_39_io_out ? io_r_33_b : _GEN_8132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8134 = 8'h22 == r_count_39_io_out ? io_r_34_b : _GEN_8133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8135 = 8'h23 == r_count_39_io_out ? io_r_35_b : _GEN_8134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8136 = 8'h24 == r_count_39_io_out ? io_r_36_b : _GEN_8135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8137 = 8'h25 == r_count_39_io_out ? io_r_37_b : _GEN_8136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8138 = 8'h26 == r_count_39_io_out ? io_r_38_b : _GEN_8137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8139 = 8'h27 == r_count_39_io_out ? io_r_39_b : _GEN_8138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8140 = 8'h28 == r_count_39_io_out ? io_r_40_b : _GEN_8139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8141 = 8'h29 == r_count_39_io_out ? io_r_41_b : _GEN_8140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8142 = 8'h2a == r_count_39_io_out ? io_r_42_b : _GEN_8141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8143 = 8'h2b == r_count_39_io_out ? io_r_43_b : _GEN_8142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8144 = 8'h2c == r_count_39_io_out ? io_r_44_b : _GEN_8143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8145 = 8'h2d == r_count_39_io_out ? io_r_45_b : _GEN_8144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8146 = 8'h2e == r_count_39_io_out ? io_r_46_b : _GEN_8145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8147 = 8'h2f == r_count_39_io_out ? io_r_47_b : _GEN_8146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8148 = 8'h30 == r_count_39_io_out ? io_r_48_b : _GEN_8147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8149 = 8'h31 == r_count_39_io_out ? io_r_49_b : _GEN_8148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8150 = 8'h32 == r_count_39_io_out ? io_r_50_b : _GEN_8149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8151 = 8'h33 == r_count_39_io_out ? io_r_51_b : _GEN_8150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8152 = 8'h34 == r_count_39_io_out ? io_r_52_b : _GEN_8151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8153 = 8'h35 == r_count_39_io_out ? io_r_53_b : _GEN_8152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8154 = 8'h36 == r_count_39_io_out ? io_r_54_b : _GEN_8153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8155 = 8'h37 == r_count_39_io_out ? io_r_55_b : _GEN_8154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8156 = 8'h38 == r_count_39_io_out ? io_r_56_b : _GEN_8155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8157 = 8'h39 == r_count_39_io_out ? io_r_57_b : _GEN_8156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8158 = 8'h3a == r_count_39_io_out ? io_r_58_b : _GEN_8157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8159 = 8'h3b == r_count_39_io_out ? io_r_59_b : _GEN_8158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8160 = 8'h3c == r_count_39_io_out ? io_r_60_b : _GEN_8159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8161 = 8'h3d == r_count_39_io_out ? io_r_61_b : _GEN_8160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8162 = 8'h3e == r_count_39_io_out ? io_r_62_b : _GEN_8161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8163 = 8'h3f == r_count_39_io_out ? io_r_63_b : _GEN_8162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8164 = 8'h40 == r_count_39_io_out ? io_r_64_b : _GEN_8163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8165 = 8'h41 == r_count_39_io_out ? io_r_65_b : _GEN_8164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8166 = 8'h42 == r_count_39_io_out ? io_r_66_b : _GEN_8165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8167 = 8'h43 == r_count_39_io_out ? io_r_67_b : _GEN_8166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8168 = 8'h44 == r_count_39_io_out ? io_r_68_b : _GEN_8167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8169 = 8'h45 == r_count_39_io_out ? io_r_69_b : _GEN_8168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8170 = 8'h46 == r_count_39_io_out ? io_r_70_b : _GEN_8169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8171 = 8'h47 == r_count_39_io_out ? io_r_71_b : _GEN_8170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8172 = 8'h48 == r_count_39_io_out ? io_r_72_b : _GEN_8171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8173 = 8'h49 == r_count_39_io_out ? io_r_73_b : _GEN_8172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8174 = 8'h4a == r_count_39_io_out ? io_r_74_b : _GEN_8173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8175 = 8'h4b == r_count_39_io_out ? io_r_75_b : _GEN_8174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8176 = 8'h4c == r_count_39_io_out ? io_r_76_b : _GEN_8175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8177 = 8'h4d == r_count_39_io_out ? io_r_77_b : _GEN_8176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8178 = 8'h4e == r_count_39_io_out ? io_r_78_b : _GEN_8177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8179 = 8'h4f == r_count_39_io_out ? io_r_79_b : _GEN_8178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8180 = 8'h50 == r_count_39_io_out ? io_r_80_b : _GEN_8179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8181 = 8'h51 == r_count_39_io_out ? io_r_81_b : _GEN_8180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8182 = 8'h52 == r_count_39_io_out ? io_r_82_b : _GEN_8181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8183 = 8'h53 == r_count_39_io_out ? io_r_83_b : _GEN_8182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8184 = 8'h54 == r_count_39_io_out ? io_r_84_b : _GEN_8183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8185 = 8'h55 == r_count_39_io_out ? io_r_85_b : _GEN_8184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8186 = 8'h56 == r_count_39_io_out ? io_r_86_b : _GEN_8185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8187 = 8'h57 == r_count_39_io_out ? io_r_87_b : _GEN_8186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8188 = 8'h58 == r_count_39_io_out ? io_r_88_b : _GEN_8187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8189 = 8'h59 == r_count_39_io_out ? io_r_89_b : _GEN_8188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8190 = 8'h5a == r_count_39_io_out ? io_r_90_b : _GEN_8189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8191 = 8'h5b == r_count_39_io_out ? io_r_91_b : _GEN_8190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8192 = 8'h5c == r_count_39_io_out ? io_r_92_b : _GEN_8191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8193 = 8'h5d == r_count_39_io_out ? io_r_93_b : _GEN_8192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8194 = 8'h5e == r_count_39_io_out ? io_r_94_b : _GEN_8193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8195 = 8'h5f == r_count_39_io_out ? io_r_95_b : _GEN_8194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8196 = 8'h60 == r_count_39_io_out ? io_r_96_b : _GEN_8195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8197 = 8'h61 == r_count_39_io_out ? io_r_97_b : _GEN_8196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8198 = 8'h62 == r_count_39_io_out ? io_r_98_b : _GEN_8197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8199 = 8'h63 == r_count_39_io_out ? io_r_99_b : _GEN_8198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8200 = 8'h64 == r_count_39_io_out ? io_r_100_b : _GEN_8199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8201 = 8'h65 == r_count_39_io_out ? io_r_101_b : _GEN_8200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8202 = 8'h66 == r_count_39_io_out ? io_r_102_b : _GEN_8201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8203 = 8'h67 == r_count_39_io_out ? io_r_103_b : _GEN_8202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8204 = 8'h68 == r_count_39_io_out ? io_r_104_b : _GEN_8203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8205 = 8'h69 == r_count_39_io_out ? io_r_105_b : _GEN_8204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8206 = 8'h6a == r_count_39_io_out ? io_r_106_b : _GEN_8205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8207 = 8'h6b == r_count_39_io_out ? io_r_107_b : _GEN_8206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8208 = 8'h6c == r_count_39_io_out ? io_r_108_b : _GEN_8207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8209 = 8'h6d == r_count_39_io_out ? io_r_109_b : _GEN_8208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8210 = 8'h6e == r_count_39_io_out ? io_r_110_b : _GEN_8209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8211 = 8'h6f == r_count_39_io_out ? io_r_111_b : _GEN_8210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8212 = 8'h70 == r_count_39_io_out ? io_r_112_b : _GEN_8211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8213 = 8'h71 == r_count_39_io_out ? io_r_113_b : _GEN_8212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8214 = 8'h72 == r_count_39_io_out ? io_r_114_b : _GEN_8213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8215 = 8'h73 == r_count_39_io_out ? io_r_115_b : _GEN_8214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8216 = 8'h74 == r_count_39_io_out ? io_r_116_b : _GEN_8215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8217 = 8'h75 == r_count_39_io_out ? io_r_117_b : _GEN_8216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8218 = 8'h76 == r_count_39_io_out ? io_r_118_b : _GEN_8217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8219 = 8'h77 == r_count_39_io_out ? io_r_119_b : _GEN_8218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8220 = 8'h78 == r_count_39_io_out ? io_r_120_b : _GEN_8219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8221 = 8'h79 == r_count_39_io_out ? io_r_121_b : _GEN_8220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8222 = 8'h7a == r_count_39_io_out ? io_r_122_b : _GEN_8221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8223 = 8'h7b == r_count_39_io_out ? io_r_123_b : _GEN_8222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8224 = 8'h7c == r_count_39_io_out ? io_r_124_b : _GEN_8223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8225 = 8'h7d == r_count_39_io_out ? io_r_125_b : _GEN_8224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8226 = 8'h7e == r_count_39_io_out ? io_r_126_b : _GEN_8225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8227 = 8'h7f == r_count_39_io_out ? io_r_127_b : _GEN_8226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8228 = 8'h80 == r_count_39_io_out ? io_r_128_b : _GEN_8227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8229 = 8'h81 == r_count_39_io_out ? io_r_129_b : _GEN_8228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8230 = 8'h82 == r_count_39_io_out ? io_r_130_b : _GEN_8229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8231 = 8'h83 == r_count_39_io_out ? io_r_131_b : _GEN_8230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8232 = 8'h84 == r_count_39_io_out ? io_r_132_b : _GEN_8231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8233 = 8'h85 == r_count_39_io_out ? io_r_133_b : _GEN_8232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8234 = 8'h86 == r_count_39_io_out ? io_r_134_b : _GEN_8233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8235 = 8'h87 == r_count_39_io_out ? io_r_135_b : _GEN_8234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8236 = 8'h88 == r_count_39_io_out ? io_r_136_b : _GEN_8235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8237 = 8'h89 == r_count_39_io_out ? io_r_137_b : _GEN_8236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8238 = 8'h8a == r_count_39_io_out ? io_r_138_b : _GEN_8237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8239 = 8'h8b == r_count_39_io_out ? io_r_139_b : _GEN_8238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8240 = 8'h8c == r_count_39_io_out ? io_r_140_b : _GEN_8239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8241 = 8'h8d == r_count_39_io_out ? io_r_141_b : _GEN_8240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8242 = 8'h8e == r_count_39_io_out ? io_r_142_b : _GEN_8241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8243 = 8'h8f == r_count_39_io_out ? io_r_143_b : _GEN_8242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8244 = 8'h90 == r_count_39_io_out ? io_r_144_b : _GEN_8243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8245 = 8'h91 == r_count_39_io_out ? io_r_145_b : _GEN_8244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8246 = 8'h92 == r_count_39_io_out ? io_r_146_b : _GEN_8245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8247 = 8'h93 == r_count_39_io_out ? io_r_147_b : _GEN_8246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8248 = 8'h94 == r_count_39_io_out ? io_r_148_b : _GEN_8247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8249 = 8'h95 == r_count_39_io_out ? io_r_149_b : _GEN_8248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8250 = 8'h96 == r_count_39_io_out ? io_r_150_b : _GEN_8249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8251 = 8'h97 == r_count_39_io_out ? io_r_151_b : _GEN_8250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8252 = 8'h98 == r_count_39_io_out ? io_r_152_b : _GEN_8251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8253 = 8'h99 == r_count_39_io_out ? io_r_153_b : _GEN_8252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8254 = 8'h9a == r_count_39_io_out ? io_r_154_b : _GEN_8253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8255 = 8'h9b == r_count_39_io_out ? io_r_155_b : _GEN_8254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8256 = 8'h9c == r_count_39_io_out ? io_r_156_b : _GEN_8255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8257 = 8'h9d == r_count_39_io_out ? io_r_157_b : _GEN_8256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8258 = 8'h9e == r_count_39_io_out ? io_r_158_b : _GEN_8257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8259 = 8'h9f == r_count_39_io_out ? io_r_159_b : _GEN_8258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8260 = 8'ha0 == r_count_39_io_out ? io_r_160_b : _GEN_8259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8261 = 8'ha1 == r_count_39_io_out ? io_r_161_b : _GEN_8260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8262 = 8'ha2 == r_count_39_io_out ? io_r_162_b : _GEN_8261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8263 = 8'ha3 == r_count_39_io_out ? io_r_163_b : _GEN_8262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8264 = 8'ha4 == r_count_39_io_out ? io_r_164_b : _GEN_8263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8265 = 8'ha5 == r_count_39_io_out ? io_r_165_b : _GEN_8264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8266 = 8'ha6 == r_count_39_io_out ? io_r_166_b : _GEN_8265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8267 = 8'ha7 == r_count_39_io_out ? io_r_167_b : _GEN_8266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8268 = 8'ha8 == r_count_39_io_out ? io_r_168_b : _GEN_8267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8269 = 8'ha9 == r_count_39_io_out ? io_r_169_b : _GEN_8268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8270 = 8'haa == r_count_39_io_out ? io_r_170_b : _GEN_8269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8271 = 8'hab == r_count_39_io_out ? io_r_171_b : _GEN_8270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8272 = 8'hac == r_count_39_io_out ? io_r_172_b : _GEN_8271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8273 = 8'had == r_count_39_io_out ? io_r_173_b : _GEN_8272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8274 = 8'hae == r_count_39_io_out ? io_r_174_b : _GEN_8273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8275 = 8'haf == r_count_39_io_out ? io_r_175_b : _GEN_8274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8276 = 8'hb0 == r_count_39_io_out ? io_r_176_b : _GEN_8275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8277 = 8'hb1 == r_count_39_io_out ? io_r_177_b : _GEN_8276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8278 = 8'hb2 == r_count_39_io_out ? io_r_178_b : _GEN_8277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8279 = 8'hb3 == r_count_39_io_out ? io_r_179_b : _GEN_8278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8280 = 8'hb4 == r_count_39_io_out ? io_r_180_b : _GEN_8279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8281 = 8'hb5 == r_count_39_io_out ? io_r_181_b : _GEN_8280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8282 = 8'hb6 == r_count_39_io_out ? io_r_182_b : _GEN_8281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8283 = 8'hb7 == r_count_39_io_out ? io_r_183_b : _GEN_8282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8284 = 8'hb8 == r_count_39_io_out ? io_r_184_b : _GEN_8283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8285 = 8'hb9 == r_count_39_io_out ? io_r_185_b : _GEN_8284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8286 = 8'hba == r_count_39_io_out ? io_r_186_b : _GEN_8285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8287 = 8'hbb == r_count_39_io_out ? io_r_187_b : _GEN_8286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8288 = 8'hbc == r_count_39_io_out ? io_r_188_b : _GEN_8287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8289 = 8'hbd == r_count_39_io_out ? io_r_189_b : _GEN_8288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8290 = 8'hbe == r_count_39_io_out ? io_r_190_b : _GEN_8289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8291 = 8'hbf == r_count_39_io_out ? io_r_191_b : _GEN_8290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8292 = 8'hc0 == r_count_39_io_out ? io_r_192_b : _GEN_8291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8293 = 8'hc1 == r_count_39_io_out ? io_r_193_b : _GEN_8292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8294 = 8'hc2 == r_count_39_io_out ? io_r_194_b : _GEN_8293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8295 = 8'hc3 == r_count_39_io_out ? io_r_195_b : _GEN_8294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8296 = 8'hc4 == r_count_39_io_out ? io_r_196_b : _GEN_8295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8297 = 8'hc5 == r_count_39_io_out ? io_r_197_b : _GEN_8296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8298 = 8'hc6 == r_count_39_io_out ? io_r_198_b : _GEN_8297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8301 = 8'h1 == r_count_40_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8302 = 8'h2 == r_count_40_io_out ? io_r_2_b : _GEN_8301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8303 = 8'h3 == r_count_40_io_out ? io_r_3_b : _GEN_8302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8304 = 8'h4 == r_count_40_io_out ? io_r_4_b : _GEN_8303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8305 = 8'h5 == r_count_40_io_out ? io_r_5_b : _GEN_8304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8306 = 8'h6 == r_count_40_io_out ? io_r_6_b : _GEN_8305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8307 = 8'h7 == r_count_40_io_out ? io_r_7_b : _GEN_8306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8308 = 8'h8 == r_count_40_io_out ? io_r_8_b : _GEN_8307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8309 = 8'h9 == r_count_40_io_out ? io_r_9_b : _GEN_8308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8310 = 8'ha == r_count_40_io_out ? io_r_10_b : _GEN_8309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8311 = 8'hb == r_count_40_io_out ? io_r_11_b : _GEN_8310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8312 = 8'hc == r_count_40_io_out ? io_r_12_b : _GEN_8311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8313 = 8'hd == r_count_40_io_out ? io_r_13_b : _GEN_8312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8314 = 8'he == r_count_40_io_out ? io_r_14_b : _GEN_8313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8315 = 8'hf == r_count_40_io_out ? io_r_15_b : _GEN_8314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8316 = 8'h10 == r_count_40_io_out ? io_r_16_b : _GEN_8315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8317 = 8'h11 == r_count_40_io_out ? io_r_17_b : _GEN_8316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8318 = 8'h12 == r_count_40_io_out ? io_r_18_b : _GEN_8317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8319 = 8'h13 == r_count_40_io_out ? io_r_19_b : _GEN_8318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8320 = 8'h14 == r_count_40_io_out ? io_r_20_b : _GEN_8319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8321 = 8'h15 == r_count_40_io_out ? io_r_21_b : _GEN_8320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8322 = 8'h16 == r_count_40_io_out ? io_r_22_b : _GEN_8321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8323 = 8'h17 == r_count_40_io_out ? io_r_23_b : _GEN_8322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8324 = 8'h18 == r_count_40_io_out ? io_r_24_b : _GEN_8323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8325 = 8'h19 == r_count_40_io_out ? io_r_25_b : _GEN_8324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8326 = 8'h1a == r_count_40_io_out ? io_r_26_b : _GEN_8325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8327 = 8'h1b == r_count_40_io_out ? io_r_27_b : _GEN_8326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8328 = 8'h1c == r_count_40_io_out ? io_r_28_b : _GEN_8327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8329 = 8'h1d == r_count_40_io_out ? io_r_29_b : _GEN_8328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8330 = 8'h1e == r_count_40_io_out ? io_r_30_b : _GEN_8329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8331 = 8'h1f == r_count_40_io_out ? io_r_31_b : _GEN_8330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8332 = 8'h20 == r_count_40_io_out ? io_r_32_b : _GEN_8331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8333 = 8'h21 == r_count_40_io_out ? io_r_33_b : _GEN_8332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8334 = 8'h22 == r_count_40_io_out ? io_r_34_b : _GEN_8333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8335 = 8'h23 == r_count_40_io_out ? io_r_35_b : _GEN_8334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8336 = 8'h24 == r_count_40_io_out ? io_r_36_b : _GEN_8335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8337 = 8'h25 == r_count_40_io_out ? io_r_37_b : _GEN_8336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8338 = 8'h26 == r_count_40_io_out ? io_r_38_b : _GEN_8337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8339 = 8'h27 == r_count_40_io_out ? io_r_39_b : _GEN_8338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8340 = 8'h28 == r_count_40_io_out ? io_r_40_b : _GEN_8339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8341 = 8'h29 == r_count_40_io_out ? io_r_41_b : _GEN_8340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8342 = 8'h2a == r_count_40_io_out ? io_r_42_b : _GEN_8341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8343 = 8'h2b == r_count_40_io_out ? io_r_43_b : _GEN_8342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8344 = 8'h2c == r_count_40_io_out ? io_r_44_b : _GEN_8343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8345 = 8'h2d == r_count_40_io_out ? io_r_45_b : _GEN_8344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8346 = 8'h2e == r_count_40_io_out ? io_r_46_b : _GEN_8345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8347 = 8'h2f == r_count_40_io_out ? io_r_47_b : _GEN_8346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8348 = 8'h30 == r_count_40_io_out ? io_r_48_b : _GEN_8347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8349 = 8'h31 == r_count_40_io_out ? io_r_49_b : _GEN_8348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8350 = 8'h32 == r_count_40_io_out ? io_r_50_b : _GEN_8349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8351 = 8'h33 == r_count_40_io_out ? io_r_51_b : _GEN_8350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8352 = 8'h34 == r_count_40_io_out ? io_r_52_b : _GEN_8351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8353 = 8'h35 == r_count_40_io_out ? io_r_53_b : _GEN_8352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8354 = 8'h36 == r_count_40_io_out ? io_r_54_b : _GEN_8353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8355 = 8'h37 == r_count_40_io_out ? io_r_55_b : _GEN_8354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8356 = 8'h38 == r_count_40_io_out ? io_r_56_b : _GEN_8355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8357 = 8'h39 == r_count_40_io_out ? io_r_57_b : _GEN_8356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8358 = 8'h3a == r_count_40_io_out ? io_r_58_b : _GEN_8357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8359 = 8'h3b == r_count_40_io_out ? io_r_59_b : _GEN_8358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8360 = 8'h3c == r_count_40_io_out ? io_r_60_b : _GEN_8359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8361 = 8'h3d == r_count_40_io_out ? io_r_61_b : _GEN_8360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8362 = 8'h3e == r_count_40_io_out ? io_r_62_b : _GEN_8361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8363 = 8'h3f == r_count_40_io_out ? io_r_63_b : _GEN_8362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8364 = 8'h40 == r_count_40_io_out ? io_r_64_b : _GEN_8363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8365 = 8'h41 == r_count_40_io_out ? io_r_65_b : _GEN_8364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8366 = 8'h42 == r_count_40_io_out ? io_r_66_b : _GEN_8365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8367 = 8'h43 == r_count_40_io_out ? io_r_67_b : _GEN_8366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8368 = 8'h44 == r_count_40_io_out ? io_r_68_b : _GEN_8367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8369 = 8'h45 == r_count_40_io_out ? io_r_69_b : _GEN_8368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8370 = 8'h46 == r_count_40_io_out ? io_r_70_b : _GEN_8369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8371 = 8'h47 == r_count_40_io_out ? io_r_71_b : _GEN_8370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8372 = 8'h48 == r_count_40_io_out ? io_r_72_b : _GEN_8371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8373 = 8'h49 == r_count_40_io_out ? io_r_73_b : _GEN_8372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8374 = 8'h4a == r_count_40_io_out ? io_r_74_b : _GEN_8373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8375 = 8'h4b == r_count_40_io_out ? io_r_75_b : _GEN_8374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8376 = 8'h4c == r_count_40_io_out ? io_r_76_b : _GEN_8375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8377 = 8'h4d == r_count_40_io_out ? io_r_77_b : _GEN_8376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8378 = 8'h4e == r_count_40_io_out ? io_r_78_b : _GEN_8377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8379 = 8'h4f == r_count_40_io_out ? io_r_79_b : _GEN_8378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8380 = 8'h50 == r_count_40_io_out ? io_r_80_b : _GEN_8379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8381 = 8'h51 == r_count_40_io_out ? io_r_81_b : _GEN_8380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8382 = 8'h52 == r_count_40_io_out ? io_r_82_b : _GEN_8381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8383 = 8'h53 == r_count_40_io_out ? io_r_83_b : _GEN_8382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8384 = 8'h54 == r_count_40_io_out ? io_r_84_b : _GEN_8383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8385 = 8'h55 == r_count_40_io_out ? io_r_85_b : _GEN_8384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8386 = 8'h56 == r_count_40_io_out ? io_r_86_b : _GEN_8385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8387 = 8'h57 == r_count_40_io_out ? io_r_87_b : _GEN_8386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8388 = 8'h58 == r_count_40_io_out ? io_r_88_b : _GEN_8387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8389 = 8'h59 == r_count_40_io_out ? io_r_89_b : _GEN_8388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8390 = 8'h5a == r_count_40_io_out ? io_r_90_b : _GEN_8389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8391 = 8'h5b == r_count_40_io_out ? io_r_91_b : _GEN_8390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8392 = 8'h5c == r_count_40_io_out ? io_r_92_b : _GEN_8391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8393 = 8'h5d == r_count_40_io_out ? io_r_93_b : _GEN_8392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8394 = 8'h5e == r_count_40_io_out ? io_r_94_b : _GEN_8393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8395 = 8'h5f == r_count_40_io_out ? io_r_95_b : _GEN_8394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8396 = 8'h60 == r_count_40_io_out ? io_r_96_b : _GEN_8395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8397 = 8'h61 == r_count_40_io_out ? io_r_97_b : _GEN_8396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8398 = 8'h62 == r_count_40_io_out ? io_r_98_b : _GEN_8397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8399 = 8'h63 == r_count_40_io_out ? io_r_99_b : _GEN_8398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8400 = 8'h64 == r_count_40_io_out ? io_r_100_b : _GEN_8399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8401 = 8'h65 == r_count_40_io_out ? io_r_101_b : _GEN_8400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8402 = 8'h66 == r_count_40_io_out ? io_r_102_b : _GEN_8401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8403 = 8'h67 == r_count_40_io_out ? io_r_103_b : _GEN_8402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8404 = 8'h68 == r_count_40_io_out ? io_r_104_b : _GEN_8403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8405 = 8'h69 == r_count_40_io_out ? io_r_105_b : _GEN_8404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8406 = 8'h6a == r_count_40_io_out ? io_r_106_b : _GEN_8405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8407 = 8'h6b == r_count_40_io_out ? io_r_107_b : _GEN_8406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8408 = 8'h6c == r_count_40_io_out ? io_r_108_b : _GEN_8407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8409 = 8'h6d == r_count_40_io_out ? io_r_109_b : _GEN_8408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8410 = 8'h6e == r_count_40_io_out ? io_r_110_b : _GEN_8409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8411 = 8'h6f == r_count_40_io_out ? io_r_111_b : _GEN_8410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8412 = 8'h70 == r_count_40_io_out ? io_r_112_b : _GEN_8411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8413 = 8'h71 == r_count_40_io_out ? io_r_113_b : _GEN_8412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8414 = 8'h72 == r_count_40_io_out ? io_r_114_b : _GEN_8413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8415 = 8'h73 == r_count_40_io_out ? io_r_115_b : _GEN_8414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8416 = 8'h74 == r_count_40_io_out ? io_r_116_b : _GEN_8415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8417 = 8'h75 == r_count_40_io_out ? io_r_117_b : _GEN_8416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8418 = 8'h76 == r_count_40_io_out ? io_r_118_b : _GEN_8417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8419 = 8'h77 == r_count_40_io_out ? io_r_119_b : _GEN_8418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8420 = 8'h78 == r_count_40_io_out ? io_r_120_b : _GEN_8419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8421 = 8'h79 == r_count_40_io_out ? io_r_121_b : _GEN_8420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8422 = 8'h7a == r_count_40_io_out ? io_r_122_b : _GEN_8421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8423 = 8'h7b == r_count_40_io_out ? io_r_123_b : _GEN_8422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8424 = 8'h7c == r_count_40_io_out ? io_r_124_b : _GEN_8423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8425 = 8'h7d == r_count_40_io_out ? io_r_125_b : _GEN_8424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8426 = 8'h7e == r_count_40_io_out ? io_r_126_b : _GEN_8425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8427 = 8'h7f == r_count_40_io_out ? io_r_127_b : _GEN_8426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8428 = 8'h80 == r_count_40_io_out ? io_r_128_b : _GEN_8427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8429 = 8'h81 == r_count_40_io_out ? io_r_129_b : _GEN_8428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8430 = 8'h82 == r_count_40_io_out ? io_r_130_b : _GEN_8429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8431 = 8'h83 == r_count_40_io_out ? io_r_131_b : _GEN_8430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8432 = 8'h84 == r_count_40_io_out ? io_r_132_b : _GEN_8431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8433 = 8'h85 == r_count_40_io_out ? io_r_133_b : _GEN_8432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8434 = 8'h86 == r_count_40_io_out ? io_r_134_b : _GEN_8433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8435 = 8'h87 == r_count_40_io_out ? io_r_135_b : _GEN_8434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8436 = 8'h88 == r_count_40_io_out ? io_r_136_b : _GEN_8435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8437 = 8'h89 == r_count_40_io_out ? io_r_137_b : _GEN_8436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8438 = 8'h8a == r_count_40_io_out ? io_r_138_b : _GEN_8437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8439 = 8'h8b == r_count_40_io_out ? io_r_139_b : _GEN_8438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8440 = 8'h8c == r_count_40_io_out ? io_r_140_b : _GEN_8439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8441 = 8'h8d == r_count_40_io_out ? io_r_141_b : _GEN_8440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8442 = 8'h8e == r_count_40_io_out ? io_r_142_b : _GEN_8441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8443 = 8'h8f == r_count_40_io_out ? io_r_143_b : _GEN_8442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8444 = 8'h90 == r_count_40_io_out ? io_r_144_b : _GEN_8443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8445 = 8'h91 == r_count_40_io_out ? io_r_145_b : _GEN_8444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8446 = 8'h92 == r_count_40_io_out ? io_r_146_b : _GEN_8445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8447 = 8'h93 == r_count_40_io_out ? io_r_147_b : _GEN_8446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8448 = 8'h94 == r_count_40_io_out ? io_r_148_b : _GEN_8447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8449 = 8'h95 == r_count_40_io_out ? io_r_149_b : _GEN_8448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8450 = 8'h96 == r_count_40_io_out ? io_r_150_b : _GEN_8449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8451 = 8'h97 == r_count_40_io_out ? io_r_151_b : _GEN_8450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8452 = 8'h98 == r_count_40_io_out ? io_r_152_b : _GEN_8451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8453 = 8'h99 == r_count_40_io_out ? io_r_153_b : _GEN_8452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8454 = 8'h9a == r_count_40_io_out ? io_r_154_b : _GEN_8453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8455 = 8'h9b == r_count_40_io_out ? io_r_155_b : _GEN_8454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8456 = 8'h9c == r_count_40_io_out ? io_r_156_b : _GEN_8455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8457 = 8'h9d == r_count_40_io_out ? io_r_157_b : _GEN_8456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8458 = 8'h9e == r_count_40_io_out ? io_r_158_b : _GEN_8457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8459 = 8'h9f == r_count_40_io_out ? io_r_159_b : _GEN_8458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8460 = 8'ha0 == r_count_40_io_out ? io_r_160_b : _GEN_8459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8461 = 8'ha1 == r_count_40_io_out ? io_r_161_b : _GEN_8460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8462 = 8'ha2 == r_count_40_io_out ? io_r_162_b : _GEN_8461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8463 = 8'ha3 == r_count_40_io_out ? io_r_163_b : _GEN_8462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8464 = 8'ha4 == r_count_40_io_out ? io_r_164_b : _GEN_8463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8465 = 8'ha5 == r_count_40_io_out ? io_r_165_b : _GEN_8464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8466 = 8'ha6 == r_count_40_io_out ? io_r_166_b : _GEN_8465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8467 = 8'ha7 == r_count_40_io_out ? io_r_167_b : _GEN_8466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8468 = 8'ha8 == r_count_40_io_out ? io_r_168_b : _GEN_8467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8469 = 8'ha9 == r_count_40_io_out ? io_r_169_b : _GEN_8468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8470 = 8'haa == r_count_40_io_out ? io_r_170_b : _GEN_8469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8471 = 8'hab == r_count_40_io_out ? io_r_171_b : _GEN_8470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8472 = 8'hac == r_count_40_io_out ? io_r_172_b : _GEN_8471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8473 = 8'had == r_count_40_io_out ? io_r_173_b : _GEN_8472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8474 = 8'hae == r_count_40_io_out ? io_r_174_b : _GEN_8473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8475 = 8'haf == r_count_40_io_out ? io_r_175_b : _GEN_8474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8476 = 8'hb0 == r_count_40_io_out ? io_r_176_b : _GEN_8475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8477 = 8'hb1 == r_count_40_io_out ? io_r_177_b : _GEN_8476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8478 = 8'hb2 == r_count_40_io_out ? io_r_178_b : _GEN_8477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8479 = 8'hb3 == r_count_40_io_out ? io_r_179_b : _GEN_8478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8480 = 8'hb4 == r_count_40_io_out ? io_r_180_b : _GEN_8479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8481 = 8'hb5 == r_count_40_io_out ? io_r_181_b : _GEN_8480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8482 = 8'hb6 == r_count_40_io_out ? io_r_182_b : _GEN_8481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8483 = 8'hb7 == r_count_40_io_out ? io_r_183_b : _GEN_8482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8484 = 8'hb8 == r_count_40_io_out ? io_r_184_b : _GEN_8483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8485 = 8'hb9 == r_count_40_io_out ? io_r_185_b : _GEN_8484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8486 = 8'hba == r_count_40_io_out ? io_r_186_b : _GEN_8485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8487 = 8'hbb == r_count_40_io_out ? io_r_187_b : _GEN_8486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8488 = 8'hbc == r_count_40_io_out ? io_r_188_b : _GEN_8487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8489 = 8'hbd == r_count_40_io_out ? io_r_189_b : _GEN_8488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8490 = 8'hbe == r_count_40_io_out ? io_r_190_b : _GEN_8489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8491 = 8'hbf == r_count_40_io_out ? io_r_191_b : _GEN_8490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8492 = 8'hc0 == r_count_40_io_out ? io_r_192_b : _GEN_8491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8493 = 8'hc1 == r_count_40_io_out ? io_r_193_b : _GEN_8492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8494 = 8'hc2 == r_count_40_io_out ? io_r_194_b : _GEN_8493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8495 = 8'hc3 == r_count_40_io_out ? io_r_195_b : _GEN_8494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8496 = 8'hc4 == r_count_40_io_out ? io_r_196_b : _GEN_8495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8497 = 8'hc5 == r_count_40_io_out ? io_r_197_b : _GEN_8496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8498 = 8'hc6 == r_count_40_io_out ? io_r_198_b : _GEN_8497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8501 = 8'h1 == r_count_41_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8502 = 8'h2 == r_count_41_io_out ? io_r_2_b : _GEN_8501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8503 = 8'h3 == r_count_41_io_out ? io_r_3_b : _GEN_8502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8504 = 8'h4 == r_count_41_io_out ? io_r_4_b : _GEN_8503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8505 = 8'h5 == r_count_41_io_out ? io_r_5_b : _GEN_8504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8506 = 8'h6 == r_count_41_io_out ? io_r_6_b : _GEN_8505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8507 = 8'h7 == r_count_41_io_out ? io_r_7_b : _GEN_8506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8508 = 8'h8 == r_count_41_io_out ? io_r_8_b : _GEN_8507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8509 = 8'h9 == r_count_41_io_out ? io_r_9_b : _GEN_8508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8510 = 8'ha == r_count_41_io_out ? io_r_10_b : _GEN_8509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8511 = 8'hb == r_count_41_io_out ? io_r_11_b : _GEN_8510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8512 = 8'hc == r_count_41_io_out ? io_r_12_b : _GEN_8511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8513 = 8'hd == r_count_41_io_out ? io_r_13_b : _GEN_8512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8514 = 8'he == r_count_41_io_out ? io_r_14_b : _GEN_8513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8515 = 8'hf == r_count_41_io_out ? io_r_15_b : _GEN_8514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8516 = 8'h10 == r_count_41_io_out ? io_r_16_b : _GEN_8515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8517 = 8'h11 == r_count_41_io_out ? io_r_17_b : _GEN_8516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8518 = 8'h12 == r_count_41_io_out ? io_r_18_b : _GEN_8517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8519 = 8'h13 == r_count_41_io_out ? io_r_19_b : _GEN_8518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8520 = 8'h14 == r_count_41_io_out ? io_r_20_b : _GEN_8519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8521 = 8'h15 == r_count_41_io_out ? io_r_21_b : _GEN_8520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8522 = 8'h16 == r_count_41_io_out ? io_r_22_b : _GEN_8521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8523 = 8'h17 == r_count_41_io_out ? io_r_23_b : _GEN_8522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8524 = 8'h18 == r_count_41_io_out ? io_r_24_b : _GEN_8523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8525 = 8'h19 == r_count_41_io_out ? io_r_25_b : _GEN_8524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8526 = 8'h1a == r_count_41_io_out ? io_r_26_b : _GEN_8525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8527 = 8'h1b == r_count_41_io_out ? io_r_27_b : _GEN_8526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8528 = 8'h1c == r_count_41_io_out ? io_r_28_b : _GEN_8527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8529 = 8'h1d == r_count_41_io_out ? io_r_29_b : _GEN_8528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8530 = 8'h1e == r_count_41_io_out ? io_r_30_b : _GEN_8529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8531 = 8'h1f == r_count_41_io_out ? io_r_31_b : _GEN_8530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8532 = 8'h20 == r_count_41_io_out ? io_r_32_b : _GEN_8531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8533 = 8'h21 == r_count_41_io_out ? io_r_33_b : _GEN_8532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8534 = 8'h22 == r_count_41_io_out ? io_r_34_b : _GEN_8533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8535 = 8'h23 == r_count_41_io_out ? io_r_35_b : _GEN_8534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8536 = 8'h24 == r_count_41_io_out ? io_r_36_b : _GEN_8535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8537 = 8'h25 == r_count_41_io_out ? io_r_37_b : _GEN_8536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8538 = 8'h26 == r_count_41_io_out ? io_r_38_b : _GEN_8537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8539 = 8'h27 == r_count_41_io_out ? io_r_39_b : _GEN_8538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8540 = 8'h28 == r_count_41_io_out ? io_r_40_b : _GEN_8539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8541 = 8'h29 == r_count_41_io_out ? io_r_41_b : _GEN_8540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8542 = 8'h2a == r_count_41_io_out ? io_r_42_b : _GEN_8541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8543 = 8'h2b == r_count_41_io_out ? io_r_43_b : _GEN_8542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8544 = 8'h2c == r_count_41_io_out ? io_r_44_b : _GEN_8543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8545 = 8'h2d == r_count_41_io_out ? io_r_45_b : _GEN_8544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8546 = 8'h2e == r_count_41_io_out ? io_r_46_b : _GEN_8545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8547 = 8'h2f == r_count_41_io_out ? io_r_47_b : _GEN_8546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8548 = 8'h30 == r_count_41_io_out ? io_r_48_b : _GEN_8547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8549 = 8'h31 == r_count_41_io_out ? io_r_49_b : _GEN_8548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8550 = 8'h32 == r_count_41_io_out ? io_r_50_b : _GEN_8549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8551 = 8'h33 == r_count_41_io_out ? io_r_51_b : _GEN_8550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8552 = 8'h34 == r_count_41_io_out ? io_r_52_b : _GEN_8551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8553 = 8'h35 == r_count_41_io_out ? io_r_53_b : _GEN_8552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8554 = 8'h36 == r_count_41_io_out ? io_r_54_b : _GEN_8553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8555 = 8'h37 == r_count_41_io_out ? io_r_55_b : _GEN_8554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8556 = 8'h38 == r_count_41_io_out ? io_r_56_b : _GEN_8555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8557 = 8'h39 == r_count_41_io_out ? io_r_57_b : _GEN_8556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8558 = 8'h3a == r_count_41_io_out ? io_r_58_b : _GEN_8557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8559 = 8'h3b == r_count_41_io_out ? io_r_59_b : _GEN_8558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8560 = 8'h3c == r_count_41_io_out ? io_r_60_b : _GEN_8559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8561 = 8'h3d == r_count_41_io_out ? io_r_61_b : _GEN_8560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8562 = 8'h3e == r_count_41_io_out ? io_r_62_b : _GEN_8561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8563 = 8'h3f == r_count_41_io_out ? io_r_63_b : _GEN_8562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8564 = 8'h40 == r_count_41_io_out ? io_r_64_b : _GEN_8563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8565 = 8'h41 == r_count_41_io_out ? io_r_65_b : _GEN_8564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8566 = 8'h42 == r_count_41_io_out ? io_r_66_b : _GEN_8565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8567 = 8'h43 == r_count_41_io_out ? io_r_67_b : _GEN_8566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8568 = 8'h44 == r_count_41_io_out ? io_r_68_b : _GEN_8567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8569 = 8'h45 == r_count_41_io_out ? io_r_69_b : _GEN_8568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8570 = 8'h46 == r_count_41_io_out ? io_r_70_b : _GEN_8569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8571 = 8'h47 == r_count_41_io_out ? io_r_71_b : _GEN_8570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8572 = 8'h48 == r_count_41_io_out ? io_r_72_b : _GEN_8571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8573 = 8'h49 == r_count_41_io_out ? io_r_73_b : _GEN_8572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8574 = 8'h4a == r_count_41_io_out ? io_r_74_b : _GEN_8573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8575 = 8'h4b == r_count_41_io_out ? io_r_75_b : _GEN_8574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8576 = 8'h4c == r_count_41_io_out ? io_r_76_b : _GEN_8575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8577 = 8'h4d == r_count_41_io_out ? io_r_77_b : _GEN_8576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8578 = 8'h4e == r_count_41_io_out ? io_r_78_b : _GEN_8577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8579 = 8'h4f == r_count_41_io_out ? io_r_79_b : _GEN_8578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8580 = 8'h50 == r_count_41_io_out ? io_r_80_b : _GEN_8579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8581 = 8'h51 == r_count_41_io_out ? io_r_81_b : _GEN_8580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8582 = 8'h52 == r_count_41_io_out ? io_r_82_b : _GEN_8581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8583 = 8'h53 == r_count_41_io_out ? io_r_83_b : _GEN_8582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8584 = 8'h54 == r_count_41_io_out ? io_r_84_b : _GEN_8583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8585 = 8'h55 == r_count_41_io_out ? io_r_85_b : _GEN_8584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8586 = 8'h56 == r_count_41_io_out ? io_r_86_b : _GEN_8585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8587 = 8'h57 == r_count_41_io_out ? io_r_87_b : _GEN_8586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8588 = 8'h58 == r_count_41_io_out ? io_r_88_b : _GEN_8587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8589 = 8'h59 == r_count_41_io_out ? io_r_89_b : _GEN_8588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8590 = 8'h5a == r_count_41_io_out ? io_r_90_b : _GEN_8589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8591 = 8'h5b == r_count_41_io_out ? io_r_91_b : _GEN_8590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8592 = 8'h5c == r_count_41_io_out ? io_r_92_b : _GEN_8591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8593 = 8'h5d == r_count_41_io_out ? io_r_93_b : _GEN_8592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8594 = 8'h5e == r_count_41_io_out ? io_r_94_b : _GEN_8593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8595 = 8'h5f == r_count_41_io_out ? io_r_95_b : _GEN_8594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8596 = 8'h60 == r_count_41_io_out ? io_r_96_b : _GEN_8595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8597 = 8'h61 == r_count_41_io_out ? io_r_97_b : _GEN_8596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8598 = 8'h62 == r_count_41_io_out ? io_r_98_b : _GEN_8597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8599 = 8'h63 == r_count_41_io_out ? io_r_99_b : _GEN_8598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8600 = 8'h64 == r_count_41_io_out ? io_r_100_b : _GEN_8599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8601 = 8'h65 == r_count_41_io_out ? io_r_101_b : _GEN_8600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8602 = 8'h66 == r_count_41_io_out ? io_r_102_b : _GEN_8601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8603 = 8'h67 == r_count_41_io_out ? io_r_103_b : _GEN_8602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8604 = 8'h68 == r_count_41_io_out ? io_r_104_b : _GEN_8603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8605 = 8'h69 == r_count_41_io_out ? io_r_105_b : _GEN_8604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8606 = 8'h6a == r_count_41_io_out ? io_r_106_b : _GEN_8605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8607 = 8'h6b == r_count_41_io_out ? io_r_107_b : _GEN_8606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8608 = 8'h6c == r_count_41_io_out ? io_r_108_b : _GEN_8607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8609 = 8'h6d == r_count_41_io_out ? io_r_109_b : _GEN_8608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8610 = 8'h6e == r_count_41_io_out ? io_r_110_b : _GEN_8609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8611 = 8'h6f == r_count_41_io_out ? io_r_111_b : _GEN_8610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8612 = 8'h70 == r_count_41_io_out ? io_r_112_b : _GEN_8611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8613 = 8'h71 == r_count_41_io_out ? io_r_113_b : _GEN_8612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8614 = 8'h72 == r_count_41_io_out ? io_r_114_b : _GEN_8613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8615 = 8'h73 == r_count_41_io_out ? io_r_115_b : _GEN_8614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8616 = 8'h74 == r_count_41_io_out ? io_r_116_b : _GEN_8615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8617 = 8'h75 == r_count_41_io_out ? io_r_117_b : _GEN_8616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8618 = 8'h76 == r_count_41_io_out ? io_r_118_b : _GEN_8617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8619 = 8'h77 == r_count_41_io_out ? io_r_119_b : _GEN_8618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8620 = 8'h78 == r_count_41_io_out ? io_r_120_b : _GEN_8619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8621 = 8'h79 == r_count_41_io_out ? io_r_121_b : _GEN_8620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8622 = 8'h7a == r_count_41_io_out ? io_r_122_b : _GEN_8621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8623 = 8'h7b == r_count_41_io_out ? io_r_123_b : _GEN_8622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8624 = 8'h7c == r_count_41_io_out ? io_r_124_b : _GEN_8623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8625 = 8'h7d == r_count_41_io_out ? io_r_125_b : _GEN_8624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8626 = 8'h7e == r_count_41_io_out ? io_r_126_b : _GEN_8625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8627 = 8'h7f == r_count_41_io_out ? io_r_127_b : _GEN_8626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8628 = 8'h80 == r_count_41_io_out ? io_r_128_b : _GEN_8627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8629 = 8'h81 == r_count_41_io_out ? io_r_129_b : _GEN_8628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8630 = 8'h82 == r_count_41_io_out ? io_r_130_b : _GEN_8629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8631 = 8'h83 == r_count_41_io_out ? io_r_131_b : _GEN_8630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8632 = 8'h84 == r_count_41_io_out ? io_r_132_b : _GEN_8631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8633 = 8'h85 == r_count_41_io_out ? io_r_133_b : _GEN_8632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8634 = 8'h86 == r_count_41_io_out ? io_r_134_b : _GEN_8633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8635 = 8'h87 == r_count_41_io_out ? io_r_135_b : _GEN_8634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8636 = 8'h88 == r_count_41_io_out ? io_r_136_b : _GEN_8635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8637 = 8'h89 == r_count_41_io_out ? io_r_137_b : _GEN_8636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8638 = 8'h8a == r_count_41_io_out ? io_r_138_b : _GEN_8637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8639 = 8'h8b == r_count_41_io_out ? io_r_139_b : _GEN_8638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8640 = 8'h8c == r_count_41_io_out ? io_r_140_b : _GEN_8639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8641 = 8'h8d == r_count_41_io_out ? io_r_141_b : _GEN_8640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8642 = 8'h8e == r_count_41_io_out ? io_r_142_b : _GEN_8641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8643 = 8'h8f == r_count_41_io_out ? io_r_143_b : _GEN_8642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8644 = 8'h90 == r_count_41_io_out ? io_r_144_b : _GEN_8643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8645 = 8'h91 == r_count_41_io_out ? io_r_145_b : _GEN_8644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8646 = 8'h92 == r_count_41_io_out ? io_r_146_b : _GEN_8645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8647 = 8'h93 == r_count_41_io_out ? io_r_147_b : _GEN_8646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8648 = 8'h94 == r_count_41_io_out ? io_r_148_b : _GEN_8647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8649 = 8'h95 == r_count_41_io_out ? io_r_149_b : _GEN_8648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8650 = 8'h96 == r_count_41_io_out ? io_r_150_b : _GEN_8649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8651 = 8'h97 == r_count_41_io_out ? io_r_151_b : _GEN_8650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8652 = 8'h98 == r_count_41_io_out ? io_r_152_b : _GEN_8651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8653 = 8'h99 == r_count_41_io_out ? io_r_153_b : _GEN_8652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8654 = 8'h9a == r_count_41_io_out ? io_r_154_b : _GEN_8653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8655 = 8'h9b == r_count_41_io_out ? io_r_155_b : _GEN_8654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8656 = 8'h9c == r_count_41_io_out ? io_r_156_b : _GEN_8655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8657 = 8'h9d == r_count_41_io_out ? io_r_157_b : _GEN_8656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8658 = 8'h9e == r_count_41_io_out ? io_r_158_b : _GEN_8657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8659 = 8'h9f == r_count_41_io_out ? io_r_159_b : _GEN_8658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8660 = 8'ha0 == r_count_41_io_out ? io_r_160_b : _GEN_8659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8661 = 8'ha1 == r_count_41_io_out ? io_r_161_b : _GEN_8660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8662 = 8'ha2 == r_count_41_io_out ? io_r_162_b : _GEN_8661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8663 = 8'ha3 == r_count_41_io_out ? io_r_163_b : _GEN_8662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8664 = 8'ha4 == r_count_41_io_out ? io_r_164_b : _GEN_8663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8665 = 8'ha5 == r_count_41_io_out ? io_r_165_b : _GEN_8664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8666 = 8'ha6 == r_count_41_io_out ? io_r_166_b : _GEN_8665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8667 = 8'ha7 == r_count_41_io_out ? io_r_167_b : _GEN_8666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8668 = 8'ha8 == r_count_41_io_out ? io_r_168_b : _GEN_8667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8669 = 8'ha9 == r_count_41_io_out ? io_r_169_b : _GEN_8668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8670 = 8'haa == r_count_41_io_out ? io_r_170_b : _GEN_8669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8671 = 8'hab == r_count_41_io_out ? io_r_171_b : _GEN_8670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8672 = 8'hac == r_count_41_io_out ? io_r_172_b : _GEN_8671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8673 = 8'had == r_count_41_io_out ? io_r_173_b : _GEN_8672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8674 = 8'hae == r_count_41_io_out ? io_r_174_b : _GEN_8673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8675 = 8'haf == r_count_41_io_out ? io_r_175_b : _GEN_8674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8676 = 8'hb0 == r_count_41_io_out ? io_r_176_b : _GEN_8675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8677 = 8'hb1 == r_count_41_io_out ? io_r_177_b : _GEN_8676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8678 = 8'hb2 == r_count_41_io_out ? io_r_178_b : _GEN_8677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8679 = 8'hb3 == r_count_41_io_out ? io_r_179_b : _GEN_8678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8680 = 8'hb4 == r_count_41_io_out ? io_r_180_b : _GEN_8679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8681 = 8'hb5 == r_count_41_io_out ? io_r_181_b : _GEN_8680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8682 = 8'hb6 == r_count_41_io_out ? io_r_182_b : _GEN_8681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8683 = 8'hb7 == r_count_41_io_out ? io_r_183_b : _GEN_8682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8684 = 8'hb8 == r_count_41_io_out ? io_r_184_b : _GEN_8683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8685 = 8'hb9 == r_count_41_io_out ? io_r_185_b : _GEN_8684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8686 = 8'hba == r_count_41_io_out ? io_r_186_b : _GEN_8685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8687 = 8'hbb == r_count_41_io_out ? io_r_187_b : _GEN_8686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8688 = 8'hbc == r_count_41_io_out ? io_r_188_b : _GEN_8687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8689 = 8'hbd == r_count_41_io_out ? io_r_189_b : _GEN_8688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8690 = 8'hbe == r_count_41_io_out ? io_r_190_b : _GEN_8689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8691 = 8'hbf == r_count_41_io_out ? io_r_191_b : _GEN_8690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8692 = 8'hc0 == r_count_41_io_out ? io_r_192_b : _GEN_8691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8693 = 8'hc1 == r_count_41_io_out ? io_r_193_b : _GEN_8692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8694 = 8'hc2 == r_count_41_io_out ? io_r_194_b : _GEN_8693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8695 = 8'hc3 == r_count_41_io_out ? io_r_195_b : _GEN_8694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8696 = 8'hc4 == r_count_41_io_out ? io_r_196_b : _GEN_8695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8697 = 8'hc5 == r_count_41_io_out ? io_r_197_b : _GEN_8696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8698 = 8'hc6 == r_count_41_io_out ? io_r_198_b : _GEN_8697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8701 = 8'h1 == r_count_42_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8702 = 8'h2 == r_count_42_io_out ? io_r_2_b : _GEN_8701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8703 = 8'h3 == r_count_42_io_out ? io_r_3_b : _GEN_8702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8704 = 8'h4 == r_count_42_io_out ? io_r_4_b : _GEN_8703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8705 = 8'h5 == r_count_42_io_out ? io_r_5_b : _GEN_8704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8706 = 8'h6 == r_count_42_io_out ? io_r_6_b : _GEN_8705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8707 = 8'h7 == r_count_42_io_out ? io_r_7_b : _GEN_8706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8708 = 8'h8 == r_count_42_io_out ? io_r_8_b : _GEN_8707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8709 = 8'h9 == r_count_42_io_out ? io_r_9_b : _GEN_8708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8710 = 8'ha == r_count_42_io_out ? io_r_10_b : _GEN_8709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8711 = 8'hb == r_count_42_io_out ? io_r_11_b : _GEN_8710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8712 = 8'hc == r_count_42_io_out ? io_r_12_b : _GEN_8711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8713 = 8'hd == r_count_42_io_out ? io_r_13_b : _GEN_8712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8714 = 8'he == r_count_42_io_out ? io_r_14_b : _GEN_8713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8715 = 8'hf == r_count_42_io_out ? io_r_15_b : _GEN_8714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8716 = 8'h10 == r_count_42_io_out ? io_r_16_b : _GEN_8715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8717 = 8'h11 == r_count_42_io_out ? io_r_17_b : _GEN_8716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8718 = 8'h12 == r_count_42_io_out ? io_r_18_b : _GEN_8717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8719 = 8'h13 == r_count_42_io_out ? io_r_19_b : _GEN_8718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8720 = 8'h14 == r_count_42_io_out ? io_r_20_b : _GEN_8719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8721 = 8'h15 == r_count_42_io_out ? io_r_21_b : _GEN_8720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8722 = 8'h16 == r_count_42_io_out ? io_r_22_b : _GEN_8721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8723 = 8'h17 == r_count_42_io_out ? io_r_23_b : _GEN_8722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8724 = 8'h18 == r_count_42_io_out ? io_r_24_b : _GEN_8723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8725 = 8'h19 == r_count_42_io_out ? io_r_25_b : _GEN_8724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8726 = 8'h1a == r_count_42_io_out ? io_r_26_b : _GEN_8725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8727 = 8'h1b == r_count_42_io_out ? io_r_27_b : _GEN_8726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8728 = 8'h1c == r_count_42_io_out ? io_r_28_b : _GEN_8727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8729 = 8'h1d == r_count_42_io_out ? io_r_29_b : _GEN_8728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8730 = 8'h1e == r_count_42_io_out ? io_r_30_b : _GEN_8729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8731 = 8'h1f == r_count_42_io_out ? io_r_31_b : _GEN_8730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8732 = 8'h20 == r_count_42_io_out ? io_r_32_b : _GEN_8731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8733 = 8'h21 == r_count_42_io_out ? io_r_33_b : _GEN_8732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8734 = 8'h22 == r_count_42_io_out ? io_r_34_b : _GEN_8733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8735 = 8'h23 == r_count_42_io_out ? io_r_35_b : _GEN_8734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8736 = 8'h24 == r_count_42_io_out ? io_r_36_b : _GEN_8735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8737 = 8'h25 == r_count_42_io_out ? io_r_37_b : _GEN_8736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8738 = 8'h26 == r_count_42_io_out ? io_r_38_b : _GEN_8737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8739 = 8'h27 == r_count_42_io_out ? io_r_39_b : _GEN_8738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8740 = 8'h28 == r_count_42_io_out ? io_r_40_b : _GEN_8739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8741 = 8'h29 == r_count_42_io_out ? io_r_41_b : _GEN_8740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8742 = 8'h2a == r_count_42_io_out ? io_r_42_b : _GEN_8741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8743 = 8'h2b == r_count_42_io_out ? io_r_43_b : _GEN_8742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8744 = 8'h2c == r_count_42_io_out ? io_r_44_b : _GEN_8743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8745 = 8'h2d == r_count_42_io_out ? io_r_45_b : _GEN_8744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8746 = 8'h2e == r_count_42_io_out ? io_r_46_b : _GEN_8745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8747 = 8'h2f == r_count_42_io_out ? io_r_47_b : _GEN_8746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8748 = 8'h30 == r_count_42_io_out ? io_r_48_b : _GEN_8747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8749 = 8'h31 == r_count_42_io_out ? io_r_49_b : _GEN_8748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8750 = 8'h32 == r_count_42_io_out ? io_r_50_b : _GEN_8749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8751 = 8'h33 == r_count_42_io_out ? io_r_51_b : _GEN_8750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8752 = 8'h34 == r_count_42_io_out ? io_r_52_b : _GEN_8751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8753 = 8'h35 == r_count_42_io_out ? io_r_53_b : _GEN_8752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8754 = 8'h36 == r_count_42_io_out ? io_r_54_b : _GEN_8753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8755 = 8'h37 == r_count_42_io_out ? io_r_55_b : _GEN_8754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8756 = 8'h38 == r_count_42_io_out ? io_r_56_b : _GEN_8755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8757 = 8'h39 == r_count_42_io_out ? io_r_57_b : _GEN_8756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8758 = 8'h3a == r_count_42_io_out ? io_r_58_b : _GEN_8757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8759 = 8'h3b == r_count_42_io_out ? io_r_59_b : _GEN_8758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8760 = 8'h3c == r_count_42_io_out ? io_r_60_b : _GEN_8759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8761 = 8'h3d == r_count_42_io_out ? io_r_61_b : _GEN_8760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8762 = 8'h3e == r_count_42_io_out ? io_r_62_b : _GEN_8761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8763 = 8'h3f == r_count_42_io_out ? io_r_63_b : _GEN_8762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8764 = 8'h40 == r_count_42_io_out ? io_r_64_b : _GEN_8763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8765 = 8'h41 == r_count_42_io_out ? io_r_65_b : _GEN_8764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8766 = 8'h42 == r_count_42_io_out ? io_r_66_b : _GEN_8765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8767 = 8'h43 == r_count_42_io_out ? io_r_67_b : _GEN_8766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8768 = 8'h44 == r_count_42_io_out ? io_r_68_b : _GEN_8767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8769 = 8'h45 == r_count_42_io_out ? io_r_69_b : _GEN_8768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8770 = 8'h46 == r_count_42_io_out ? io_r_70_b : _GEN_8769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8771 = 8'h47 == r_count_42_io_out ? io_r_71_b : _GEN_8770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8772 = 8'h48 == r_count_42_io_out ? io_r_72_b : _GEN_8771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8773 = 8'h49 == r_count_42_io_out ? io_r_73_b : _GEN_8772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8774 = 8'h4a == r_count_42_io_out ? io_r_74_b : _GEN_8773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8775 = 8'h4b == r_count_42_io_out ? io_r_75_b : _GEN_8774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8776 = 8'h4c == r_count_42_io_out ? io_r_76_b : _GEN_8775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8777 = 8'h4d == r_count_42_io_out ? io_r_77_b : _GEN_8776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8778 = 8'h4e == r_count_42_io_out ? io_r_78_b : _GEN_8777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8779 = 8'h4f == r_count_42_io_out ? io_r_79_b : _GEN_8778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8780 = 8'h50 == r_count_42_io_out ? io_r_80_b : _GEN_8779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8781 = 8'h51 == r_count_42_io_out ? io_r_81_b : _GEN_8780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8782 = 8'h52 == r_count_42_io_out ? io_r_82_b : _GEN_8781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8783 = 8'h53 == r_count_42_io_out ? io_r_83_b : _GEN_8782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8784 = 8'h54 == r_count_42_io_out ? io_r_84_b : _GEN_8783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8785 = 8'h55 == r_count_42_io_out ? io_r_85_b : _GEN_8784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8786 = 8'h56 == r_count_42_io_out ? io_r_86_b : _GEN_8785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8787 = 8'h57 == r_count_42_io_out ? io_r_87_b : _GEN_8786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8788 = 8'h58 == r_count_42_io_out ? io_r_88_b : _GEN_8787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8789 = 8'h59 == r_count_42_io_out ? io_r_89_b : _GEN_8788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8790 = 8'h5a == r_count_42_io_out ? io_r_90_b : _GEN_8789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8791 = 8'h5b == r_count_42_io_out ? io_r_91_b : _GEN_8790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8792 = 8'h5c == r_count_42_io_out ? io_r_92_b : _GEN_8791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8793 = 8'h5d == r_count_42_io_out ? io_r_93_b : _GEN_8792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8794 = 8'h5e == r_count_42_io_out ? io_r_94_b : _GEN_8793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8795 = 8'h5f == r_count_42_io_out ? io_r_95_b : _GEN_8794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8796 = 8'h60 == r_count_42_io_out ? io_r_96_b : _GEN_8795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8797 = 8'h61 == r_count_42_io_out ? io_r_97_b : _GEN_8796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8798 = 8'h62 == r_count_42_io_out ? io_r_98_b : _GEN_8797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8799 = 8'h63 == r_count_42_io_out ? io_r_99_b : _GEN_8798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8800 = 8'h64 == r_count_42_io_out ? io_r_100_b : _GEN_8799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8801 = 8'h65 == r_count_42_io_out ? io_r_101_b : _GEN_8800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8802 = 8'h66 == r_count_42_io_out ? io_r_102_b : _GEN_8801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8803 = 8'h67 == r_count_42_io_out ? io_r_103_b : _GEN_8802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8804 = 8'h68 == r_count_42_io_out ? io_r_104_b : _GEN_8803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8805 = 8'h69 == r_count_42_io_out ? io_r_105_b : _GEN_8804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8806 = 8'h6a == r_count_42_io_out ? io_r_106_b : _GEN_8805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8807 = 8'h6b == r_count_42_io_out ? io_r_107_b : _GEN_8806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8808 = 8'h6c == r_count_42_io_out ? io_r_108_b : _GEN_8807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8809 = 8'h6d == r_count_42_io_out ? io_r_109_b : _GEN_8808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8810 = 8'h6e == r_count_42_io_out ? io_r_110_b : _GEN_8809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8811 = 8'h6f == r_count_42_io_out ? io_r_111_b : _GEN_8810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8812 = 8'h70 == r_count_42_io_out ? io_r_112_b : _GEN_8811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8813 = 8'h71 == r_count_42_io_out ? io_r_113_b : _GEN_8812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8814 = 8'h72 == r_count_42_io_out ? io_r_114_b : _GEN_8813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8815 = 8'h73 == r_count_42_io_out ? io_r_115_b : _GEN_8814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8816 = 8'h74 == r_count_42_io_out ? io_r_116_b : _GEN_8815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8817 = 8'h75 == r_count_42_io_out ? io_r_117_b : _GEN_8816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8818 = 8'h76 == r_count_42_io_out ? io_r_118_b : _GEN_8817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8819 = 8'h77 == r_count_42_io_out ? io_r_119_b : _GEN_8818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8820 = 8'h78 == r_count_42_io_out ? io_r_120_b : _GEN_8819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8821 = 8'h79 == r_count_42_io_out ? io_r_121_b : _GEN_8820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8822 = 8'h7a == r_count_42_io_out ? io_r_122_b : _GEN_8821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8823 = 8'h7b == r_count_42_io_out ? io_r_123_b : _GEN_8822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8824 = 8'h7c == r_count_42_io_out ? io_r_124_b : _GEN_8823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8825 = 8'h7d == r_count_42_io_out ? io_r_125_b : _GEN_8824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8826 = 8'h7e == r_count_42_io_out ? io_r_126_b : _GEN_8825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8827 = 8'h7f == r_count_42_io_out ? io_r_127_b : _GEN_8826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8828 = 8'h80 == r_count_42_io_out ? io_r_128_b : _GEN_8827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8829 = 8'h81 == r_count_42_io_out ? io_r_129_b : _GEN_8828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8830 = 8'h82 == r_count_42_io_out ? io_r_130_b : _GEN_8829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8831 = 8'h83 == r_count_42_io_out ? io_r_131_b : _GEN_8830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8832 = 8'h84 == r_count_42_io_out ? io_r_132_b : _GEN_8831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8833 = 8'h85 == r_count_42_io_out ? io_r_133_b : _GEN_8832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8834 = 8'h86 == r_count_42_io_out ? io_r_134_b : _GEN_8833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8835 = 8'h87 == r_count_42_io_out ? io_r_135_b : _GEN_8834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8836 = 8'h88 == r_count_42_io_out ? io_r_136_b : _GEN_8835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8837 = 8'h89 == r_count_42_io_out ? io_r_137_b : _GEN_8836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8838 = 8'h8a == r_count_42_io_out ? io_r_138_b : _GEN_8837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8839 = 8'h8b == r_count_42_io_out ? io_r_139_b : _GEN_8838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8840 = 8'h8c == r_count_42_io_out ? io_r_140_b : _GEN_8839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8841 = 8'h8d == r_count_42_io_out ? io_r_141_b : _GEN_8840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8842 = 8'h8e == r_count_42_io_out ? io_r_142_b : _GEN_8841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8843 = 8'h8f == r_count_42_io_out ? io_r_143_b : _GEN_8842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8844 = 8'h90 == r_count_42_io_out ? io_r_144_b : _GEN_8843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8845 = 8'h91 == r_count_42_io_out ? io_r_145_b : _GEN_8844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8846 = 8'h92 == r_count_42_io_out ? io_r_146_b : _GEN_8845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8847 = 8'h93 == r_count_42_io_out ? io_r_147_b : _GEN_8846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8848 = 8'h94 == r_count_42_io_out ? io_r_148_b : _GEN_8847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8849 = 8'h95 == r_count_42_io_out ? io_r_149_b : _GEN_8848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8850 = 8'h96 == r_count_42_io_out ? io_r_150_b : _GEN_8849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8851 = 8'h97 == r_count_42_io_out ? io_r_151_b : _GEN_8850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8852 = 8'h98 == r_count_42_io_out ? io_r_152_b : _GEN_8851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8853 = 8'h99 == r_count_42_io_out ? io_r_153_b : _GEN_8852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8854 = 8'h9a == r_count_42_io_out ? io_r_154_b : _GEN_8853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8855 = 8'h9b == r_count_42_io_out ? io_r_155_b : _GEN_8854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8856 = 8'h9c == r_count_42_io_out ? io_r_156_b : _GEN_8855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8857 = 8'h9d == r_count_42_io_out ? io_r_157_b : _GEN_8856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8858 = 8'h9e == r_count_42_io_out ? io_r_158_b : _GEN_8857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8859 = 8'h9f == r_count_42_io_out ? io_r_159_b : _GEN_8858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8860 = 8'ha0 == r_count_42_io_out ? io_r_160_b : _GEN_8859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8861 = 8'ha1 == r_count_42_io_out ? io_r_161_b : _GEN_8860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8862 = 8'ha2 == r_count_42_io_out ? io_r_162_b : _GEN_8861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8863 = 8'ha3 == r_count_42_io_out ? io_r_163_b : _GEN_8862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8864 = 8'ha4 == r_count_42_io_out ? io_r_164_b : _GEN_8863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8865 = 8'ha5 == r_count_42_io_out ? io_r_165_b : _GEN_8864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8866 = 8'ha6 == r_count_42_io_out ? io_r_166_b : _GEN_8865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8867 = 8'ha7 == r_count_42_io_out ? io_r_167_b : _GEN_8866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8868 = 8'ha8 == r_count_42_io_out ? io_r_168_b : _GEN_8867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8869 = 8'ha9 == r_count_42_io_out ? io_r_169_b : _GEN_8868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8870 = 8'haa == r_count_42_io_out ? io_r_170_b : _GEN_8869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8871 = 8'hab == r_count_42_io_out ? io_r_171_b : _GEN_8870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8872 = 8'hac == r_count_42_io_out ? io_r_172_b : _GEN_8871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8873 = 8'had == r_count_42_io_out ? io_r_173_b : _GEN_8872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8874 = 8'hae == r_count_42_io_out ? io_r_174_b : _GEN_8873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8875 = 8'haf == r_count_42_io_out ? io_r_175_b : _GEN_8874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8876 = 8'hb0 == r_count_42_io_out ? io_r_176_b : _GEN_8875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8877 = 8'hb1 == r_count_42_io_out ? io_r_177_b : _GEN_8876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8878 = 8'hb2 == r_count_42_io_out ? io_r_178_b : _GEN_8877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8879 = 8'hb3 == r_count_42_io_out ? io_r_179_b : _GEN_8878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8880 = 8'hb4 == r_count_42_io_out ? io_r_180_b : _GEN_8879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8881 = 8'hb5 == r_count_42_io_out ? io_r_181_b : _GEN_8880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8882 = 8'hb6 == r_count_42_io_out ? io_r_182_b : _GEN_8881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8883 = 8'hb7 == r_count_42_io_out ? io_r_183_b : _GEN_8882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8884 = 8'hb8 == r_count_42_io_out ? io_r_184_b : _GEN_8883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8885 = 8'hb9 == r_count_42_io_out ? io_r_185_b : _GEN_8884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8886 = 8'hba == r_count_42_io_out ? io_r_186_b : _GEN_8885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8887 = 8'hbb == r_count_42_io_out ? io_r_187_b : _GEN_8886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8888 = 8'hbc == r_count_42_io_out ? io_r_188_b : _GEN_8887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8889 = 8'hbd == r_count_42_io_out ? io_r_189_b : _GEN_8888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8890 = 8'hbe == r_count_42_io_out ? io_r_190_b : _GEN_8889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8891 = 8'hbf == r_count_42_io_out ? io_r_191_b : _GEN_8890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8892 = 8'hc0 == r_count_42_io_out ? io_r_192_b : _GEN_8891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8893 = 8'hc1 == r_count_42_io_out ? io_r_193_b : _GEN_8892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8894 = 8'hc2 == r_count_42_io_out ? io_r_194_b : _GEN_8893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8895 = 8'hc3 == r_count_42_io_out ? io_r_195_b : _GEN_8894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8896 = 8'hc4 == r_count_42_io_out ? io_r_196_b : _GEN_8895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8897 = 8'hc5 == r_count_42_io_out ? io_r_197_b : _GEN_8896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8898 = 8'hc6 == r_count_42_io_out ? io_r_198_b : _GEN_8897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8901 = 8'h1 == r_count_43_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8902 = 8'h2 == r_count_43_io_out ? io_r_2_b : _GEN_8901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8903 = 8'h3 == r_count_43_io_out ? io_r_3_b : _GEN_8902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8904 = 8'h4 == r_count_43_io_out ? io_r_4_b : _GEN_8903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8905 = 8'h5 == r_count_43_io_out ? io_r_5_b : _GEN_8904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8906 = 8'h6 == r_count_43_io_out ? io_r_6_b : _GEN_8905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8907 = 8'h7 == r_count_43_io_out ? io_r_7_b : _GEN_8906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8908 = 8'h8 == r_count_43_io_out ? io_r_8_b : _GEN_8907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8909 = 8'h9 == r_count_43_io_out ? io_r_9_b : _GEN_8908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8910 = 8'ha == r_count_43_io_out ? io_r_10_b : _GEN_8909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8911 = 8'hb == r_count_43_io_out ? io_r_11_b : _GEN_8910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8912 = 8'hc == r_count_43_io_out ? io_r_12_b : _GEN_8911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8913 = 8'hd == r_count_43_io_out ? io_r_13_b : _GEN_8912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8914 = 8'he == r_count_43_io_out ? io_r_14_b : _GEN_8913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8915 = 8'hf == r_count_43_io_out ? io_r_15_b : _GEN_8914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8916 = 8'h10 == r_count_43_io_out ? io_r_16_b : _GEN_8915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8917 = 8'h11 == r_count_43_io_out ? io_r_17_b : _GEN_8916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8918 = 8'h12 == r_count_43_io_out ? io_r_18_b : _GEN_8917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8919 = 8'h13 == r_count_43_io_out ? io_r_19_b : _GEN_8918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8920 = 8'h14 == r_count_43_io_out ? io_r_20_b : _GEN_8919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8921 = 8'h15 == r_count_43_io_out ? io_r_21_b : _GEN_8920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8922 = 8'h16 == r_count_43_io_out ? io_r_22_b : _GEN_8921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8923 = 8'h17 == r_count_43_io_out ? io_r_23_b : _GEN_8922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8924 = 8'h18 == r_count_43_io_out ? io_r_24_b : _GEN_8923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8925 = 8'h19 == r_count_43_io_out ? io_r_25_b : _GEN_8924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8926 = 8'h1a == r_count_43_io_out ? io_r_26_b : _GEN_8925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8927 = 8'h1b == r_count_43_io_out ? io_r_27_b : _GEN_8926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8928 = 8'h1c == r_count_43_io_out ? io_r_28_b : _GEN_8927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8929 = 8'h1d == r_count_43_io_out ? io_r_29_b : _GEN_8928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8930 = 8'h1e == r_count_43_io_out ? io_r_30_b : _GEN_8929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8931 = 8'h1f == r_count_43_io_out ? io_r_31_b : _GEN_8930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8932 = 8'h20 == r_count_43_io_out ? io_r_32_b : _GEN_8931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8933 = 8'h21 == r_count_43_io_out ? io_r_33_b : _GEN_8932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8934 = 8'h22 == r_count_43_io_out ? io_r_34_b : _GEN_8933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8935 = 8'h23 == r_count_43_io_out ? io_r_35_b : _GEN_8934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8936 = 8'h24 == r_count_43_io_out ? io_r_36_b : _GEN_8935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8937 = 8'h25 == r_count_43_io_out ? io_r_37_b : _GEN_8936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8938 = 8'h26 == r_count_43_io_out ? io_r_38_b : _GEN_8937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8939 = 8'h27 == r_count_43_io_out ? io_r_39_b : _GEN_8938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8940 = 8'h28 == r_count_43_io_out ? io_r_40_b : _GEN_8939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8941 = 8'h29 == r_count_43_io_out ? io_r_41_b : _GEN_8940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8942 = 8'h2a == r_count_43_io_out ? io_r_42_b : _GEN_8941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8943 = 8'h2b == r_count_43_io_out ? io_r_43_b : _GEN_8942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8944 = 8'h2c == r_count_43_io_out ? io_r_44_b : _GEN_8943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8945 = 8'h2d == r_count_43_io_out ? io_r_45_b : _GEN_8944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8946 = 8'h2e == r_count_43_io_out ? io_r_46_b : _GEN_8945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8947 = 8'h2f == r_count_43_io_out ? io_r_47_b : _GEN_8946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8948 = 8'h30 == r_count_43_io_out ? io_r_48_b : _GEN_8947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8949 = 8'h31 == r_count_43_io_out ? io_r_49_b : _GEN_8948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8950 = 8'h32 == r_count_43_io_out ? io_r_50_b : _GEN_8949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8951 = 8'h33 == r_count_43_io_out ? io_r_51_b : _GEN_8950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8952 = 8'h34 == r_count_43_io_out ? io_r_52_b : _GEN_8951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8953 = 8'h35 == r_count_43_io_out ? io_r_53_b : _GEN_8952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8954 = 8'h36 == r_count_43_io_out ? io_r_54_b : _GEN_8953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8955 = 8'h37 == r_count_43_io_out ? io_r_55_b : _GEN_8954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8956 = 8'h38 == r_count_43_io_out ? io_r_56_b : _GEN_8955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8957 = 8'h39 == r_count_43_io_out ? io_r_57_b : _GEN_8956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8958 = 8'h3a == r_count_43_io_out ? io_r_58_b : _GEN_8957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8959 = 8'h3b == r_count_43_io_out ? io_r_59_b : _GEN_8958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8960 = 8'h3c == r_count_43_io_out ? io_r_60_b : _GEN_8959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8961 = 8'h3d == r_count_43_io_out ? io_r_61_b : _GEN_8960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8962 = 8'h3e == r_count_43_io_out ? io_r_62_b : _GEN_8961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8963 = 8'h3f == r_count_43_io_out ? io_r_63_b : _GEN_8962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8964 = 8'h40 == r_count_43_io_out ? io_r_64_b : _GEN_8963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8965 = 8'h41 == r_count_43_io_out ? io_r_65_b : _GEN_8964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8966 = 8'h42 == r_count_43_io_out ? io_r_66_b : _GEN_8965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8967 = 8'h43 == r_count_43_io_out ? io_r_67_b : _GEN_8966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8968 = 8'h44 == r_count_43_io_out ? io_r_68_b : _GEN_8967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8969 = 8'h45 == r_count_43_io_out ? io_r_69_b : _GEN_8968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8970 = 8'h46 == r_count_43_io_out ? io_r_70_b : _GEN_8969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8971 = 8'h47 == r_count_43_io_out ? io_r_71_b : _GEN_8970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8972 = 8'h48 == r_count_43_io_out ? io_r_72_b : _GEN_8971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8973 = 8'h49 == r_count_43_io_out ? io_r_73_b : _GEN_8972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8974 = 8'h4a == r_count_43_io_out ? io_r_74_b : _GEN_8973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8975 = 8'h4b == r_count_43_io_out ? io_r_75_b : _GEN_8974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8976 = 8'h4c == r_count_43_io_out ? io_r_76_b : _GEN_8975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8977 = 8'h4d == r_count_43_io_out ? io_r_77_b : _GEN_8976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8978 = 8'h4e == r_count_43_io_out ? io_r_78_b : _GEN_8977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8979 = 8'h4f == r_count_43_io_out ? io_r_79_b : _GEN_8978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8980 = 8'h50 == r_count_43_io_out ? io_r_80_b : _GEN_8979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8981 = 8'h51 == r_count_43_io_out ? io_r_81_b : _GEN_8980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8982 = 8'h52 == r_count_43_io_out ? io_r_82_b : _GEN_8981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8983 = 8'h53 == r_count_43_io_out ? io_r_83_b : _GEN_8982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8984 = 8'h54 == r_count_43_io_out ? io_r_84_b : _GEN_8983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8985 = 8'h55 == r_count_43_io_out ? io_r_85_b : _GEN_8984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8986 = 8'h56 == r_count_43_io_out ? io_r_86_b : _GEN_8985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8987 = 8'h57 == r_count_43_io_out ? io_r_87_b : _GEN_8986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8988 = 8'h58 == r_count_43_io_out ? io_r_88_b : _GEN_8987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8989 = 8'h59 == r_count_43_io_out ? io_r_89_b : _GEN_8988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8990 = 8'h5a == r_count_43_io_out ? io_r_90_b : _GEN_8989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8991 = 8'h5b == r_count_43_io_out ? io_r_91_b : _GEN_8990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8992 = 8'h5c == r_count_43_io_out ? io_r_92_b : _GEN_8991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8993 = 8'h5d == r_count_43_io_out ? io_r_93_b : _GEN_8992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8994 = 8'h5e == r_count_43_io_out ? io_r_94_b : _GEN_8993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8995 = 8'h5f == r_count_43_io_out ? io_r_95_b : _GEN_8994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8996 = 8'h60 == r_count_43_io_out ? io_r_96_b : _GEN_8995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8997 = 8'h61 == r_count_43_io_out ? io_r_97_b : _GEN_8996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8998 = 8'h62 == r_count_43_io_out ? io_r_98_b : _GEN_8997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8999 = 8'h63 == r_count_43_io_out ? io_r_99_b : _GEN_8998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9000 = 8'h64 == r_count_43_io_out ? io_r_100_b : _GEN_8999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9001 = 8'h65 == r_count_43_io_out ? io_r_101_b : _GEN_9000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9002 = 8'h66 == r_count_43_io_out ? io_r_102_b : _GEN_9001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9003 = 8'h67 == r_count_43_io_out ? io_r_103_b : _GEN_9002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9004 = 8'h68 == r_count_43_io_out ? io_r_104_b : _GEN_9003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9005 = 8'h69 == r_count_43_io_out ? io_r_105_b : _GEN_9004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9006 = 8'h6a == r_count_43_io_out ? io_r_106_b : _GEN_9005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9007 = 8'h6b == r_count_43_io_out ? io_r_107_b : _GEN_9006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9008 = 8'h6c == r_count_43_io_out ? io_r_108_b : _GEN_9007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9009 = 8'h6d == r_count_43_io_out ? io_r_109_b : _GEN_9008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9010 = 8'h6e == r_count_43_io_out ? io_r_110_b : _GEN_9009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9011 = 8'h6f == r_count_43_io_out ? io_r_111_b : _GEN_9010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9012 = 8'h70 == r_count_43_io_out ? io_r_112_b : _GEN_9011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9013 = 8'h71 == r_count_43_io_out ? io_r_113_b : _GEN_9012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9014 = 8'h72 == r_count_43_io_out ? io_r_114_b : _GEN_9013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9015 = 8'h73 == r_count_43_io_out ? io_r_115_b : _GEN_9014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9016 = 8'h74 == r_count_43_io_out ? io_r_116_b : _GEN_9015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9017 = 8'h75 == r_count_43_io_out ? io_r_117_b : _GEN_9016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9018 = 8'h76 == r_count_43_io_out ? io_r_118_b : _GEN_9017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9019 = 8'h77 == r_count_43_io_out ? io_r_119_b : _GEN_9018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9020 = 8'h78 == r_count_43_io_out ? io_r_120_b : _GEN_9019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9021 = 8'h79 == r_count_43_io_out ? io_r_121_b : _GEN_9020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9022 = 8'h7a == r_count_43_io_out ? io_r_122_b : _GEN_9021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9023 = 8'h7b == r_count_43_io_out ? io_r_123_b : _GEN_9022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9024 = 8'h7c == r_count_43_io_out ? io_r_124_b : _GEN_9023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9025 = 8'h7d == r_count_43_io_out ? io_r_125_b : _GEN_9024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9026 = 8'h7e == r_count_43_io_out ? io_r_126_b : _GEN_9025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9027 = 8'h7f == r_count_43_io_out ? io_r_127_b : _GEN_9026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9028 = 8'h80 == r_count_43_io_out ? io_r_128_b : _GEN_9027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9029 = 8'h81 == r_count_43_io_out ? io_r_129_b : _GEN_9028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9030 = 8'h82 == r_count_43_io_out ? io_r_130_b : _GEN_9029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9031 = 8'h83 == r_count_43_io_out ? io_r_131_b : _GEN_9030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9032 = 8'h84 == r_count_43_io_out ? io_r_132_b : _GEN_9031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9033 = 8'h85 == r_count_43_io_out ? io_r_133_b : _GEN_9032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9034 = 8'h86 == r_count_43_io_out ? io_r_134_b : _GEN_9033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9035 = 8'h87 == r_count_43_io_out ? io_r_135_b : _GEN_9034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9036 = 8'h88 == r_count_43_io_out ? io_r_136_b : _GEN_9035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9037 = 8'h89 == r_count_43_io_out ? io_r_137_b : _GEN_9036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9038 = 8'h8a == r_count_43_io_out ? io_r_138_b : _GEN_9037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9039 = 8'h8b == r_count_43_io_out ? io_r_139_b : _GEN_9038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9040 = 8'h8c == r_count_43_io_out ? io_r_140_b : _GEN_9039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9041 = 8'h8d == r_count_43_io_out ? io_r_141_b : _GEN_9040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9042 = 8'h8e == r_count_43_io_out ? io_r_142_b : _GEN_9041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9043 = 8'h8f == r_count_43_io_out ? io_r_143_b : _GEN_9042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9044 = 8'h90 == r_count_43_io_out ? io_r_144_b : _GEN_9043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9045 = 8'h91 == r_count_43_io_out ? io_r_145_b : _GEN_9044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9046 = 8'h92 == r_count_43_io_out ? io_r_146_b : _GEN_9045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9047 = 8'h93 == r_count_43_io_out ? io_r_147_b : _GEN_9046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9048 = 8'h94 == r_count_43_io_out ? io_r_148_b : _GEN_9047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9049 = 8'h95 == r_count_43_io_out ? io_r_149_b : _GEN_9048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9050 = 8'h96 == r_count_43_io_out ? io_r_150_b : _GEN_9049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9051 = 8'h97 == r_count_43_io_out ? io_r_151_b : _GEN_9050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9052 = 8'h98 == r_count_43_io_out ? io_r_152_b : _GEN_9051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9053 = 8'h99 == r_count_43_io_out ? io_r_153_b : _GEN_9052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9054 = 8'h9a == r_count_43_io_out ? io_r_154_b : _GEN_9053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9055 = 8'h9b == r_count_43_io_out ? io_r_155_b : _GEN_9054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9056 = 8'h9c == r_count_43_io_out ? io_r_156_b : _GEN_9055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9057 = 8'h9d == r_count_43_io_out ? io_r_157_b : _GEN_9056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9058 = 8'h9e == r_count_43_io_out ? io_r_158_b : _GEN_9057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9059 = 8'h9f == r_count_43_io_out ? io_r_159_b : _GEN_9058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9060 = 8'ha0 == r_count_43_io_out ? io_r_160_b : _GEN_9059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9061 = 8'ha1 == r_count_43_io_out ? io_r_161_b : _GEN_9060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9062 = 8'ha2 == r_count_43_io_out ? io_r_162_b : _GEN_9061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9063 = 8'ha3 == r_count_43_io_out ? io_r_163_b : _GEN_9062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9064 = 8'ha4 == r_count_43_io_out ? io_r_164_b : _GEN_9063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9065 = 8'ha5 == r_count_43_io_out ? io_r_165_b : _GEN_9064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9066 = 8'ha6 == r_count_43_io_out ? io_r_166_b : _GEN_9065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9067 = 8'ha7 == r_count_43_io_out ? io_r_167_b : _GEN_9066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9068 = 8'ha8 == r_count_43_io_out ? io_r_168_b : _GEN_9067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9069 = 8'ha9 == r_count_43_io_out ? io_r_169_b : _GEN_9068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9070 = 8'haa == r_count_43_io_out ? io_r_170_b : _GEN_9069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9071 = 8'hab == r_count_43_io_out ? io_r_171_b : _GEN_9070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9072 = 8'hac == r_count_43_io_out ? io_r_172_b : _GEN_9071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9073 = 8'had == r_count_43_io_out ? io_r_173_b : _GEN_9072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9074 = 8'hae == r_count_43_io_out ? io_r_174_b : _GEN_9073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9075 = 8'haf == r_count_43_io_out ? io_r_175_b : _GEN_9074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9076 = 8'hb0 == r_count_43_io_out ? io_r_176_b : _GEN_9075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9077 = 8'hb1 == r_count_43_io_out ? io_r_177_b : _GEN_9076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9078 = 8'hb2 == r_count_43_io_out ? io_r_178_b : _GEN_9077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9079 = 8'hb3 == r_count_43_io_out ? io_r_179_b : _GEN_9078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9080 = 8'hb4 == r_count_43_io_out ? io_r_180_b : _GEN_9079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9081 = 8'hb5 == r_count_43_io_out ? io_r_181_b : _GEN_9080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9082 = 8'hb6 == r_count_43_io_out ? io_r_182_b : _GEN_9081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9083 = 8'hb7 == r_count_43_io_out ? io_r_183_b : _GEN_9082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9084 = 8'hb8 == r_count_43_io_out ? io_r_184_b : _GEN_9083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9085 = 8'hb9 == r_count_43_io_out ? io_r_185_b : _GEN_9084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9086 = 8'hba == r_count_43_io_out ? io_r_186_b : _GEN_9085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9087 = 8'hbb == r_count_43_io_out ? io_r_187_b : _GEN_9086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9088 = 8'hbc == r_count_43_io_out ? io_r_188_b : _GEN_9087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9089 = 8'hbd == r_count_43_io_out ? io_r_189_b : _GEN_9088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9090 = 8'hbe == r_count_43_io_out ? io_r_190_b : _GEN_9089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9091 = 8'hbf == r_count_43_io_out ? io_r_191_b : _GEN_9090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9092 = 8'hc0 == r_count_43_io_out ? io_r_192_b : _GEN_9091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9093 = 8'hc1 == r_count_43_io_out ? io_r_193_b : _GEN_9092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9094 = 8'hc2 == r_count_43_io_out ? io_r_194_b : _GEN_9093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9095 = 8'hc3 == r_count_43_io_out ? io_r_195_b : _GEN_9094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9096 = 8'hc4 == r_count_43_io_out ? io_r_196_b : _GEN_9095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9097 = 8'hc5 == r_count_43_io_out ? io_r_197_b : _GEN_9096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9098 = 8'hc6 == r_count_43_io_out ? io_r_198_b : _GEN_9097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9101 = 8'h1 == r_count_44_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9102 = 8'h2 == r_count_44_io_out ? io_r_2_b : _GEN_9101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9103 = 8'h3 == r_count_44_io_out ? io_r_3_b : _GEN_9102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9104 = 8'h4 == r_count_44_io_out ? io_r_4_b : _GEN_9103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9105 = 8'h5 == r_count_44_io_out ? io_r_5_b : _GEN_9104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9106 = 8'h6 == r_count_44_io_out ? io_r_6_b : _GEN_9105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9107 = 8'h7 == r_count_44_io_out ? io_r_7_b : _GEN_9106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9108 = 8'h8 == r_count_44_io_out ? io_r_8_b : _GEN_9107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9109 = 8'h9 == r_count_44_io_out ? io_r_9_b : _GEN_9108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9110 = 8'ha == r_count_44_io_out ? io_r_10_b : _GEN_9109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9111 = 8'hb == r_count_44_io_out ? io_r_11_b : _GEN_9110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9112 = 8'hc == r_count_44_io_out ? io_r_12_b : _GEN_9111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9113 = 8'hd == r_count_44_io_out ? io_r_13_b : _GEN_9112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9114 = 8'he == r_count_44_io_out ? io_r_14_b : _GEN_9113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9115 = 8'hf == r_count_44_io_out ? io_r_15_b : _GEN_9114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9116 = 8'h10 == r_count_44_io_out ? io_r_16_b : _GEN_9115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9117 = 8'h11 == r_count_44_io_out ? io_r_17_b : _GEN_9116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9118 = 8'h12 == r_count_44_io_out ? io_r_18_b : _GEN_9117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9119 = 8'h13 == r_count_44_io_out ? io_r_19_b : _GEN_9118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9120 = 8'h14 == r_count_44_io_out ? io_r_20_b : _GEN_9119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9121 = 8'h15 == r_count_44_io_out ? io_r_21_b : _GEN_9120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9122 = 8'h16 == r_count_44_io_out ? io_r_22_b : _GEN_9121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9123 = 8'h17 == r_count_44_io_out ? io_r_23_b : _GEN_9122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9124 = 8'h18 == r_count_44_io_out ? io_r_24_b : _GEN_9123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9125 = 8'h19 == r_count_44_io_out ? io_r_25_b : _GEN_9124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9126 = 8'h1a == r_count_44_io_out ? io_r_26_b : _GEN_9125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9127 = 8'h1b == r_count_44_io_out ? io_r_27_b : _GEN_9126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9128 = 8'h1c == r_count_44_io_out ? io_r_28_b : _GEN_9127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9129 = 8'h1d == r_count_44_io_out ? io_r_29_b : _GEN_9128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9130 = 8'h1e == r_count_44_io_out ? io_r_30_b : _GEN_9129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9131 = 8'h1f == r_count_44_io_out ? io_r_31_b : _GEN_9130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9132 = 8'h20 == r_count_44_io_out ? io_r_32_b : _GEN_9131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9133 = 8'h21 == r_count_44_io_out ? io_r_33_b : _GEN_9132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9134 = 8'h22 == r_count_44_io_out ? io_r_34_b : _GEN_9133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9135 = 8'h23 == r_count_44_io_out ? io_r_35_b : _GEN_9134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9136 = 8'h24 == r_count_44_io_out ? io_r_36_b : _GEN_9135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9137 = 8'h25 == r_count_44_io_out ? io_r_37_b : _GEN_9136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9138 = 8'h26 == r_count_44_io_out ? io_r_38_b : _GEN_9137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9139 = 8'h27 == r_count_44_io_out ? io_r_39_b : _GEN_9138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9140 = 8'h28 == r_count_44_io_out ? io_r_40_b : _GEN_9139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9141 = 8'h29 == r_count_44_io_out ? io_r_41_b : _GEN_9140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9142 = 8'h2a == r_count_44_io_out ? io_r_42_b : _GEN_9141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9143 = 8'h2b == r_count_44_io_out ? io_r_43_b : _GEN_9142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9144 = 8'h2c == r_count_44_io_out ? io_r_44_b : _GEN_9143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9145 = 8'h2d == r_count_44_io_out ? io_r_45_b : _GEN_9144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9146 = 8'h2e == r_count_44_io_out ? io_r_46_b : _GEN_9145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9147 = 8'h2f == r_count_44_io_out ? io_r_47_b : _GEN_9146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9148 = 8'h30 == r_count_44_io_out ? io_r_48_b : _GEN_9147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9149 = 8'h31 == r_count_44_io_out ? io_r_49_b : _GEN_9148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9150 = 8'h32 == r_count_44_io_out ? io_r_50_b : _GEN_9149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9151 = 8'h33 == r_count_44_io_out ? io_r_51_b : _GEN_9150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9152 = 8'h34 == r_count_44_io_out ? io_r_52_b : _GEN_9151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9153 = 8'h35 == r_count_44_io_out ? io_r_53_b : _GEN_9152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9154 = 8'h36 == r_count_44_io_out ? io_r_54_b : _GEN_9153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9155 = 8'h37 == r_count_44_io_out ? io_r_55_b : _GEN_9154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9156 = 8'h38 == r_count_44_io_out ? io_r_56_b : _GEN_9155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9157 = 8'h39 == r_count_44_io_out ? io_r_57_b : _GEN_9156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9158 = 8'h3a == r_count_44_io_out ? io_r_58_b : _GEN_9157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9159 = 8'h3b == r_count_44_io_out ? io_r_59_b : _GEN_9158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9160 = 8'h3c == r_count_44_io_out ? io_r_60_b : _GEN_9159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9161 = 8'h3d == r_count_44_io_out ? io_r_61_b : _GEN_9160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9162 = 8'h3e == r_count_44_io_out ? io_r_62_b : _GEN_9161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9163 = 8'h3f == r_count_44_io_out ? io_r_63_b : _GEN_9162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9164 = 8'h40 == r_count_44_io_out ? io_r_64_b : _GEN_9163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9165 = 8'h41 == r_count_44_io_out ? io_r_65_b : _GEN_9164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9166 = 8'h42 == r_count_44_io_out ? io_r_66_b : _GEN_9165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9167 = 8'h43 == r_count_44_io_out ? io_r_67_b : _GEN_9166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9168 = 8'h44 == r_count_44_io_out ? io_r_68_b : _GEN_9167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9169 = 8'h45 == r_count_44_io_out ? io_r_69_b : _GEN_9168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9170 = 8'h46 == r_count_44_io_out ? io_r_70_b : _GEN_9169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9171 = 8'h47 == r_count_44_io_out ? io_r_71_b : _GEN_9170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9172 = 8'h48 == r_count_44_io_out ? io_r_72_b : _GEN_9171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9173 = 8'h49 == r_count_44_io_out ? io_r_73_b : _GEN_9172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9174 = 8'h4a == r_count_44_io_out ? io_r_74_b : _GEN_9173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9175 = 8'h4b == r_count_44_io_out ? io_r_75_b : _GEN_9174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9176 = 8'h4c == r_count_44_io_out ? io_r_76_b : _GEN_9175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9177 = 8'h4d == r_count_44_io_out ? io_r_77_b : _GEN_9176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9178 = 8'h4e == r_count_44_io_out ? io_r_78_b : _GEN_9177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9179 = 8'h4f == r_count_44_io_out ? io_r_79_b : _GEN_9178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9180 = 8'h50 == r_count_44_io_out ? io_r_80_b : _GEN_9179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9181 = 8'h51 == r_count_44_io_out ? io_r_81_b : _GEN_9180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9182 = 8'h52 == r_count_44_io_out ? io_r_82_b : _GEN_9181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9183 = 8'h53 == r_count_44_io_out ? io_r_83_b : _GEN_9182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9184 = 8'h54 == r_count_44_io_out ? io_r_84_b : _GEN_9183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9185 = 8'h55 == r_count_44_io_out ? io_r_85_b : _GEN_9184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9186 = 8'h56 == r_count_44_io_out ? io_r_86_b : _GEN_9185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9187 = 8'h57 == r_count_44_io_out ? io_r_87_b : _GEN_9186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9188 = 8'h58 == r_count_44_io_out ? io_r_88_b : _GEN_9187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9189 = 8'h59 == r_count_44_io_out ? io_r_89_b : _GEN_9188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9190 = 8'h5a == r_count_44_io_out ? io_r_90_b : _GEN_9189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9191 = 8'h5b == r_count_44_io_out ? io_r_91_b : _GEN_9190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9192 = 8'h5c == r_count_44_io_out ? io_r_92_b : _GEN_9191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9193 = 8'h5d == r_count_44_io_out ? io_r_93_b : _GEN_9192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9194 = 8'h5e == r_count_44_io_out ? io_r_94_b : _GEN_9193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9195 = 8'h5f == r_count_44_io_out ? io_r_95_b : _GEN_9194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9196 = 8'h60 == r_count_44_io_out ? io_r_96_b : _GEN_9195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9197 = 8'h61 == r_count_44_io_out ? io_r_97_b : _GEN_9196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9198 = 8'h62 == r_count_44_io_out ? io_r_98_b : _GEN_9197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9199 = 8'h63 == r_count_44_io_out ? io_r_99_b : _GEN_9198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9200 = 8'h64 == r_count_44_io_out ? io_r_100_b : _GEN_9199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9201 = 8'h65 == r_count_44_io_out ? io_r_101_b : _GEN_9200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9202 = 8'h66 == r_count_44_io_out ? io_r_102_b : _GEN_9201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9203 = 8'h67 == r_count_44_io_out ? io_r_103_b : _GEN_9202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9204 = 8'h68 == r_count_44_io_out ? io_r_104_b : _GEN_9203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9205 = 8'h69 == r_count_44_io_out ? io_r_105_b : _GEN_9204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9206 = 8'h6a == r_count_44_io_out ? io_r_106_b : _GEN_9205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9207 = 8'h6b == r_count_44_io_out ? io_r_107_b : _GEN_9206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9208 = 8'h6c == r_count_44_io_out ? io_r_108_b : _GEN_9207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9209 = 8'h6d == r_count_44_io_out ? io_r_109_b : _GEN_9208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9210 = 8'h6e == r_count_44_io_out ? io_r_110_b : _GEN_9209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9211 = 8'h6f == r_count_44_io_out ? io_r_111_b : _GEN_9210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9212 = 8'h70 == r_count_44_io_out ? io_r_112_b : _GEN_9211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9213 = 8'h71 == r_count_44_io_out ? io_r_113_b : _GEN_9212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9214 = 8'h72 == r_count_44_io_out ? io_r_114_b : _GEN_9213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9215 = 8'h73 == r_count_44_io_out ? io_r_115_b : _GEN_9214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9216 = 8'h74 == r_count_44_io_out ? io_r_116_b : _GEN_9215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9217 = 8'h75 == r_count_44_io_out ? io_r_117_b : _GEN_9216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9218 = 8'h76 == r_count_44_io_out ? io_r_118_b : _GEN_9217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9219 = 8'h77 == r_count_44_io_out ? io_r_119_b : _GEN_9218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9220 = 8'h78 == r_count_44_io_out ? io_r_120_b : _GEN_9219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9221 = 8'h79 == r_count_44_io_out ? io_r_121_b : _GEN_9220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9222 = 8'h7a == r_count_44_io_out ? io_r_122_b : _GEN_9221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9223 = 8'h7b == r_count_44_io_out ? io_r_123_b : _GEN_9222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9224 = 8'h7c == r_count_44_io_out ? io_r_124_b : _GEN_9223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9225 = 8'h7d == r_count_44_io_out ? io_r_125_b : _GEN_9224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9226 = 8'h7e == r_count_44_io_out ? io_r_126_b : _GEN_9225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9227 = 8'h7f == r_count_44_io_out ? io_r_127_b : _GEN_9226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9228 = 8'h80 == r_count_44_io_out ? io_r_128_b : _GEN_9227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9229 = 8'h81 == r_count_44_io_out ? io_r_129_b : _GEN_9228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9230 = 8'h82 == r_count_44_io_out ? io_r_130_b : _GEN_9229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9231 = 8'h83 == r_count_44_io_out ? io_r_131_b : _GEN_9230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9232 = 8'h84 == r_count_44_io_out ? io_r_132_b : _GEN_9231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9233 = 8'h85 == r_count_44_io_out ? io_r_133_b : _GEN_9232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9234 = 8'h86 == r_count_44_io_out ? io_r_134_b : _GEN_9233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9235 = 8'h87 == r_count_44_io_out ? io_r_135_b : _GEN_9234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9236 = 8'h88 == r_count_44_io_out ? io_r_136_b : _GEN_9235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9237 = 8'h89 == r_count_44_io_out ? io_r_137_b : _GEN_9236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9238 = 8'h8a == r_count_44_io_out ? io_r_138_b : _GEN_9237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9239 = 8'h8b == r_count_44_io_out ? io_r_139_b : _GEN_9238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9240 = 8'h8c == r_count_44_io_out ? io_r_140_b : _GEN_9239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9241 = 8'h8d == r_count_44_io_out ? io_r_141_b : _GEN_9240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9242 = 8'h8e == r_count_44_io_out ? io_r_142_b : _GEN_9241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9243 = 8'h8f == r_count_44_io_out ? io_r_143_b : _GEN_9242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9244 = 8'h90 == r_count_44_io_out ? io_r_144_b : _GEN_9243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9245 = 8'h91 == r_count_44_io_out ? io_r_145_b : _GEN_9244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9246 = 8'h92 == r_count_44_io_out ? io_r_146_b : _GEN_9245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9247 = 8'h93 == r_count_44_io_out ? io_r_147_b : _GEN_9246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9248 = 8'h94 == r_count_44_io_out ? io_r_148_b : _GEN_9247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9249 = 8'h95 == r_count_44_io_out ? io_r_149_b : _GEN_9248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9250 = 8'h96 == r_count_44_io_out ? io_r_150_b : _GEN_9249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9251 = 8'h97 == r_count_44_io_out ? io_r_151_b : _GEN_9250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9252 = 8'h98 == r_count_44_io_out ? io_r_152_b : _GEN_9251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9253 = 8'h99 == r_count_44_io_out ? io_r_153_b : _GEN_9252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9254 = 8'h9a == r_count_44_io_out ? io_r_154_b : _GEN_9253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9255 = 8'h9b == r_count_44_io_out ? io_r_155_b : _GEN_9254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9256 = 8'h9c == r_count_44_io_out ? io_r_156_b : _GEN_9255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9257 = 8'h9d == r_count_44_io_out ? io_r_157_b : _GEN_9256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9258 = 8'h9e == r_count_44_io_out ? io_r_158_b : _GEN_9257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9259 = 8'h9f == r_count_44_io_out ? io_r_159_b : _GEN_9258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9260 = 8'ha0 == r_count_44_io_out ? io_r_160_b : _GEN_9259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9261 = 8'ha1 == r_count_44_io_out ? io_r_161_b : _GEN_9260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9262 = 8'ha2 == r_count_44_io_out ? io_r_162_b : _GEN_9261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9263 = 8'ha3 == r_count_44_io_out ? io_r_163_b : _GEN_9262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9264 = 8'ha4 == r_count_44_io_out ? io_r_164_b : _GEN_9263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9265 = 8'ha5 == r_count_44_io_out ? io_r_165_b : _GEN_9264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9266 = 8'ha6 == r_count_44_io_out ? io_r_166_b : _GEN_9265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9267 = 8'ha7 == r_count_44_io_out ? io_r_167_b : _GEN_9266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9268 = 8'ha8 == r_count_44_io_out ? io_r_168_b : _GEN_9267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9269 = 8'ha9 == r_count_44_io_out ? io_r_169_b : _GEN_9268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9270 = 8'haa == r_count_44_io_out ? io_r_170_b : _GEN_9269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9271 = 8'hab == r_count_44_io_out ? io_r_171_b : _GEN_9270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9272 = 8'hac == r_count_44_io_out ? io_r_172_b : _GEN_9271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9273 = 8'had == r_count_44_io_out ? io_r_173_b : _GEN_9272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9274 = 8'hae == r_count_44_io_out ? io_r_174_b : _GEN_9273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9275 = 8'haf == r_count_44_io_out ? io_r_175_b : _GEN_9274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9276 = 8'hb0 == r_count_44_io_out ? io_r_176_b : _GEN_9275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9277 = 8'hb1 == r_count_44_io_out ? io_r_177_b : _GEN_9276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9278 = 8'hb2 == r_count_44_io_out ? io_r_178_b : _GEN_9277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9279 = 8'hb3 == r_count_44_io_out ? io_r_179_b : _GEN_9278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9280 = 8'hb4 == r_count_44_io_out ? io_r_180_b : _GEN_9279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9281 = 8'hb5 == r_count_44_io_out ? io_r_181_b : _GEN_9280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9282 = 8'hb6 == r_count_44_io_out ? io_r_182_b : _GEN_9281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9283 = 8'hb7 == r_count_44_io_out ? io_r_183_b : _GEN_9282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9284 = 8'hb8 == r_count_44_io_out ? io_r_184_b : _GEN_9283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9285 = 8'hb9 == r_count_44_io_out ? io_r_185_b : _GEN_9284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9286 = 8'hba == r_count_44_io_out ? io_r_186_b : _GEN_9285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9287 = 8'hbb == r_count_44_io_out ? io_r_187_b : _GEN_9286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9288 = 8'hbc == r_count_44_io_out ? io_r_188_b : _GEN_9287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9289 = 8'hbd == r_count_44_io_out ? io_r_189_b : _GEN_9288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9290 = 8'hbe == r_count_44_io_out ? io_r_190_b : _GEN_9289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9291 = 8'hbf == r_count_44_io_out ? io_r_191_b : _GEN_9290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9292 = 8'hc0 == r_count_44_io_out ? io_r_192_b : _GEN_9291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9293 = 8'hc1 == r_count_44_io_out ? io_r_193_b : _GEN_9292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9294 = 8'hc2 == r_count_44_io_out ? io_r_194_b : _GEN_9293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9295 = 8'hc3 == r_count_44_io_out ? io_r_195_b : _GEN_9294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9296 = 8'hc4 == r_count_44_io_out ? io_r_196_b : _GEN_9295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9297 = 8'hc5 == r_count_44_io_out ? io_r_197_b : _GEN_9296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9298 = 8'hc6 == r_count_44_io_out ? io_r_198_b : _GEN_9297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9301 = 8'h1 == r_count_45_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9302 = 8'h2 == r_count_45_io_out ? io_r_2_b : _GEN_9301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9303 = 8'h3 == r_count_45_io_out ? io_r_3_b : _GEN_9302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9304 = 8'h4 == r_count_45_io_out ? io_r_4_b : _GEN_9303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9305 = 8'h5 == r_count_45_io_out ? io_r_5_b : _GEN_9304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9306 = 8'h6 == r_count_45_io_out ? io_r_6_b : _GEN_9305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9307 = 8'h7 == r_count_45_io_out ? io_r_7_b : _GEN_9306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9308 = 8'h8 == r_count_45_io_out ? io_r_8_b : _GEN_9307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9309 = 8'h9 == r_count_45_io_out ? io_r_9_b : _GEN_9308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9310 = 8'ha == r_count_45_io_out ? io_r_10_b : _GEN_9309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9311 = 8'hb == r_count_45_io_out ? io_r_11_b : _GEN_9310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9312 = 8'hc == r_count_45_io_out ? io_r_12_b : _GEN_9311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9313 = 8'hd == r_count_45_io_out ? io_r_13_b : _GEN_9312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9314 = 8'he == r_count_45_io_out ? io_r_14_b : _GEN_9313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9315 = 8'hf == r_count_45_io_out ? io_r_15_b : _GEN_9314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9316 = 8'h10 == r_count_45_io_out ? io_r_16_b : _GEN_9315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9317 = 8'h11 == r_count_45_io_out ? io_r_17_b : _GEN_9316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9318 = 8'h12 == r_count_45_io_out ? io_r_18_b : _GEN_9317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9319 = 8'h13 == r_count_45_io_out ? io_r_19_b : _GEN_9318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9320 = 8'h14 == r_count_45_io_out ? io_r_20_b : _GEN_9319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9321 = 8'h15 == r_count_45_io_out ? io_r_21_b : _GEN_9320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9322 = 8'h16 == r_count_45_io_out ? io_r_22_b : _GEN_9321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9323 = 8'h17 == r_count_45_io_out ? io_r_23_b : _GEN_9322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9324 = 8'h18 == r_count_45_io_out ? io_r_24_b : _GEN_9323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9325 = 8'h19 == r_count_45_io_out ? io_r_25_b : _GEN_9324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9326 = 8'h1a == r_count_45_io_out ? io_r_26_b : _GEN_9325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9327 = 8'h1b == r_count_45_io_out ? io_r_27_b : _GEN_9326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9328 = 8'h1c == r_count_45_io_out ? io_r_28_b : _GEN_9327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9329 = 8'h1d == r_count_45_io_out ? io_r_29_b : _GEN_9328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9330 = 8'h1e == r_count_45_io_out ? io_r_30_b : _GEN_9329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9331 = 8'h1f == r_count_45_io_out ? io_r_31_b : _GEN_9330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9332 = 8'h20 == r_count_45_io_out ? io_r_32_b : _GEN_9331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9333 = 8'h21 == r_count_45_io_out ? io_r_33_b : _GEN_9332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9334 = 8'h22 == r_count_45_io_out ? io_r_34_b : _GEN_9333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9335 = 8'h23 == r_count_45_io_out ? io_r_35_b : _GEN_9334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9336 = 8'h24 == r_count_45_io_out ? io_r_36_b : _GEN_9335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9337 = 8'h25 == r_count_45_io_out ? io_r_37_b : _GEN_9336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9338 = 8'h26 == r_count_45_io_out ? io_r_38_b : _GEN_9337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9339 = 8'h27 == r_count_45_io_out ? io_r_39_b : _GEN_9338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9340 = 8'h28 == r_count_45_io_out ? io_r_40_b : _GEN_9339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9341 = 8'h29 == r_count_45_io_out ? io_r_41_b : _GEN_9340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9342 = 8'h2a == r_count_45_io_out ? io_r_42_b : _GEN_9341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9343 = 8'h2b == r_count_45_io_out ? io_r_43_b : _GEN_9342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9344 = 8'h2c == r_count_45_io_out ? io_r_44_b : _GEN_9343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9345 = 8'h2d == r_count_45_io_out ? io_r_45_b : _GEN_9344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9346 = 8'h2e == r_count_45_io_out ? io_r_46_b : _GEN_9345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9347 = 8'h2f == r_count_45_io_out ? io_r_47_b : _GEN_9346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9348 = 8'h30 == r_count_45_io_out ? io_r_48_b : _GEN_9347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9349 = 8'h31 == r_count_45_io_out ? io_r_49_b : _GEN_9348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9350 = 8'h32 == r_count_45_io_out ? io_r_50_b : _GEN_9349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9351 = 8'h33 == r_count_45_io_out ? io_r_51_b : _GEN_9350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9352 = 8'h34 == r_count_45_io_out ? io_r_52_b : _GEN_9351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9353 = 8'h35 == r_count_45_io_out ? io_r_53_b : _GEN_9352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9354 = 8'h36 == r_count_45_io_out ? io_r_54_b : _GEN_9353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9355 = 8'h37 == r_count_45_io_out ? io_r_55_b : _GEN_9354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9356 = 8'h38 == r_count_45_io_out ? io_r_56_b : _GEN_9355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9357 = 8'h39 == r_count_45_io_out ? io_r_57_b : _GEN_9356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9358 = 8'h3a == r_count_45_io_out ? io_r_58_b : _GEN_9357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9359 = 8'h3b == r_count_45_io_out ? io_r_59_b : _GEN_9358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9360 = 8'h3c == r_count_45_io_out ? io_r_60_b : _GEN_9359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9361 = 8'h3d == r_count_45_io_out ? io_r_61_b : _GEN_9360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9362 = 8'h3e == r_count_45_io_out ? io_r_62_b : _GEN_9361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9363 = 8'h3f == r_count_45_io_out ? io_r_63_b : _GEN_9362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9364 = 8'h40 == r_count_45_io_out ? io_r_64_b : _GEN_9363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9365 = 8'h41 == r_count_45_io_out ? io_r_65_b : _GEN_9364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9366 = 8'h42 == r_count_45_io_out ? io_r_66_b : _GEN_9365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9367 = 8'h43 == r_count_45_io_out ? io_r_67_b : _GEN_9366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9368 = 8'h44 == r_count_45_io_out ? io_r_68_b : _GEN_9367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9369 = 8'h45 == r_count_45_io_out ? io_r_69_b : _GEN_9368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9370 = 8'h46 == r_count_45_io_out ? io_r_70_b : _GEN_9369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9371 = 8'h47 == r_count_45_io_out ? io_r_71_b : _GEN_9370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9372 = 8'h48 == r_count_45_io_out ? io_r_72_b : _GEN_9371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9373 = 8'h49 == r_count_45_io_out ? io_r_73_b : _GEN_9372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9374 = 8'h4a == r_count_45_io_out ? io_r_74_b : _GEN_9373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9375 = 8'h4b == r_count_45_io_out ? io_r_75_b : _GEN_9374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9376 = 8'h4c == r_count_45_io_out ? io_r_76_b : _GEN_9375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9377 = 8'h4d == r_count_45_io_out ? io_r_77_b : _GEN_9376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9378 = 8'h4e == r_count_45_io_out ? io_r_78_b : _GEN_9377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9379 = 8'h4f == r_count_45_io_out ? io_r_79_b : _GEN_9378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9380 = 8'h50 == r_count_45_io_out ? io_r_80_b : _GEN_9379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9381 = 8'h51 == r_count_45_io_out ? io_r_81_b : _GEN_9380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9382 = 8'h52 == r_count_45_io_out ? io_r_82_b : _GEN_9381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9383 = 8'h53 == r_count_45_io_out ? io_r_83_b : _GEN_9382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9384 = 8'h54 == r_count_45_io_out ? io_r_84_b : _GEN_9383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9385 = 8'h55 == r_count_45_io_out ? io_r_85_b : _GEN_9384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9386 = 8'h56 == r_count_45_io_out ? io_r_86_b : _GEN_9385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9387 = 8'h57 == r_count_45_io_out ? io_r_87_b : _GEN_9386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9388 = 8'h58 == r_count_45_io_out ? io_r_88_b : _GEN_9387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9389 = 8'h59 == r_count_45_io_out ? io_r_89_b : _GEN_9388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9390 = 8'h5a == r_count_45_io_out ? io_r_90_b : _GEN_9389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9391 = 8'h5b == r_count_45_io_out ? io_r_91_b : _GEN_9390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9392 = 8'h5c == r_count_45_io_out ? io_r_92_b : _GEN_9391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9393 = 8'h5d == r_count_45_io_out ? io_r_93_b : _GEN_9392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9394 = 8'h5e == r_count_45_io_out ? io_r_94_b : _GEN_9393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9395 = 8'h5f == r_count_45_io_out ? io_r_95_b : _GEN_9394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9396 = 8'h60 == r_count_45_io_out ? io_r_96_b : _GEN_9395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9397 = 8'h61 == r_count_45_io_out ? io_r_97_b : _GEN_9396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9398 = 8'h62 == r_count_45_io_out ? io_r_98_b : _GEN_9397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9399 = 8'h63 == r_count_45_io_out ? io_r_99_b : _GEN_9398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9400 = 8'h64 == r_count_45_io_out ? io_r_100_b : _GEN_9399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9401 = 8'h65 == r_count_45_io_out ? io_r_101_b : _GEN_9400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9402 = 8'h66 == r_count_45_io_out ? io_r_102_b : _GEN_9401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9403 = 8'h67 == r_count_45_io_out ? io_r_103_b : _GEN_9402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9404 = 8'h68 == r_count_45_io_out ? io_r_104_b : _GEN_9403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9405 = 8'h69 == r_count_45_io_out ? io_r_105_b : _GEN_9404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9406 = 8'h6a == r_count_45_io_out ? io_r_106_b : _GEN_9405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9407 = 8'h6b == r_count_45_io_out ? io_r_107_b : _GEN_9406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9408 = 8'h6c == r_count_45_io_out ? io_r_108_b : _GEN_9407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9409 = 8'h6d == r_count_45_io_out ? io_r_109_b : _GEN_9408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9410 = 8'h6e == r_count_45_io_out ? io_r_110_b : _GEN_9409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9411 = 8'h6f == r_count_45_io_out ? io_r_111_b : _GEN_9410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9412 = 8'h70 == r_count_45_io_out ? io_r_112_b : _GEN_9411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9413 = 8'h71 == r_count_45_io_out ? io_r_113_b : _GEN_9412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9414 = 8'h72 == r_count_45_io_out ? io_r_114_b : _GEN_9413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9415 = 8'h73 == r_count_45_io_out ? io_r_115_b : _GEN_9414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9416 = 8'h74 == r_count_45_io_out ? io_r_116_b : _GEN_9415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9417 = 8'h75 == r_count_45_io_out ? io_r_117_b : _GEN_9416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9418 = 8'h76 == r_count_45_io_out ? io_r_118_b : _GEN_9417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9419 = 8'h77 == r_count_45_io_out ? io_r_119_b : _GEN_9418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9420 = 8'h78 == r_count_45_io_out ? io_r_120_b : _GEN_9419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9421 = 8'h79 == r_count_45_io_out ? io_r_121_b : _GEN_9420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9422 = 8'h7a == r_count_45_io_out ? io_r_122_b : _GEN_9421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9423 = 8'h7b == r_count_45_io_out ? io_r_123_b : _GEN_9422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9424 = 8'h7c == r_count_45_io_out ? io_r_124_b : _GEN_9423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9425 = 8'h7d == r_count_45_io_out ? io_r_125_b : _GEN_9424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9426 = 8'h7e == r_count_45_io_out ? io_r_126_b : _GEN_9425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9427 = 8'h7f == r_count_45_io_out ? io_r_127_b : _GEN_9426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9428 = 8'h80 == r_count_45_io_out ? io_r_128_b : _GEN_9427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9429 = 8'h81 == r_count_45_io_out ? io_r_129_b : _GEN_9428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9430 = 8'h82 == r_count_45_io_out ? io_r_130_b : _GEN_9429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9431 = 8'h83 == r_count_45_io_out ? io_r_131_b : _GEN_9430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9432 = 8'h84 == r_count_45_io_out ? io_r_132_b : _GEN_9431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9433 = 8'h85 == r_count_45_io_out ? io_r_133_b : _GEN_9432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9434 = 8'h86 == r_count_45_io_out ? io_r_134_b : _GEN_9433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9435 = 8'h87 == r_count_45_io_out ? io_r_135_b : _GEN_9434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9436 = 8'h88 == r_count_45_io_out ? io_r_136_b : _GEN_9435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9437 = 8'h89 == r_count_45_io_out ? io_r_137_b : _GEN_9436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9438 = 8'h8a == r_count_45_io_out ? io_r_138_b : _GEN_9437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9439 = 8'h8b == r_count_45_io_out ? io_r_139_b : _GEN_9438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9440 = 8'h8c == r_count_45_io_out ? io_r_140_b : _GEN_9439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9441 = 8'h8d == r_count_45_io_out ? io_r_141_b : _GEN_9440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9442 = 8'h8e == r_count_45_io_out ? io_r_142_b : _GEN_9441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9443 = 8'h8f == r_count_45_io_out ? io_r_143_b : _GEN_9442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9444 = 8'h90 == r_count_45_io_out ? io_r_144_b : _GEN_9443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9445 = 8'h91 == r_count_45_io_out ? io_r_145_b : _GEN_9444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9446 = 8'h92 == r_count_45_io_out ? io_r_146_b : _GEN_9445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9447 = 8'h93 == r_count_45_io_out ? io_r_147_b : _GEN_9446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9448 = 8'h94 == r_count_45_io_out ? io_r_148_b : _GEN_9447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9449 = 8'h95 == r_count_45_io_out ? io_r_149_b : _GEN_9448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9450 = 8'h96 == r_count_45_io_out ? io_r_150_b : _GEN_9449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9451 = 8'h97 == r_count_45_io_out ? io_r_151_b : _GEN_9450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9452 = 8'h98 == r_count_45_io_out ? io_r_152_b : _GEN_9451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9453 = 8'h99 == r_count_45_io_out ? io_r_153_b : _GEN_9452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9454 = 8'h9a == r_count_45_io_out ? io_r_154_b : _GEN_9453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9455 = 8'h9b == r_count_45_io_out ? io_r_155_b : _GEN_9454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9456 = 8'h9c == r_count_45_io_out ? io_r_156_b : _GEN_9455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9457 = 8'h9d == r_count_45_io_out ? io_r_157_b : _GEN_9456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9458 = 8'h9e == r_count_45_io_out ? io_r_158_b : _GEN_9457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9459 = 8'h9f == r_count_45_io_out ? io_r_159_b : _GEN_9458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9460 = 8'ha0 == r_count_45_io_out ? io_r_160_b : _GEN_9459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9461 = 8'ha1 == r_count_45_io_out ? io_r_161_b : _GEN_9460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9462 = 8'ha2 == r_count_45_io_out ? io_r_162_b : _GEN_9461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9463 = 8'ha3 == r_count_45_io_out ? io_r_163_b : _GEN_9462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9464 = 8'ha4 == r_count_45_io_out ? io_r_164_b : _GEN_9463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9465 = 8'ha5 == r_count_45_io_out ? io_r_165_b : _GEN_9464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9466 = 8'ha6 == r_count_45_io_out ? io_r_166_b : _GEN_9465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9467 = 8'ha7 == r_count_45_io_out ? io_r_167_b : _GEN_9466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9468 = 8'ha8 == r_count_45_io_out ? io_r_168_b : _GEN_9467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9469 = 8'ha9 == r_count_45_io_out ? io_r_169_b : _GEN_9468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9470 = 8'haa == r_count_45_io_out ? io_r_170_b : _GEN_9469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9471 = 8'hab == r_count_45_io_out ? io_r_171_b : _GEN_9470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9472 = 8'hac == r_count_45_io_out ? io_r_172_b : _GEN_9471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9473 = 8'had == r_count_45_io_out ? io_r_173_b : _GEN_9472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9474 = 8'hae == r_count_45_io_out ? io_r_174_b : _GEN_9473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9475 = 8'haf == r_count_45_io_out ? io_r_175_b : _GEN_9474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9476 = 8'hb0 == r_count_45_io_out ? io_r_176_b : _GEN_9475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9477 = 8'hb1 == r_count_45_io_out ? io_r_177_b : _GEN_9476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9478 = 8'hb2 == r_count_45_io_out ? io_r_178_b : _GEN_9477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9479 = 8'hb3 == r_count_45_io_out ? io_r_179_b : _GEN_9478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9480 = 8'hb4 == r_count_45_io_out ? io_r_180_b : _GEN_9479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9481 = 8'hb5 == r_count_45_io_out ? io_r_181_b : _GEN_9480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9482 = 8'hb6 == r_count_45_io_out ? io_r_182_b : _GEN_9481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9483 = 8'hb7 == r_count_45_io_out ? io_r_183_b : _GEN_9482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9484 = 8'hb8 == r_count_45_io_out ? io_r_184_b : _GEN_9483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9485 = 8'hb9 == r_count_45_io_out ? io_r_185_b : _GEN_9484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9486 = 8'hba == r_count_45_io_out ? io_r_186_b : _GEN_9485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9487 = 8'hbb == r_count_45_io_out ? io_r_187_b : _GEN_9486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9488 = 8'hbc == r_count_45_io_out ? io_r_188_b : _GEN_9487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9489 = 8'hbd == r_count_45_io_out ? io_r_189_b : _GEN_9488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9490 = 8'hbe == r_count_45_io_out ? io_r_190_b : _GEN_9489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9491 = 8'hbf == r_count_45_io_out ? io_r_191_b : _GEN_9490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9492 = 8'hc0 == r_count_45_io_out ? io_r_192_b : _GEN_9491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9493 = 8'hc1 == r_count_45_io_out ? io_r_193_b : _GEN_9492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9494 = 8'hc2 == r_count_45_io_out ? io_r_194_b : _GEN_9493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9495 = 8'hc3 == r_count_45_io_out ? io_r_195_b : _GEN_9494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9496 = 8'hc4 == r_count_45_io_out ? io_r_196_b : _GEN_9495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9497 = 8'hc5 == r_count_45_io_out ? io_r_197_b : _GEN_9496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9498 = 8'hc6 == r_count_45_io_out ? io_r_198_b : _GEN_9497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9501 = 8'h1 == r_count_46_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9502 = 8'h2 == r_count_46_io_out ? io_r_2_b : _GEN_9501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9503 = 8'h3 == r_count_46_io_out ? io_r_3_b : _GEN_9502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9504 = 8'h4 == r_count_46_io_out ? io_r_4_b : _GEN_9503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9505 = 8'h5 == r_count_46_io_out ? io_r_5_b : _GEN_9504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9506 = 8'h6 == r_count_46_io_out ? io_r_6_b : _GEN_9505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9507 = 8'h7 == r_count_46_io_out ? io_r_7_b : _GEN_9506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9508 = 8'h8 == r_count_46_io_out ? io_r_8_b : _GEN_9507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9509 = 8'h9 == r_count_46_io_out ? io_r_9_b : _GEN_9508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9510 = 8'ha == r_count_46_io_out ? io_r_10_b : _GEN_9509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9511 = 8'hb == r_count_46_io_out ? io_r_11_b : _GEN_9510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9512 = 8'hc == r_count_46_io_out ? io_r_12_b : _GEN_9511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9513 = 8'hd == r_count_46_io_out ? io_r_13_b : _GEN_9512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9514 = 8'he == r_count_46_io_out ? io_r_14_b : _GEN_9513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9515 = 8'hf == r_count_46_io_out ? io_r_15_b : _GEN_9514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9516 = 8'h10 == r_count_46_io_out ? io_r_16_b : _GEN_9515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9517 = 8'h11 == r_count_46_io_out ? io_r_17_b : _GEN_9516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9518 = 8'h12 == r_count_46_io_out ? io_r_18_b : _GEN_9517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9519 = 8'h13 == r_count_46_io_out ? io_r_19_b : _GEN_9518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9520 = 8'h14 == r_count_46_io_out ? io_r_20_b : _GEN_9519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9521 = 8'h15 == r_count_46_io_out ? io_r_21_b : _GEN_9520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9522 = 8'h16 == r_count_46_io_out ? io_r_22_b : _GEN_9521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9523 = 8'h17 == r_count_46_io_out ? io_r_23_b : _GEN_9522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9524 = 8'h18 == r_count_46_io_out ? io_r_24_b : _GEN_9523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9525 = 8'h19 == r_count_46_io_out ? io_r_25_b : _GEN_9524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9526 = 8'h1a == r_count_46_io_out ? io_r_26_b : _GEN_9525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9527 = 8'h1b == r_count_46_io_out ? io_r_27_b : _GEN_9526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9528 = 8'h1c == r_count_46_io_out ? io_r_28_b : _GEN_9527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9529 = 8'h1d == r_count_46_io_out ? io_r_29_b : _GEN_9528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9530 = 8'h1e == r_count_46_io_out ? io_r_30_b : _GEN_9529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9531 = 8'h1f == r_count_46_io_out ? io_r_31_b : _GEN_9530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9532 = 8'h20 == r_count_46_io_out ? io_r_32_b : _GEN_9531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9533 = 8'h21 == r_count_46_io_out ? io_r_33_b : _GEN_9532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9534 = 8'h22 == r_count_46_io_out ? io_r_34_b : _GEN_9533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9535 = 8'h23 == r_count_46_io_out ? io_r_35_b : _GEN_9534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9536 = 8'h24 == r_count_46_io_out ? io_r_36_b : _GEN_9535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9537 = 8'h25 == r_count_46_io_out ? io_r_37_b : _GEN_9536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9538 = 8'h26 == r_count_46_io_out ? io_r_38_b : _GEN_9537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9539 = 8'h27 == r_count_46_io_out ? io_r_39_b : _GEN_9538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9540 = 8'h28 == r_count_46_io_out ? io_r_40_b : _GEN_9539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9541 = 8'h29 == r_count_46_io_out ? io_r_41_b : _GEN_9540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9542 = 8'h2a == r_count_46_io_out ? io_r_42_b : _GEN_9541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9543 = 8'h2b == r_count_46_io_out ? io_r_43_b : _GEN_9542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9544 = 8'h2c == r_count_46_io_out ? io_r_44_b : _GEN_9543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9545 = 8'h2d == r_count_46_io_out ? io_r_45_b : _GEN_9544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9546 = 8'h2e == r_count_46_io_out ? io_r_46_b : _GEN_9545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9547 = 8'h2f == r_count_46_io_out ? io_r_47_b : _GEN_9546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9548 = 8'h30 == r_count_46_io_out ? io_r_48_b : _GEN_9547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9549 = 8'h31 == r_count_46_io_out ? io_r_49_b : _GEN_9548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9550 = 8'h32 == r_count_46_io_out ? io_r_50_b : _GEN_9549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9551 = 8'h33 == r_count_46_io_out ? io_r_51_b : _GEN_9550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9552 = 8'h34 == r_count_46_io_out ? io_r_52_b : _GEN_9551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9553 = 8'h35 == r_count_46_io_out ? io_r_53_b : _GEN_9552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9554 = 8'h36 == r_count_46_io_out ? io_r_54_b : _GEN_9553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9555 = 8'h37 == r_count_46_io_out ? io_r_55_b : _GEN_9554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9556 = 8'h38 == r_count_46_io_out ? io_r_56_b : _GEN_9555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9557 = 8'h39 == r_count_46_io_out ? io_r_57_b : _GEN_9556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9558 = 8'h3a == r_count_46_io_out ? io_r_58_b : _GEN_9557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9559 = 8'h3b == r_count_46_io_out ? io_r_59_b : _GEN_9558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9560 = 8'h3c == r_count_46_io_out ? io_r_60_b : _GEN_9559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9561 = 8'h3d == r_count_46_io_out ? io_r_61_b : _GEN_9560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9562 = 8'h3e == r_count_46_io_out ? io_r_62_b : _GEN_9561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9563 = 8'h3f == r_count_46_io_out ? io_r_63_b : _GEN_9562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9564 = 8'h40 == r_count_46_io_out ? io_r_64_b : _GEN_9563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9565 = 8'h41 == r_count_46_io_out ? io_r_65_b : _GEN_9564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9566 = 8'h42 == r_count_46_io_out ? io_r_66_b : _GEN_9565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9567 = 8'h43 == r_count_46_io_out ? io_r_67_b : _GEN_9566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9568 = 8'h44 == r_count_46_io_out ? io_r_68_b : _GEN_9567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9569 = 8'h45 == r_count_46_io_out ? io_r_69_b : _GEN_9568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9570 = 8'h46 == r_count_46_io_out ? io_r_70_b : _GEN_9569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9571 = 8'h47 == r_count_46_io_out ? io_r_71_b : _GEN_9570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9572 = 8'h48 == r_count_46_io_out ? io_r_72_b : _GEN_9571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9573 = 8'h49 == r_count_46_io_out ? io_r_73_b : _GEN_9572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9574 = 8'h4a == r_count_46_io_out ? io_r_74_b : _GEN_9573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9575 = 8'h4b == r_count_46_io_out ? io_r_75_b : _GEN_9574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9576 = 8'h4c == r_count_46_io_out ? io_r_76_b : _GEN_9575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9577 = 8'h4d == r_count_46_io_out ? io_r_77_b : _GEN_9576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9578 = 8'h4e == r_count_46_io_out ? io_r_78_b : _GEN_9577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9579 = 8'h4f == r_count_46_io_out ? io_r_79_b : _GEN_9578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9580 = 8'h50 == r_count_46_io_out ? io_r_80_b : _GEN_9579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9581 = 8'h51 == r_count_46_io_out ? io_r_81_b : _GEN_9580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9582 = 8'h52 == r_count_46_io_out ? io_r_82_b : _GEN_9581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9583 = 8'h53 == r_count_46_io_out ? io_r_83_b : _GEN_9582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9584 = 8'h54 == r_count_46_io_out ? io_r_84_b : _GEN_9583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9585 = 8'h55 == r_count_46_io_out ? io_r_85_b : _GEN_9584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9586 = 8'h56 == r_count_46_io_out ? io_r_86_b : _GEN_9585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9587 = 8'h57 == r_count_46_io_out ? io_r_87_b : _GEN_9586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9588 = 8'h58 == r_count_46_io_out ? io_r_88_b : _GEN_9587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9589 = 8'h59 == r_count_46_io_out ? io_r_89_b : _GEN_9588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9590 = 8'h5a == r_count_46_io_out ? io_r_90_b : _GEN_9589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9591 = 8'h5b == r_count_46_io_out ? io_r_91_b : _GEN_9590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9592 = 8'h5c == r_count_46_io_out ? io_r_92_b : _GEN_9591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9593 = 8'h5d == r_count_46_io_out ? io_r_93_b : _GEN_9592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9594 = 8'h5e == r_count_46_io_out ? io_r_94_b : _GEN_9593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9595 = 8'h5f == r_count_46_io_out ? io_r_95_b : _GEN_9594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9596 = 8'h60 == r_count_46_io_out ? io_r_96_b : _GEN_9595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9597 = 8'h61 == r_count_46_io_out ? io_r_97_b : _GEN_9596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9598 = 8'h62 == r_count_46_io_out ? io_r_98_b : _GEN_9597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9599 = 8'h63 == r_count_46_io_out ? io_r_99_b : _GEN_9598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9600 = 8'h64 == r_count_46_io_out ? io_r_100_b : _GEN_9599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9601 = 8'h65 == r_count_46_io_out ? io_r_101_b : _GEN_9600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9602 = 8'h66 == r_count_46_io_out ? io_r_102_b : _GEN_9601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9603 = 8'h67 == r_count_46_io_out ? io_r_103_b : _GEN_9602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9604 = 8'h68 == r_count_46_io_out ? io_r_104_b : _GEN_9603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9605 = 8'h69 == r_count_46_io_out ? io_r_105_b : _GEN_9604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9606 = 8'h6a == r_count_46_io_out ? io_r_106_b : _GEN_9605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9607 = 8'h6b == r_count_46_io_out ? io_r_107_b : _GEN_9606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9608 = 8'h6c == r_count_46_io_out ? io_r_108_b : _GEN_9607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9609 = 8'h6d == r_count_46_io_out ? io_r_109_b : _GEN_9608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9610 = 8'h6e == r_count_46_io_out ? io_r_110_b : _GEN_9609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9611 = 8'h6f == r_count_46_io_out ? io_r_111_b : _GEN_9610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9612 = 8'h70 == r_count_46_io_out ? io_r_112_b : _GEN_9611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9613 = 8'h71 == r_count_46_io_out ? io_r_113_b : _GEN_9612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9614 = 8'h72 == r_count_46_io_out ? io_r_114_b : _GEN_9613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9615 = 8'h73 == r_count_46_io_out ? io_r_115_b : _GEN_9614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9616 = 8'h74 == r_count_46_io_out ? io_r_116_b : _GEN_9615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9617 = 8'h75 == r_count_46_io_out ? io_r_117_b : _GEN_9616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9618 = 8'h76 == r_count_46_io_out ? io_r_118_b : _GEN_9617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9619 = 8'h77 == r_count_46_io_out ? io_r_119_b : _GEN_9618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9620 = 8'h78 == r_count_46_io_out ? io_r_120_b : _GEN_9619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9621 = 8'h79 == r_count_46_io_out ? io_r_121_b : _GEN_9620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9622 = 8'h7a == r_count_46_io_out ? io_r_122_b : _GEN_9621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9623 = 8'h7b == r_count_46_io_out ? io_r_123_b : _GEN_9622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9624 = 8'h7c == r_count_46_io_out ? io_r_124_b : _GEN_9623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9625 = 8'h7d == r_count_46_io_out ? io_r_125_b : _GEN_9624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9626 = 8'h7e == r_count_46_io_out ? io_r_126_b : _GEN_9625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9627 = 8'h7f == r_count_46_io_out ? io_r_127_b : _GEN_9626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9628 = 8'h80 == r_count_46_io_out ? io_r_128_b : _GEN_9627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9629 = 8'h81 == r_count_46_io_out ? io_r_129_b : _GEN_9628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9630 = 8'h82 == r_count_46_io_out ? io_r_130_b : _GEN_9629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9631 = 8'h83 == r_count_46_io_out ? io_r_131_b : _GEN_9630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9632 = 8'h84 == r_count_46_io_out ? io_r_132_b : _GEN_9631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9633 = 8'h85 == r_count_46_io_out ? io_r_133_b : _GEN_9632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9634 = 8'h86 == r_count_46_io_out ? io_r_134_b : _GEN_9633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9635 = 8'h87 == r_count_46_io_out ? io_r_135_b : _GEN_9634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9636 = 8'h88 == r_count_46_io_out ? io_r_136_b : _GEN_9635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9637 = 8'h89 == r_count_46_io_out ? io_r_137_b : _GEN_9636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9638 = 8'h8a == r_count_46_io_out ? io_r_138_b : _GEN_9637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9639 = 8'h8b == r_count_46_io_out ? io_r_139_b : _GEN_9638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9640 = 8'h8c == r_count_46_io_out ? io_r_140_b : _GEN_9639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9641 = 8'h8d == r_count_46_io_out ? io_r_141_b : _GEN_9640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9642 = 8'h8e == r_count_46_io_out ? io_r_142_b : _GEN_9641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9643 = 8'h8f == r_count_46_io_out ? io_r_143_b : _GEN_9642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9644 = 8'h90 == r_count_46_io_out ? io_r_144_b : _GEN_9643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9645 = 8'h91 == r_count_46_io_out ? io_r_145_b : _GEN_9644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9646 = 8'h92 == r_count_46_io_out ? io_r_146_b : _GEN_9645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9647 = 8'h93 == r_count_46_io_out ? io_r_147_b : _GEN_9646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9648 = 8'h94 == r_count_46_io_out ? io_r_148_b : _GEN_9647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9649 = 8'h95 == r_count_46_io_out ? io_r_149_b : _GEN_9648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9650 = 8'h96 == r_count_46_io_out ? io_r_150_b : _GEN_9649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9651 = 8'h97 == r_count_46_io_out ? io_r_151_b : _GEN_9650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9652 = 8'h98 == r_count_46_io_out ? io_r_152_b : _GEN_9651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9653 = 8'h99 == r_count_46_io_out ? io_r_153_b : _GEN_9652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9654 = 8'h9a == r_count_46_io_out ? io_r_154_b : _GEN_9653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9655 = 8'h9b == r_count_46_io_out ? io_r_155_b : _GEN_9654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9656 = 8'h9c == r_count_46_io_out ? io_r_156_b : _GEN_9655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9657 = 8'h9d == r_count_46_io_out ? io_r_157_b : _GEN_9656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9658 = 8'h9e == r_count_46_io_out ? io_r_158_b : _GEN_9657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9659 = 8'h9f == r_count_46_io_out ? io_r_159_b : _GEN_9658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9660 = 8'ha0 == r_count_46_io_out ? io_r_160_b : _GEN_9659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9661 = 8'ha1 == r_count_46_io_out ? io_r_161_b : _GEN_9660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9662 = 8'ha2 == r_count_46_io_out ? io_r_162_b : _GEN_9661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9663 = 8'ha3 == r_count_46_io_out ? io_r_163_b : _GEN_9662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9664 = 8'ha4 == r_count_46_io_out ? io_r_164_b : _GEN_9663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9665 = 8'ha5 == r_count_46_io_out ? io_r_165_b : _GEN_9664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9666 = 8'ha6 == r_count_46_io_out ? io_r_166_b : _GEN_9665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9667 = 8'ha7 == r_count_46_io_out ? io_r_167_b : _GEN_9666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9668 = 8'ha8 == r_count_46_io_out ? io_r_168_b : _GEN_9667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9669 = 8'ha9 == r_count_46_io_out ? io_r_169_b : _GEN_9668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9670 = 8'haa == r_count_46_io_out ? io_r_170_b : _GEN_9669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9671 = 8'hab == r_count_46_io_out ? io_r_171_b : _GEN_9670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9672 = 8'hac == r_count_46_io_out ? io_r_172_b : _GEN_9671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9673 = 8'had == r_count_46_io_out ? io_r_173_b : _GEN_9672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9674 = 8'hae == r_count_46_io_out ? io_r_174_b : _GEN_9673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9675 = 8'haf == r_count_46_io_out ? io_r_175_b : _GEN_9674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9676 = 8'hb0 == r_count_46_io_out ? io_r_176_b : _GEN_9675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9677 = 8'hb1 == r_count_46_io_out ? io_r_177_b : _GEN_9676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9678 = 8'hb2 == r_count_46_io_out ? io_r_178_b : _GEN_9677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9679 = 8'hb3 == r_count_46_io_out ? io_r_179_b : _GEN_9678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9680 = 8'hb4 == r_count_46_io_out ? io_r_180_b : _GEN_9679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9681 = 8'hb5 == r_count_46_io_out ? io_r_181_b : _GEN_9680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9682 = 8'hb6 == r_count_46_io_out ? io_r_182_b : _GEN_9681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9683 = 8'hb7 == r_count_46_io_out ? io_r_183_b : _GEN_9682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9684 = 8'hb8 == r_count_46_io_out ? io_r_184_b : _GEN_9683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9685 = 8'hb9 == r_count_46_io_out ? io_r_185_b : _GEN_9684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9686 = 8'hba == r_count_46_io_out ? io_r_186_b : _GEN_9685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9687 = 8'hbb == r_count_46_io_out ? io_r_187_b : _GEN_9686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9688 = 8'hbc == r_count_46_io_out ? io_r_188_b : _GEN_9687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9689 = 8'hbd == r_count_46_io_out ? io_r_189_b : _GEN_9688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9690 = 8'hbe == r_count_46_io_out ? io_r_190_b : _GEN_9689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9691 = 8'hbf == r_count_46_io_out ? io_r_191_b : _GEN_9690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9692 = 8'hc0 == r_count_46_io_out ? io_r_192_b : _GEN_9691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9693 = 8'hc1 == r_count_46_io_out ? io_r_193_b : _GEN_9692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9694 = 8'hc2 == r_count_46_io_out ? io_r_194_b : _GEN_9693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9695 = 8'hc3 == r_count_46_io_out ? io_r_195_b : _GEN_9694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9696 = 8'hc4 == r_count_46_io_out ? io_r_196_b : _GEN_9695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9697 = 8'hc5 == r_count_46_io_out ? io_r_197_b : _GEN_9696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9698 = 8'hc6 == r_count_46_io_out ? io_r_198_b : _GEN_9697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9701 = 8'h1 == r_count_47_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9702 = 8'h2 == r_count_47_io_out ? io_r_2_b : _GEN_9701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9703 = 8'h3 == r_count_47_io_out ? io_r_3_b : _GEN_9702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9704 = 8'h4 == r_count_47_io_out ? io_r_4_b : _GEN_9703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9705 = 8'h5 == r_count_47_io_out ? io_r_5_b : _GEN_9704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9706 = 8'h6 == r_count_47_io_out ? io_r_6_b : _GEN_9705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9707 = 8'h7 == r_count_47_io_out ? io_r_7_b : _GEN_9706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9708 = 8'h8 == r_count_47_io_out ? io_r_8_b : _GEN_9707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9709 = 8'h9 == r_count_47_io_out ? io_r_9_b : _GEN_9708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9710 = 8'ha == r_count_47_io_out ? io_r_10_b : _GEN_9709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9711 = 8'hb == r_count_47_io_out ? io_r_11_b : _GEN_9710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9712 = 8'hc == r_count_47_io_out ? io_r_12_b : _GEN_9711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9713 = 8'hd == r_count_47_io_out ? io_r_13_b : _GEN_9712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9714 = 8'he == r_count_47_io_out ? io_r_14_b : _GEN_9713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9715 = 8'hf == r_count_47_io_out ? io_r_15_b : _GEN_9714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9716 = 8'h10 == r_count_47_io_out ? io_r_16_b : _GEN_9715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9717 = 8'h11 == r_count_47_io_out ? io_r_17_b : _GEN_9716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9718 = 8'h12 == r_count_47_io_out ? io_r_18_b : _GEN_9717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9719 = 8'h13 == r_count_47_io_out ? io_r_19_b : _GEN_9718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9720 = 8'h14 == r_count_47_io_out ? io_r_20_b : _GEN_9719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9721 = 8'h15 == r_count_47_io_out ? io_r_21_b : _GEN_9720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9722 = 8'h16 == r_count_47_io_out ? io_r_22_b : _GEN_9721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9723 = 8'h17 == r_count_47_io_out ? io_r_23_b : _GEN_9722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9724 = 8'h18 == r_count_47_io_out ? io_r_24_b : _GEN_9723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9725 = 8'h19 == r_count_47_io_out ? io_r_25_b : _GEN_9724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9726 = 8'h1a == r_count_47_io_out ? io_r_26_b : _GEN_9725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9727 = 8'h1b == r_count_47_io_out ? io_r_27_b : _GEN_9726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9728 = 8'h1c == r_count_47_io_out ? io_r_28_b : _GEN_9727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9729 = 8'h1d == r_count_47_io_out ? io_r_29_b : _GEN_9728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9730 = 8'h1e == r_count_47_io_out ? io_r_30_b : _GEN_9729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9731 = 8'h1f == r_count_47_io_out ? io_r_31_b : _GEN_9730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9732 = 8'h20 == r_count_47_io_out ? io_r_32_b : _GEN_9731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9733 = 8'h21 == r_count_47_io_out ? io_r_33_b : _GEN_9732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9734 = 8'h22 == r_count_47_io_out ? io_r_34_b : _GEN_9733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9735 = 8'h23 == r_count_47_io_out ? io_r_35_b : _GEN_9734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9736 = 8'h24 == r_count_47_io_out ? io_r_36_b : _GEN_9735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9737 = 8'h25 == r_count_47_io_out ? io_r_37_b : _GEN_9736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9738 = 8'h26 == r_count_47_io_out ? io_r_38_b : _GEN_9737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9739 = 8'h27 == r_count_47_io_out ? io_r_39_b : _GEN_9738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9740 = 8'h28 == r_count_47_io_out ? io_r_40_b : _GEN_9739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9741 = 8'h29 == r_count_47_io_out ? io_r_41_b : _GEN_9740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9742 = 8'h2a == r_count_47_io_out ? io_r_42_b : _GEN_9741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9743 = 8'h2b == r_count_47_io_out ? io_r_43_b : _GEN_9742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9744 = 8'h2c == r_count_47_io_out ? io_r_44_b : _GEN_9743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9745 = 8'h2d == r_count_47_io_out ? io_r_45_b : _GEN_9744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9746 = 8'h2e == r_count_47_io_out ? io_r_46_b : _GEN_9745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9747 = 8'h2f == r_count_47_io_out ? io_r_47_b : _GEN_9746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9748 = 8'h30 == r_count_47_io_out ? io_r_48_b : _GEN_9747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9749 = 8'h31 == r_count_47_io_out ? io_r_49_b : _GEN_9748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9750 = 8'h32 == r_count_47_io_out ? io_r_50_b : _GEN_9749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9751 = 8'h33 == r_count_47_io_out ? io_r_51_b : _GEN_9750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9752 = 8'h34 == r_count_47_io_out ? io_r_52_b : _GEN_9751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9753 = 8'h35 == r_count_47_io_out ? io_r_53_b : _GEN_9752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9754 = 8'h36 == r_count_47_io_out ? io_r_54_b : _GEN_9753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9755 = 8'h37 == r_count_47_io_out ? io_r_55_b : _GEN_9754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9756 = 8'h38 == r_count_47_io_out ? io_r_56_b : _GEN_9755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9757 = 8'h39 == r_count_47_io_out ? io_r_57_b : _GEN_9756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9758 = 8'h3a == r_count_47_io_out ? io_r_58_b : _GEN_9757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9759 = 8'h3b == r_count_47_io_out ? io_r_59_b : _GEN_9758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9760 = 8'h3c == r_count_47_io_out ? io_r_60_b : _GEN_9759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9761 = 8'h3d == r_count_47_io_out ? io_r_61_b : _GEN_9760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9762 = 8'h3e == r_count_47_io_out ? io_r_62_b : _GEN_9761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9763 = 8'h3f == r_count_47_io_out ? io_r_63_b : _GEN_9762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9764 = 8'h40 == r_count_47_io_out ? io_r_64_b : _GEN_9763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9765 = 8'h41 == r_count_47_io_out ? io_r_65_b : _GEN_9764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9766 = 8'h42 == r_count_47_io_out ? io_r_66_b : _GEN_9765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9767 = 8'h43 == r_count_47_io_out ? io_r_67_b : _GEN_9766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9768 = 8'h44 == r_count_47_io_out ? io_r_68_b : _GEN_9767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9769 = 8'h45 == r_count_47_io_out ? io_r_69_b : _GEN_9768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9770 = 8'h46 == r_count_47_io_out ? io_r_70_b : _GEN_9769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9771 = 8'h47 == r_count_47_io_out ? io_r_71_b : _GEN_9770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9772 = 8'h48 == r_count_47_io_out ? io_r_72_b : _GEN_9771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9773 = 8'h49 == r_count_47_io_out ? io_r_73_b : _GEN_9772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9774 = 8'h4a == r_count_47_io_out ? io_r_74_b : _GEN_9773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9775 = 8'h4b == r_count_47_io_out ? io_r_75_b : _GEN_9774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9776 = 8'h4c == r_count_47_io_out ? io_r_76_b : _GEN_9775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9777 = 8'h4d == r_count_47_io_out ? io_r_77_b : _GEN_9776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9778 = 8'h4e == r_count_47_io_out ? io_r_78_b : _GEN_9777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9779 = 8'h4f == r_count_47_io_out ? io_r_79_b : _GEN_9778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9780 = 8'h50 == r_count_47_io_out ? io_r_80_b : _GEN_9779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9781 = 8'h51 == r_count_47_io_out ? io_r_81_b : _GEN_9780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9782 = 8'h52 == r_count_47_io_out ? io_r_82_b : _GEN_9781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9783 = 8'h53 == r_count_47_io_out ? io_r_83_b : _GEN_9782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9784 = 8'h54 == r_count_47_io_out ? io_r_84_b : _GEN_9783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9785 = 8'h55 == r_count_47_io_out ? io_r_85_b : _GEN_9784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9786 = 8'h56 == r_count_47_io_out ? io_r_86_b : _GEN_9785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9787 = 8'h57 == r_count_47_io_out ? io_r_87_b : _GEN_9786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9788 = 8'h58 == r_count_47_io_out ? io_r_88_b : _GEN_9787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9789 = 8'h59 == r_count_47_io_out ? io_r_89_b : _GEN_9788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9790 = 8'h5a == r_count_47_io_out ? io_r_90_b : _GEN_9789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9791 = 8'h5b == r_count_47_io_out ? io_r_91_b : _GEN_9790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9792 = 8'h5c == r_count_47_io_out ? io_r_92_b : _GEN_9791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9793 = 8'h5d == r_count_47_io_out ? io_r_93_b : _GEN_9792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9794 = 8'h5e == r_count_47_io_out ? io_r_94_b : _GEN_9793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9795 = 8'h5f == r_count_47_io_out ? io_r_95_b : _GEN_9794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9796 = 8'h60 == r_count_47_io_out ? io_r_96_b : _GEN_9795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9797 = 8'h61 == r_count_47_io_out ? io_r_97_b : _GEN_9796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9798 = 8'h62 == r_count_47_io_out ? io_r_98_b : _GEN_9797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9799 = 8'h63 == r_count_47_io_out ? io_r_99_b : _GEN_9798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9800 = 8'h64 == r_count_47_io_out ? io_r_100_b : _GEN_9799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9801 = 8'h65 == r_count_47_io_out ? io_r_101_b : _GEN_9800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9802 = 8'h66 == r_count_47_io_out ? io_r_102_b : _GEN_9801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9803 = 8'h67 == r_count_47_io_out ? io_r_103_b : _GEN_9802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9804 = 8'h68 == r_count_47_io_out ? io_r_104_b : _GEN_9803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9805 = 8'h69 == r_count_47_io_out ? io_r_105_b : _GEN_9804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9806 = 8'h6a == r_count_47_io_out ? io_r_106_b : _GEN_9805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9807 = 8'h6b == r_count_47_io_out ? io_r_107_b : _GEN_9806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9808 = 8'h6c == r_count_47_io_out ? io_r_108_b : _GEN_9807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9809 = 8'h6d == r_count_47_io_out ? io_r_109_b : _GEN_9808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9810 = 8'h6e == r_count_47_io_out ? io_r_110_b : _GEN_9809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9811 = 8'h6f == r_count_47_io_out ? io_r_111_b : _GEN_9810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9812 = 8'h70 == r_count_47_io_out ? io_r_112_b : _GEN_9811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9813 = 8'h71 == r_count_47_io_out ? io_r_113_b : _GEN_9812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9814 = 8'h72 == r_count_47_io_out ? io_r_114_b : _GEN_9813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9815 = 8'h73 == r_count_47_io_out ? io_r_115_b : _GEN_9814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9816 = 8'h74 == r_count_47_io_out ? io_r_116_b : _GEN_9815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9817 = 8'h75 == r_count_47_io_out ? io_r_117_b : _GEN_9816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9818 = 8'h76 == r_count_47_io_out ? io_r_118_b : _GEN_9817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9819 = 8'h77 == r_count_47_io_out ? io_r_119_b : _GEN_9818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9820 = 8'h78 == r_count_47_io_out ? io_r_120_b : _GEN_9819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9821 = 8'h79 == r_count_47_io_out ? io_r_121_b : _GEN_9820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9822 = 8'h7a == r_count_47_io_out ? io_r_122_b : _GEN_9821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9823 = 8'h7b == r_count_47_io_out ? io_r_123_b : _GEN_9822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9824 = 8'h7c == r_count_47_io_out ? io_r_124_b : _GEN_9823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9825 = 8'h7d == r_count_47_io_out ? io_r_125_b : _GEN_9824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9826 = 8'h7e == r_count_47_io_out ? io_r_126_b : _GEN_9825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9827 = 8'h7f == r_count_47_io_out ? io_r_127_b : _GEN_9826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9828 = 8'h80 == r_count_47_io_out ? io_r_128_b : _GEN_9827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9829 = 8'h81 == r_count_47_io_out ? io_r_129_b : _GEN_9828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9830 = 8'h82 == r_count_47_io_out ? io_r_130_b : _GEN_9829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9831 = 8'h83 == r_count_47_io_out ? io_r_131_b : _GEN_9830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9832 = 8'h84 == r_count_47_io_out ? io_r_132_b : _GEN_9831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9833 = 8'h85 == r_count_47_io_out ? io_r_133_b : _GEN_9832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9834 = 8'h86 == r_count_47_io_out ? io_r_134_b : _GEN_9833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9835 = 8'h87 == r_count_47_io_out ? io_r_135_b : _GEN_9834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9836 = 8'h88 == r_count_47_io_out ? io_r_136_b : _GEN_9835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9837 = 8'h89 == r_count_47_io_out ? io_r_137_b : _GEN_9836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9838 = 8'h8a == r_count_47_io_out ? io_r_138_b : _GEN_9837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9839 = 8'h8b == r_count_47_io_out ? io_r_139_b : _GEN_9838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9840 = 8'h8c == r_count_47_io_out ? io_r_140_b : _GEN_9839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9841 = 8'h8d == r_count_47_io_out ? io_r_141_b : _GEN_9840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9842 = 8'h8e == r_count_47_io_out ? io_r_142_b : _GEN_9841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9843 = 8'h8f == r_count_47_io_out ? io_r_143_b : _GEN_9842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9844 = 8'h90 == r_count_47_io_out ? io_r_144_b : _GEN_9843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9845 = 8'h91 == r_count_47_io_out ? io_r_145_b : _GEN_9844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9846 = 8'h92 == r_count_47_io_out ? io_r_146_b : _GEN_9845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9847 = 8'h93 == r_count_47_io_out ? io_r_147_b : _GEN_9846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9848 = 8'h94 == r_count_47_io_out ? io_r_148_b : _GEN_9847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9849 = 8'h95 == r_count_47_io_out ? io_r_149_b : _GEN_9848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9850 = 8'h96 == r_count_47_io_out ? io_r_150_b : _GEN_9849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9851 = 8'h97 == r_count_47_io_out ? io_r_151_b : _GEN_9850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9852 = 8'h98 == r_count_47_io_out ? io_r_152_b : _GEN_9851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9853 = 8'h99 == r_count_47_io_out ? io_r_153_b : _GEN_9852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9854 = 8'h9a == r_count_47_io_out ? io_r_154_b : _GEN_9853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9855 = 8'h9b == r_count_47_io_out ? io_r_155_b : _GEN_9854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9856 = 8'h9c == r_count_47_io_out ? io_r_156_b : _GEN_9855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9857 = 8'h9d == r_count_47_io_out ? io_r_157_b : _GEN_9856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9858 = 8'h9e == r_count_47_io_out ? io_r_158_b : _GEN_9857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9859 = 8'h9f == r_count_47_io_out ? io_r_159_b : _GEN_9858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9860 = 8'ha0 == r_count_47_io_out ? io_r_160_b : _GEN_9859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9861 = 8'ha1 == r_count_47_io_out ? io_r_161_b : _GEN_9860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9862 = 8'ha2 == r_count_47_io_out ? io_r_162_b : _GEN_9861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9863 = 8'ha3 == r_count_47_io_out ? io_r_163_b : _GEN_9862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9864 = 8'ha4 == r_count_47_io_out ? io_r_164_b : _GEN_9863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9865 = 8'ha5 == r_count_47_io_out ? io_r_165_b : _GEN_9864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9866 = 8'ha6 == r_count_47_io_out ? io_r_166_b : _GEN_9865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9867 = 8'ha7 == r_count_47_io_out ? io_r_167_b : _GEN_9866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9868 = 8'ha8 == r_count_47_io_out ? io_r_168_b : _GEN_9867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9869 = 8'ha9 == r_count_47_io_out ? io_r_169_b : _GEN_9868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9870 = 8'haa == r_count_47_io_out ? io_r_170_b : _GEN_9869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9871 = 8'hab == r_count_47_io_out ? io_r_171_b : _GEN_9870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9872 = 8'hac == r_count_47_io_out ? io_r_172_b : _GEN_9871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9873 = 8'had == r_count_47_io_out ? io_r_173_b : _GEN_9872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9874 = 8'hae == r_count_47_io_out ? io_r_174_b : _GEN_9873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9875 = 8'haf == r_count_47_io_out ? io_r_175_b : _GEN_9874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9876 = 8'hb0 == r_count_47_io_out ? io_r_176_b : _GEN_9875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9877 = 8'hb1 == r_count_47_io_out ? io_r_177_b : _GEN_9876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9878 = 8'hb2 == r_count_47_io_out ? io_r_178_b : _GEN_9877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9879 = 8'hb3 == r_count_47_io_out ? io_r_179_b : _GEN_9878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9880 = 8'hb4 == r_count_47_io_out ? io_r_180_b : _GEN_9879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9881 = 8'hb5 == r_count_47_io_out ? io_r_181_b : _GEN_9880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9882 = 8'hb6 == r_count_47_io_out ? io_r_182_b : _GEN_9881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9883 = 8'hb7 == r_count_47_io_out ? io_r_183_b : _GEN_9882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9884 = 8'hb8 == r_count_47_io_out ? io_r_184_b : _GEN_9883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9885 = 8'hb9 == r_count_47_io_out ? io_r_185_b : _GEN_9884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9886 = 8'hba == r_count_47_io_out ? io_r_186_b : _GEN_9885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9887 = 8'hbb == r_count_47_io_out ? io_r_187_b : _GEN_9886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9888 = 8'hbc == r_count_47_io_out ? io_r_188_b : _GEN_9887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9889 = 8'hbd == r_count_47_io_out ? io_r_189_b : _GEN_9888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9890 = 8'hbe == r_count_47_io_out ? io_r_190_b : _GEN_9889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9891 = 8'hbf == r_count_47_io_out ? io_r_191_b : _GEN_9890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9892 = 8'hc0 == r_count_47_io_out ? io_r_192_b : _GEN_9891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9893 = 8'hc1 == r_count_47_io_out ? io_r_193_b : _GEN_9892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9894 = 8'hc2 == r_count_47_io_out ? io_r_194_b : _GEN_9893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9895 = 8'hc3 == r_count_47_io_out ? io_r_195_b : _GEN_9894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9896 = 8'hc4 == r_count_47_io_out ? io_r_196_b : _GEN_9895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9897 = 8'hc5 == r_count_47_io_out ? io_r_197_b : _GEN_9896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9898 = 8'hc6 == r_count_47_io_out ? io_r_198_b : _GEN_9897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9901 = 8'h1 == r_count_48_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9902 = 8'h2 == r_count_48_io_out ? io_r_2_b : _GEN_9901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9903 = 8'h3 == r_count_48_io_out ? io_r_3_b : _GEN_9902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9904 = 8'h4 == r_count_48_io_out ? io_r_4_b : _GEN_9903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9905 = 8'h5 == r_count_48_io_out ? io_r_5_b : _GEN_9904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9906 = 8'h6 == r_count_48_io_out ? io_r_6_b : _GEN_9905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9907 = 8'h7 == r_count_48_io_out ? io_r_7_b : _GEN_9906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9908 = 8'h8 == r_count_48_io_out ? io_r_8_b : _GEN_9907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9909 = 8'h9 == r_count_48_io_out ? io_r_9_b : _GEN_9908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9910 = 8'ha == r_count_48_io_out ? io_r_10_b : _GEN_9909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9911 = 8'hb == r_count_48_io_out ? io_r_11_b : _GEN_9910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9912 = 8'hc == r_count_48_io_out ? io_r_12_b : _GEN_9911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9913 = 8'hd == r_count_48_io_out ? io_r_13_b : _GEN_9912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9914 = 8'he == r_count_48_io_out ? io_r_14_b : _GEN_9913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9915 = 8'hf == r_count_48_io_out ? io_r_15_b : _GEN_9914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9916 = 8'h10 == r_count_48_io_out ? io_r_16_b : _GEN_9915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9917 = 8'h11 == r_count_48_io_out ? io_r_17_b : _GEN_9916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9918 = 8'h12 == r_count_48_io_out ? io_r_18_b : _GEN_9917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9919 = 8'h13 == r_count_48_io_out ? io_r_19_b : _GEN_9918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9920 = 8'h14 == r_count_48_io_out ? io_r_20_b : _GEN_9919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9921 = 8'h15 == r_count_48_io_out ? io_r_21_b : _GEN_9920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9922 = 8'h16 == r_count_48_io_out ? io_r_22_b : _GEN_9921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9923 = 8'h17 == r_count_48_io_out ? io_r_23_b : _GEN_9922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9924 = 8'h18 == r_count_48_io_out ? io_r_24_b : _GEN_9923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9925 = 8'h19 == r_count_48_io_out ? io_r_25_b : _GEN_9924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9926 = 8'h1a == r_count_48_io_out ? io_r_26_b : _GEN_9925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9927 = 8'h1b == r_count_48_io_out ? io_r_27_b : _GEN_9926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9928 = 8'h1c == r_count_48_io_out ? io_r_28_b : _GEN_9927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9929 = 8'h1d == r_count_48_io_out ? io_r_29_b : _GEN_9928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9930 = 8'h1e == r_count_48_io_out ? io_r_30_b : _GEN_9929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9931 = 8'h1f == r_count_48_io_out ? io_r_31_b : _GEN_9930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9932 = 8'h20 == r_count_48_io_out ? io_r_32_b : _GEN_9931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9933 = 8'h21 == r_count_48_io_out ? io_r_33_b : _GEN_9932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9934 = 8'h22 == r_count_48_io_out ? io_r_34_b : _GEN_9933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9935 = 8'h23 == r_count_48_io_out ? io_r_35_b : _GEN_9934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9936 = 8'h24 == r_count_48_io_out ? io_r_36_b : _GEN_9935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9937 = 8'h25 == r_count_48_io_out ? io_r_37_b : _GEN_9936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9938 = 8'h26 == r_count_48_io_out ? io_r_38_b : _GEN_9937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9939 = 8'h27 == r_count_48_io_out ? io_r_39_b : _GEN_9938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9940 = 8'h28 == r_count_48_io_out ? io_r_40_b : _GEN_9939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9941 = 8'h29 == r_count_48_io_out ? io_r_41_b : _GEN_9940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9942 = 8'h2a == r_count_48_io_out ? io_r_42_b : _GEN_9941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9943 = 8'h2b == r_count_48_io_out ? io_r_43_b : _GEN_9942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9944 = 8'h2c == r_count_48_io_out ? io_r_44_b : _GEN_9943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9945 = 8'h2d == r_count_48_io_out ? io_r_45_b : _GEN_9944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9946 = 8'h2e == r_count_48_io_out ? io_r_46_b : _GEN_9945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9947 = 8'h2f == r_count_48_io_out ? io_r_47_b : _GEN_9946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9948 = 8'h30 == r_count_48_io_out ? io_r_48_b : _GEN_9947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9949 = 8'h31 == r_count_48_io_out ? io_r_49_b : _GEN_9948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9950 = 8'h32 == r_count_48_io_out ? io_r_50_b : _GEN_9949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9951 = 8'h33 == r_count_48_io_out ? io_r_51_b : _GEN_9950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9952 = 8'h34 == r_count_48_io_out ? io_r_52_b : _GEN_9951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9953 = 8'h35 == r_count_48_io_out ? io_r_53_b : _GEN_9952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9954 = 8'h36 == r_count_48_io_out ? io_r_54_b : _GEN_9953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9955 = 8'h37 == r_count_48_io_out ? io_r_55_b : _GEN_9954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9956 = 8'h38 == r_count_48_io_out ? io_r_56_b : _GEN_9955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9957 = 8'h39 == r_count_48_io_out ? io_r_57_b : _GEN_9956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9958 = 8'h3a == r_count_48_io_out ? io_r_58_b : _GEN_9957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9959 = 8'h3b == r_count_48_io_out ? io_r_59_b : _GEN_9958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9960 = 8'h3c == r_count_48_io_out ? io_r_60_b : _GEN_9959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9961 = 8'h3d == r_count_48_io_out ? io_r_61_b : _GEN_9960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9962 = 8'h3e == r_count_48_io_out ? io_r_62_b : _GEN_9961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9963 = 8'h3f == r_count_48_io_out ? io_r_63_b : _GEN_9962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9964 = 8'h40 == r_count_48_io_out ? io_r_64_b : _GEN_9963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9965 = 8'h41 == r_count_48_io_out ? io_r_65_b : _GEN_9964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9966 = 8'h42 == r_count_48_io_out ? io_r_66_b : _GEN_9965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9967 = 8'h43 == r_count_48_io_out ? io_r_67_b : _GEN_9966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9968 = 8'h44 == r_count_48_io_out ? io_r_68_b : _GEN_9967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9969 = 8'h45 == r_count_48_io_out ? io_r_69_b : _GEN_9968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9970 = 8'h46 == r_count_48_io_out ? io_r_70_b : _GEN_9969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9971 = 8'h47 == r_count_48_io_out ? io_r_71_b : _GEN_9970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9972 = 8'h48 == r_count_48_io_out ? io_r_72_b : _GEN_9971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9973 = 8'h49 == r_count_48_io_out ? io_r_73_b : _GEN_9972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9974 = 8'h4a == r_count_48_io_out ? io_r_74_b : _GEN_9973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9975 = 8'h4b == r_count_48_io_out ? io_r_75_b : _GEN_9974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9976 = 8'h4c == r_count_48_io_out ? io_r_76_b : _GEN_9975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9977 = 8'h4d == r_count_48_io_out ? io_r_77_b : _GEN_9976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9978 = 8'h4e == r_count_48_io_out ? io_r_78_b : _GEN_9977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9979 = 8'h4f == r_count_48_io_out ? io_r_79_b : _GEN_9978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9980 = 8'h50 == r_count_48_io_out ? io_r_80_b : _GEN_9979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9981 = 8'h51 == r_count_48_io_out ? io_r_81_b : _GEN_9980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9982 = 8'h52 == r_count_48_io_out ? io_r_82_b : _GEN_9981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9983 = 8'h53 == r_count_48_io_out ? io_r_83_b : _GEN_9982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9984 = 8'h54 == r_count_48_io_out ? io_r_84_b : _GEN_9983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9985 = 8'h55 == r_count_48_io_out ? io_r_85_b : _GEN_9984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9986 = 8'h56 == r_count_48_io_out ? io_r_86_b : _GEN_9985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9987 = 8'h57 == r_count_48_io_out ? io_r_87_b : _GEN_9986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9988 = 8'h58 == r_count_48_io_out ? io_r_88_b : _GEN_9987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9989 = 8'h59 == r_count_48_io_out ? io_r_89_b : _GEN_9988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9990 = 8'h5a == r_count_48_io_out ? io_r_90_b : _GEN_9989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9991 = 8'h5b == r_count_48_io_out ? io_r_91_b : _GEN_9990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9992 = 8'h5c == r_count_48_io_out ? io_r_92_b : _GEN_9991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9993 = 8'h5d == r_count_48_io_out ? io_r_93_b : _GEN_9992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9994 = 8'h5e == r_count_48_io_out ? io_r_94_b : _GEN_9993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9995 = 8'h5f == r_count_48_io_out ? io_r_95_b : _GEN_9994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9996 = 8'h60 == r_count_48_io_out ? io_r_96_b : _GEN_9995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9997 = 8'h61 == r_count_48_io_out ? io_r_97_b : _GEN_9996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9998 = 8'h62 == r_count_48_io_out ? io_r_98_b : _GEN_9997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_9999 = 8'h63 == r_count_48_io_out ? io_r_99_b : _GEN_9998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10000 = 8'h64 == r_count_48_io_out ? io_r_100_b : _GEN_9999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10001 = 8'h65 == r_count_48_io_out ? io_r_101_b : _GEN_10000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10002 = 8'h66 == r_count_48_io_out ? io_r_102_b : _GEN_10001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10003 = 8'h67 == r_count_48_io_out ? io_r_103_b : _GEN_10002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10004 = 8'h68 == r_count_48_io_out ? io_r_104_b : _GEN_10003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10005 = 8'h69 == r_count_48_io_out ? io_r_105_b : _GEN_10004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10006 = 8'h6a == r_count_48_io_out ? io_r_106_b : _GEN_10005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10007 = 8'h6b == r_count_48_io_out ? io_r_107_b : _GEN_10006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10008 = 8'h6c == r_count_48_io_out ? io_r_108_b : _GEN_10007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10009 = 8'h6d == r_count_48_io_out ? io_r_109_b : _GEN_10008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10010 = 8'h6e == r_count_48_io_out ? io_r_110_b : _GEN_10009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10011 = 8'h6f == r_count_48_io_out ? io_r_111_b : _GEN_10010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10012 = 8'h70 == r_count_48_io_out ? io_r_112_b : _GEN_10011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10013 = 8'h71 == r_count_48_io_out ? io_r_113_b : _GEN_10012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10014 = 8'h72 == r_count_48_io_out ? io_r_114_b : _GEN_10013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10015 = 8'h73 == r_count_48_io_out ? io_r_115_b : _GEN_10014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10016 = 8'h74 == r_count_48_io_out ? io_r_116_b : _GEN_10015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10017 = 8'h75 == r_count_48_io_out ? io_r_117_b : _GEN_10016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10018 = 8'h76 == r_count_48_io_out ? io_r_118_b : _GEN_10017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10019 = 8'h77 == r_count_48_io_out ? io_r_119_b : _GEN_10018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10020 = 8'h78 == r_count_48_io_out ? io_r_120_b : _GEN_10019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10021 = 8'h79 == r_count_48_io_out ? io_r_121_b : _GEN_10020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10022 = 8'h7a == r_count_48_io_out ? io_r_122_b : _GEN_10021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10023 = 8'h7b == r_count_48_io_out ? io_r_123_b : _GEN_10022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10024 = 8'h7c == r_count_48_io_out ? io_r_124_b : _GEN_10023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10025 = 8'h7d == r_count_48_io_out ? io_r_125_b : _GEN_10024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10026 = 8'h7e == r_count_48_io_out ? io_r_126_b : _GEN_10025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10027 = 8'h7f == r_count_48_io_out ? io_r_127_b : _GEN_10026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10028 = 8'h80 == r_count_48_io_out ? io_r_128_b : _GEN_10027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10029 = 8'h81 == r_count_48_io_out ? io_r_129_b : _GEN_10028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10030 = 8'h82 == r_count_48_io_out ? io_r_130_b : _GEN_10029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10031 = 8'h83 == r_count_48_io_out ? io_r_131_b : _GEN_10030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10032 = 8'h84 == r_count_48_io_out ? io_r_132_b : _GEN_10031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10033 = 8'h85 == r_count_48_io_out ? io_r_133_b : _GEN_10032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10034 = 8'h86 == r_count_48_io_out ? io_r_134_b : _GEN_10033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10035 = 8'h87 == r_count_48_io_out ? io_r_135_b : _GEN_10034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10036 = 8'h88 == r_count_48_io_out ? io_r_136_b : _GEN_10035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10037 = 8'h89 == r_count_48_io_out ? io_r_137_b : _GEN_10036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10038 = 8'h8a == r_count_48_io_out ? io_r_138_b : _GEN_10037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10039 = 8'h8b == r_count_48_io_out ? io_r_139_b : _GEN_10038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10040 = 8'h8c == r_count_48_io_out ? io_r_140_b : _GEN_10039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10041 = 8'h8d == r_count_48_io_out ? io_r_141_b : _GEN_10040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10042 = 8'h8e == r_count_48_io_out ? io_r_142_b : _GEN_10041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10043 = 8'h8f == r_count_48_io_out ? io_r_143_b : _GEN_10042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10044 = 8'h90 == r_count_48_io_out ? io_r_144_b : _GEN_10043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10045 = 8'h91 == r_count_48_io_out ? io_r_145_b : _GEN_10044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10046 = 8'h92 == r_count_48_io_out ? io_r_146_b : _GEN_10045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10047 = 8'h93 == r_count_48_io_out ? io_r_147_b : _GEN_10046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10048 = 8'h94 == r_count_48_io_out ? io_r_148_b : _GEN_10047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10049 = 8'h95 == r_count_48_io_out ? io_r_149_b : _GEN_10048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10050 = 8'h96 == r_count_48_io_out ? io_r_150_b : _GEN_10049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10051 = 8'h97 == r_count_48_io_out ? io_r_151_b : _GEN_10050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10052 = 8'h98 == r_count_48_io_out ? io_r_152_b : _GEN_10051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10053 = 8'h99 == r_count_48_io_out ? io_r_153_b : _GEN_10052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10054 = 8'h9a == r_count_48_io_out ? io_r_154_b : _GEN_10053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10055 = 8'h9b == r_count_48_io_out ? io_r_155_b : _GEN_10054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10056 = 8'h9c == r_count_48_io_out ? io_r_156_b : _GEN_10055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10057 = 8'h9d == r_count_48_io_out ? io_r_157_b : _GEN_10056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10058 = 8'h9e == r_count_48_io_out ? io_r_158_b : _GEN_10057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10059 = 8'h9f == r_count_48_io_out ? io_r_159_b : _GEN_10058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10060 = 8'ha0 == r_count_48_io_out ? io_r_160_b : _GEN_10059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10061 = 8'ha1 == r_count_48_io_out ? io_r_161_b : _GEN_10060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10062 = 8'ha2 == r_count_48_io_out ? io_r_162_b : _GEN_10061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10063 = 8'ha3 == r_count_48_io_out ? io_r_163_b : _GEN_10062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10064 = 8'ha4 == r_count_48_io_out ? io_r_164_b : _GEN_10063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10065 = 8'ha5 == r_count_48_io_out ? io_r_165_b : _GEN_10064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10066 = 8'ha6 == r_count_48_io_out ? io_r_166_b : _GEN_10065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10067 = 8'ha7 == r_count_48_io_out ? io_r_167_b : _GEN_10066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10068 = 8'ha8 == r_count_48_io_out ? io_r_168_b : _GEN_10067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10069 = 8'ha9 == r_count_48_io_out ? io_r_169_b : _GEN_10068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10070 = 8'haa == r_count_48_io_out ? io_r_170_b : _GEN_10069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10071 = 8'hab == r_count_48_io_out ? io_r_171_b : _GEN_10070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10072 = 8'hac == r_count_48_io_out ? io_r_172_b : _GEN_10071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10073 = 8'had == r_count_48_io_out ? io_r_173_b : _GEN_10072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10074 = 8'hae == r_count_48_io_out ? io_r_174_b : _GEN_10073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10075 = 8'haf == r_count_48_io_out ? io_r_175_b : _GEN_10074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10076 = 8'hb0 == r_count_48_io_out ? io_r_176_b : _GEN_10075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10077 = 8'hb1 == r_count_48_io_out ? io_r_177_b : _GEN_10076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10078 = 8'hb2 == r_count_48_io_out ? io_r_178_b : _GEN_10077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10079 = 8'hb3 == r_count_48_io_out ? io_r_179_b : _GEN_10078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10080 = 8'hb4 == r_count_48_io_out ? io_r_180_b : _GEN_10079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10081 = 8'hb5 == r_count_48_io_out ? io_r_181_b : _GEN_10080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10082 = 8'hb6 == r_count_48_io_out ? io_r_182_b : _GEN_10081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10083 = 8'hb7 == r_count_48_io_out ? io_r_183_b : _GEN_10082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10084 = 8'hb8 == r_count_48_io_out ? io_r_184_b : _GEN_10083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10085 = 8'hb9 == r_count_48_io_out ? io_r_185_b : _GEN_10084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10086 = 8'hba == r_count_48_io_out ? io_r_186_b : _GEN_10085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10087 = 8'hbb == r_count_48_io_out ? io_r_187_b : _GEN_10086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10088 = 8'hbc == r_count_48_io_out ? io_r_188_b : _GEN_10087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10089 = 8'hbd == r_count_48_io_out ? io_r_189_b : _GEN_10088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10090 = 8'hbe == r_count_48_io_out ? io_r_190_b : _GEN_10089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10091 = 8'hbf == r_count_48_io_out ? io_r_191_b : _GEN_10090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10092 = 8'hc0 == r_count_48_io_out ? io_r_192_b : _GEN_10091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10093 = 8'hc1 == r_count_48_io_out ? io_r_193_b : _GEN_10092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10094 = 8'hc2 == r_count_48_io_out ? io_r_194_b : _GEN_10093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10095 = 8'hc3 == r_count_48_io_out ? io_r_195_b : _GEN_10094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10096 = 8'hc4 == r_count_48_io_out ? io_r_196_b : _GEN_10095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10097 = 8'hc5 == r_count_48_io_out ? io_r_197_b : _GEN_10096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10098 = 8'hc6 == r_count_48_io_out ? io_r_198_b : _GEN_10097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10101 = 8'h1 == r_count_49_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10102 = 8'h2 == r_count_49_io_out ? io_r_2_b : _GEN_10101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10103 = 8'h3 == r_count_49_io_out ? io_r_3_b : _GEN_10102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10104 = 8'h4 == r_count_49_io_out ? io_r_4_b : _GEN_10103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10105 = 8'h5 == r_count_49_io_out ? io_r_5_b : _GEN_10104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10106 = 8'h6 == r_count_49_io_out ? io_r_6_b : _GEN_10105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10107 = 8'h7 == r_count_49_io_out ? io_r_7_b : _GEN_10106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10108 = 8'h8 == r_count_49_io_out ? io_r_8_b : _GEN_10107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10109 = 8'h9 == r_count_49_io_out ? io_r_9_b : _GEN_10108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10110 = 8'ha == r_count_49_io_out ? io_r_10_b : _GEN_10109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10111 = 8'hb == r_count_49_io_out ? io_r_11_b : _GEN_10110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10112 = 8'hc == r_count_49_io_out ? io_r_12_b : _GEN_10111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10113 = 8'hd == r_count_49_io_out ? io_r_13_b : _GEN_10112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10114 = 8'he == r_count_49_io_out ? io_r_14_b : _GEN_10113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10115 = 8'hf == r_count_49_io_out ? io_r_15_b : _GEN_10114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10116 = 8'h10 == r_count_49_io_out ? io_r_16_b : _GEN_10115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10117 = 8'h11 == r_count_49_io_out ? io_r_17_b : _GEN_10116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10118 = 8'h12 == r_count_49_io_out ? io_r_18_b : _GEN_10117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10119 = 8'h13 == r_count_49_io_out ? io_r_19_b : _GEN_10118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10120 = 8'h14 == r_count_49_io_out ? io_r_20_b : _GEN_10119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10121 = 8'h15 == r_count_49_io_out ? io_r_21_b : _GEN_10120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10122 = 8'h16 == r_count_49_io_out ? io_r_22_b : _GEN_10121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10123 = 8'h17 == r_count_49_io_out ? io_r_23_b : _GEN_10122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10124 = 8'h18 == r_count_49_io_out ? io_r_24_b : _GEN_10123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10125 = 8'h19 == r_count_49_io_out ? io_r_25_b : _GEN_10124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10126 = 8'h1a == r_count_49_io_out ? io_r_26_b : _GEN_10125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10127 = 8'h1b == r_count_49_io_out ? io_r_27_b : _GEN_10126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10128 = 8'h1c == r_count_49_io_out ? io_r_28_b : _GEN_10127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10129 = 8'h1d == r_count_49_io_out ? io_r_29_b : _GEN_10128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10130 = 8'h1e == r_count_49_io_out ? io_r_30_b : _GEN_10129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10131 = 8'h1f == r_count_49_io_out ? io_r_31_b : _GEN_10130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10132 = 8'h20 == r_count_49_io_out ? io_r_32_b : _GEN_10131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10133 = 8'h21 == r_count_49_io_out ? io_r_33_b : _GEN_10132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10134 = 8'h22 == r_count_49_io_out ? io_r_34_b : _GEN_10133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10135 = 8'h23 == r_count_49_io_out ? io_r_35_b : _GEN_10134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10136 = 8'h24 == r_count_49_io_out ? io_r_36_b : _GEN_10135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10137 = 8'h25 == r_count_49_io_out ? io_r_37_b : _GEN_10136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10138 = 8'h26 == r_count_49_io_out ? io_r_38_b : _GEN_10137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10139 = 8'h27 == r_count_49_io_out ? io_r_39_b : _GEN_10138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10140 = 8'h28 == r_count_49_io_out ? io_r_40_b : _GEN_10139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10141 = 8'h29 == r_count_49_io_out ? io_r_41_b : _GEN_10140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10142 = 8'h2a == r_count_49_io_out ? io_r_42_b : _GEN_10141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10143 = 8'h2b == r_count_49_io_out ? io_r_43_b : _GEN_10142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10144 = 8'h2c == r_count_49_io_out ? io_r_44_b : _GEN_10143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10145 = 8'h2d == r_count_49_io_out ? io_r_45_b : _GEN_10144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10146 = 8'h2e == r_count_49_io_out ? io_r_46_b : _GEN_10145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10147 = 8'h2f == r_count_49_io_out ? io_r_47_b : _GEN_10146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10148 = 8'h30 == r_count_49_io_out ? io_r_48_b : _GEN_10147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10149 = 8'h31 == r_count_49_io_out ? io_r_49_b : _GEN_10148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10150 = 8'h32 == r_count_49_io_out ? io_r_50_b : _GEN_10149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10151 = 8'h33 == r_count_49_io_out ? io_r_51_b : _GEN_10150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10152 = 8'h34 == r_count_49_io_out ? io_r_52_b : _GEN_10151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10153 = 8'h35 == r_count_49_io_out ? io_r_53_b : _GEN_10152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10154 = 8'h36 == r_count_49_io_out ? io_r_54_b : _GEN_10153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10155 = 8'h37 == r_count_49_io_out ? io_r_55_b : _GEN_10154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10156 = 8'h38 == r_count_49_io_out ? io_r_56_b : _GEN_10155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10157 = 8'h39 == r_count_49_io_out ? io_r_57_b : _GEN_10156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10158 = 8'h3a == r_count_49_io_out ? io_r_58_b : _GEN_10157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10159 = 8'h3b == r_count_49_io_out ? io_r_59_b : _GEN_10158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10160 = 8'h3c == r_count_49_io_out ? io_r_60_b : _GEN_10159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10161 = 8'h3d == r_count_49_io_out ? io_r_61_b : _GEN_10160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10162 = 8'h3e == r_count_49_io_out ? io_r_62_b : _GEN_10161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10163 = 8'h3f == r_count_49_io_out ? io_r_63_b : _GEN_10162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10164 = 8'h40 == r_count_49_io_out ? io_r_64_b : _GEN_10163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10165 = 8'h41 == r_count_49_io_out ? io_r_65_b : _GEN_10164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10166 = 8'h42 == r_count_49_io_out ? io_r_66_b : _GEN_10165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10167 = 8'h43 == r_count_49_io_out ? io_r_67_b : _GEN_10166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10168 = 8'h44 == r_count_49_io_out ? io_r_68_b : _GEN_10167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10169 = 8'h45 == r_count_49_io_out ? io_r_69_b : _GEN_10168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10170 = 8'h46 == r_count_49_io_out ? io_r_70_b : _GEN_10169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10171 = 8'h47 == r_count_49_io_out ? io_r_71_b : _GEN_10170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10172 = 8'h48 == r_count_49_io_out ? io_r_72_b : _GEN_10171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10173 = 8'h49 == r_count_49_io_out ? io_r_73_b : _GEN_10172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10174 = 8'h4a == r_count_49_io_out ? io_r_74_b : _GEN_10173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10175 = 8'h4b == r_count_49_io_out ? io_r_75_b : _GEN_10174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10176 = 8'h4c == r_count_49_io_out ? io_r_76_b : _GEN_10175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10177 = 8'h4d == r_count_49_io_out ? io_r_77_b : _GEN_10176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10178 = 8'h4e == r_count_49_io_out ? io_r_78_b : _GEN_10177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10179 = 8'h4f == r_count_49_io_out ? io_r_79_b : _GEN_10178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10180 = 8'h50 == r_count_49_io_out ? io_r_80_b : _GEN_10179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10181 = 8'h51 == r_count_49_io_out ? io_r_81_b : _GEN_10180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10182 = 8'h52 == r_count_49_io_out ? io_r_82_b : _GEN_10181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10183 = 8'h53 == r_count_49_io_out ? io_r_83_b : _GEN_10182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10184 = 8'h54 == r_count_49_io_out ? io_r_84_b : _GEN_10183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10185 = 8'h55 == r_count_49_io_out ? io_r_85_b : _GEN_10184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10186 = 8'h56 == r_count_49_io_out ? io_r_86_b : _GEN_10185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10187 = 8'h57 == r_count_49_io_out ? io_r_87_b : _GEN_10186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10188 = 8'h58 == r_count_49_io_out ? io_r_88_b : _GEN_10187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10189 = 8'h59 == r_count_49_io_out ? io_r_89_b : _GEN_10188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10190 = 8'h5a == r_count_49_io_out ? io_r_90_b : _GEN_10189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10191 = 8'h5b == r_count_49_io_out ? io_r_91_b : _GEN_10190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10192 = 8'h5c == r_count_49_io_out ? io_r_92_b : _GEN_10191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10193 = 8'h5d == r_count_49_io_out ? io_r_93_b : _GEN_10192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10194 = 8'h5e == r_count_49_io_out ? io_r_94_b : _GEN_10193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10195 = 8'h5f == r_count_49_io_out ? io_r_95_b : _GEN_10194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10196 = 8'h60 == r_count_49_io_out ? io_r_96_b : _GEN_10195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10197 = 8'h61 == r_count_49_io_out ? io_r_97_b : _GEN_10196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10198 = 8'h62 == r_count_49_io_out ? io_r_98_b : _GEN_10197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10199 = 8'h63 == r_count_49_io_out ? io_r_99_b : _GEN_10198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10200 = 8'h64 == r_count_49_io_out ? io_r_100_b : _GEN_10199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10201 = 8'h65 == r_count_49_io_out ? io_r_101_b : _GEN_10200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10202 = 8'h66 == r_count_49_io_out ? io_r_102_b : _GEN_10201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10203 = 8'h67 == r_count_49_io_out ? io_r_103_b : _GEN_10202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10204 = 8'h68 == r_count_49_io_out ? io_r_104_b : _GEN_10203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10205 = 8'h69 == r_count_49_io_out ? io_r_105_b : _GEN_10204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10206 = 8'h6a == r_count_49_io_out ? io_r_106_b : _GEN_10205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10207 = 8'h6b == r_count_49_io_out ? io_r_107_b : _GEN_10206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10208 = 8'h6c == r_count_49_io_out ? io_r_108_b : _GEN_10207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10209 = 8'h6d == r_count_49_io_out ? io_r_109_b : _GEN_10208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10210 = 8'h6e == r_count_49_io_out ? io_r_110_b : _GEN_10209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10211 = 8'h6f == r_count_49_io_out ? io_r_111_b : _GEN_10210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10212 = 8'h70 == r_count_49_io_out ? io_r_112_b : _GEN_10211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10213 = 8'h71 == r_count_49_io_out ? io_r_113_b : _GEN_10212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10214 = 8'h72 == r_count_49_io_out ? io_r_114_b : _GEN_10213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10215 = 8'h73 == r_count_49_io_out ? io_r_115_b : _GEN_10214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10216 = 8'h74 == r_count_49_io_out ? io_r_116_b : _GEN_10215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10217 = 8'h75 == r_count_49_io_out ? io_r_117_b : _GEN_10216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10218 = 8'h76 == r_count_49_io_out ? io_r_118_b : _GEN_10217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10219 = 8'h77 == r_count_49_io_out ? io_r_119_b : _GEN_10218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10220 = 8'h78 == r_count_49_io_out ? io_r_120_b : _GEN_10219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10221 = 8'h79 == r_count_49_io_out ? io_r_121_b : _GEN_10220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10222 = 8'h7a == r_count_49_io_out ? io_r_122_b : _GEN_10221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10223 = 8'h7b == r_count_49_io_out ? io_r_123_b : _GEN_10222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10224 = 8'h7c == r_count_49_io_out ? io_r_124_b : _GEN_10223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10225 = 8'h7d == r_count_49_io_out ? io_r_125_b : _GEN_10224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10226 = 8'h7e == r_count_49_io_out ? io_r_126_b : _GEN_10225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10227 = 8'h7f == r_count_49_io_out ? io_r_127_b : _GEN_10226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10228 = 8'h80 == r_count_49_io_out ? io_r_128_b : _GEN_10227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10229 = 8'h81 == r_count_49_io_out ? io_r_129_b : _GEN_10228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10230 = 8'h82 == r_count_49_io_out ? io_r_130_b : _GEN_10229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10231 = 8'h83 == r_count_49_io_out ? io_r_131_b : _GEN_10230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10232 = 8'h84 == r_count_49_io_out ? io_r_132_b : _GEN_10231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10233 = 8'h85 == r_count_49_io_out ? io_r_133_b : _GEN_10232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10234 = 8'h86 == r_count_49_io_out ? io_r_134_b : _GEN_10233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10235 = 8'h87 == r_count_49_io_out ? io_r_135_b : _GEN_10234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10236 = 8'h88 == r_count_49_io_out ? io_r_136_b : _GEN_10235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10237 = 8'h89 == r_count_49_io_out ? io_r_137_b : _GEN_10236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10238 = 8'h8a == r_count_49_io_out ? io_r_138_b : _GEN_10237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10239 = 8'h8b == r_count_49_io_out ? io_r_139_b : _GEN_10238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10240 = 8'h8c == r_count_49_io_out ? io_r_140_b : _GEN_10239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10241 = 8'h8d == r_count_49_io_out ? io_r_141_b : _GEN_10240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10242 = 8'h8e == r_count_49_io_out ? io_r_142_b : _GEN_10241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10243 = 8'h8f == r_count_49_io_out ? io_r_143_b : _GEN_10242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10244 = 8'h90 == r_count_49_io_out ? io_r_144_b : _GEN_10243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10245 = 8'h91 == r_count_49_io_out ? io_r_145_b : _GEN_10244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10246 = 8'h92 == r_count_49_io_out ? io_r_146_b : _GEN_10245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10247 = 8'h93 == r_count_49_io_out ? io_r_147_b : _GEN_10246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10248 = 8'h94 == r_count_49_io_out ? io_r_148_b : _GEN_10247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10249 = 8'h95 == r_count_49_io_out ? io_r_149_b : _GEN_10248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10250 = 8'h96 == r_count_49_io_out ? io_r_150_b : _GEN_10249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10251 = 8'h97 == r_count_49_io_out ? io_r_151_b : _GEN_10250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10252 = 8'h98 == r_count_49_io_out ? io_r_152_b : _GEN_10251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10253 = 8'h99 == r_count_49_io_out ? io_r_153_b : _GEN_10252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10254 = 8'h9a == r_count_49_io_out ? io_r_154_b : _GEN_10253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10255 = 8'h9b == r_count_49_io_out ? io_r_155_b : _GEN_10254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10256 = 8'h9c == r_count_49_io_out ? io_r_156_b : _GEN_10255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10257 = 8'h9d == r_count_49_io_out ? io_r_157_b : _GEN_10256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10258 = 8'h9e == r_count_49_io_out ? io_r_158_b : _GEN_10257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10259 = 8'h9f == r_count_49_io_out ? io_r_159_b : _GEN_10258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10260 = 8'ha0 == r_count_49_io_out ? io_r_160_b : _GEN_10259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10261 = 8'ha1 == r_count_49_io_out ? io_r_161_b : _GEN_10260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10262 = 8'ha2 == r_count_49_io_out ? io_r_162_b : _GEN_10261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10263 = 8'ha3 == r_count_49_io_out ? io_r_163_b : _GEN_10262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10264 = 8'ha4 == r_count_49_io_out ? io_r_164_b : _GEN_10263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10265 = 8'ha5 == r_count_49_io_out ? io_r_165_b : _GEN_10264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10266 = 8'ha6 == r_count_49_io_out ? io_r_166_b : _GEN_10265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10267 = 8'ha7 == r_count_49_io_out ? io_r_167_b : _GEN_10266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10268 = 8'ha8 == r_count_49_io_out ? io_r_168_b : _GEN_10267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10269 = 8'ha9 == r_count_49_io_out ? io_r_169_b : _GEN_10268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10270 = 8'haa == r_count_49_io_out ? io_r_170_b : _GEN_10269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10271 = 8'hab == r_count_49_io_out ? io_r_171_b : _GEN_10270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10272 = 8'hac == r_count_49_io_out ? io_r_172_b : _GEN_10271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10273 = 8'had == r_count_49_io_out ? io_r_173_b : _GEN_10272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10274 = 8'hae == r_count_49_io_out ? io_r_174_b : _GEN_10273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10275 = 8'haf == r_count_49_io_out ? io_r_175_b : _GEN_10274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10276 = 8'hb0 == r_count_49_io_out ? io_r_176_b : _GEN_10275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10277 = 8'hb1 == r_count_49_io_out ? io_r_177_b : _GEN_10276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10278 = 8'hb2 == r_count_49_io_out ? io_r_178_b : _GEN_10277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10279 = 8'hb3 == r_count_49_io_out ? io_r_179_b : _GEN_10278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10280 = 8'hb4 == r_count_49_io_out ? io_r_180_b : _GEN_10279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10281 = 8'hb5 == r_count_49_io_out ? io_r_181_b : _GEN_10280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10282 = 8'hb6 == r_count_49_io_out ? io_r_182_b : _GEN_10281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10283 = 8'hb7 == r_count_49_io_out ? io_r_183_b : _GEN_10282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10284 = 8'hb8 == r_count_49_io_out ? io_r_184_b : _GEN_10283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10285 = 8'hb9 == r_count_49_io_out ? io_r_185_b : _GEN_10284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10286 = 8'hba == r_count_49_io_out ? io_r_186_b : _GEN_10285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10287 = 8'hbb == r_count_49_io_out ? io_r_187_b : _GEN_10286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10288 = 8'hbc == r_count_49_io_out ? io_r_188_b : _GEN_10287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10289 = 8'hbd == r_count_49_io_out ? io_r_189_b : _GEN_10288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10290 = 8'hbe == r_count_49_io_out ? io_r_190_b : _GEN_10289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10291 = 8'hbf == r_count_49_io_out ? io_r_191_b : _GEN_10290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10292 = 8'hc0 == r_count_49_io_out ? io_r_192_b : _GEN_10291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10293 = 8'hc1 == r_count_49_io_out ? io_r_193_b : _GEN_10292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10294 = 8'hc2 == r_count_49_io_out ? io_r_194_b : _GEN_10293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10295 = 8'hc3 == r_count_49_io_out ? io_r_195_b : _GEN_10294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10296 = 8'hc4 == r_count_49_io_out ? io_r_196_b : _GEN_10295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10297 = 8'hc5 == r_count_49_io_out ? io_r_197_b : _GEN_10296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10298 = 8'hc6 == r_count_49_io_out ? io_r_198_b : _GEN_10297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10301 = 8'h1 == r_count_50_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10302 = 8'h2 == r_count_50_io_out ? io_r_2_b : _GEN_10301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10303 = 8'h3 == r_count_50_io_out ? io_r_3_b : _GEN_10302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10304 = 8'h4 == r_count_50_io_out ? io_r_4_b : _GEN_10303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10305 = 8'h5 == r_count_50_io_out ? io_r_5_b : _GEN_10304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10306 = 8'h6 == r_count_50_io_out ? io_r_6_b : _GEN_10305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10307 = 8'h7 == r_count_50_io_out ? io_r_7_b : _GEN_10306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10308 = 8'h8 == r_count_50_io_out ? io_r_8_b : _GEN_10307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10309 = 8'h9 == r_count_50_io_out ? io_r_9_b : _GEN_10308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10310 = 8'ha == r_count_50_io_out ? io_r_10_b : _GEN_10309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10311 = 8'hb == r_count_50_io_out ? io_r_11_b : _GEN_10310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10312 = 8'hc == r_count_50_io_out ? io_r_12_b : _GEN_10311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10313 = 8'hd == r_count_50_io_out ? io_r_13_b : _GEN_10312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10314 = 8'he == r_count_50_io_out ? io_r_14_b : _GEN_10313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10315 = 8'hf == r_count_50_io_out ? io_r_15_b : _GEN_10314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10316 = 8'h10 == r_count_50_io_out ? io_r_16_b : _GEN_10315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10317 = 8'h11 == r_count_50_io_out ? io_r_17_b : _GEN_10316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10318 = 8'h12 == r_count_50_io_out ? io_r_18_b : _GEN_10317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10319 = 8'h13 == r_count_50_io_out ? io_r_19_b : _GEN_10318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10320 = 8'h14 == r_count_50_io_out ? io_r_20_b : _GEN_10319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10321 = 8'h15 == r_count_50_io_out ? io_r_21_b : _GEN_10320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10322 = 8'h16 == r_count_50_io_out ? io_r_22_b : _GEN_10321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10323 = 8'h17 == r_count_50_io_out ? io_r_23_b : _GEN_10322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10324 = 8'h18 == r_count_50_io_out ? io_r_24_b : _GEN_10323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10325 = 8'h19 == r_count_50_io_out ? io_r_25_b : _GEN_10324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10326 = 8'h1a == r_count_50_io_out ? io_r_26_b : _GEN_10325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10327 = 8'h1b == r_count_50_io_out ? io_r_27_b : _GEN_10326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10328 = 8'h1c == r_count_50_io_out ? io_r_28_b : _GEN_10327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10329 = 8'h1d == r_count_50_io_out ? io_r_29_b : _GEN_10328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10330 = 8'h1e == r_count_50_io_out ? io_r_30_b : _GEN_10329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10331 = 8'h1f == r_count_50_io_out ? io_r_31_b : _GEN_10330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10332 = 8'h20 == r_count_50_io_out ? io_r_32_b : _GEN_10331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10333 = 8'h21 == r_count_50_io_out ? io_r_33_b : _GEN_10332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10334 = 8'h22 == r_count_50_io_out ? io_r_34_b : _GEN_10333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10335 = 8'h23 == r_count_50_io_out ? io_r_35_b : _GEN_10334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10336 = 8'h24 == r_count_50_io_out ? io_r_36_b : _GEN_10335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10337 = 8'h25 == r_count_50_io_out ? io_r_37_b : _GEN_10336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10338 = 8'h26 == r_count_50_io_out ? io_r_38_b : _GEN_10337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10339 = 8'h27 == r_count_50_io_out ? io_r_39_b : _GEN_10338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10340 = 8'h28 == r_count_50_io_out ? io_r_40_b : _GEN_10339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10341 = 8'h29 == r_count_50_io_out ? io_r_41_b : _GEN_10340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10342 = 8'h2a == r_count_50_io_out ? io_r_42_b : _GEN_10341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10343 = 8'h2b == r_count_50_io_out ? io_r_43_b : _GEN_10342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10344 = 8'h2c == r_count_50_io_out ? io_r_44_b : _GEN_10343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10345 = 8'h2d == r_count_50_io_out ? io_r_45_b : _GEN_10344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10346 = 8'h2e == r_count_50_io_out ? io_r_46_b : _GEN_10345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10347 = 8'h2f == r_count_50_io_out ? io_r_47_b : _GEN_10346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10348 = 8'h30 == r_count_50_io_out ? io_r_48_b : _GEN_10347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10349 = 8'h31 == r_count_50_io_out ? io_r_49_b : _GEN_10348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10350 = 8'h32 == r_count_50_io_out ? io_r_50_b : _GEN_10349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10351 = 8'h33 == r_count_50_io_out ? io_r_51_b : _GEN_10350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10352 = 8'h34 == r_count_50_io_out ? io_r_52_b : _GEN_10351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10353 = 8'h35 == r_count_50_io_out ? io_r_53_b : _GEN_10352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10354 = 8'h36 == r_count_50_io_out ? io_r_54_b : _GEN_10353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10355 = 8'h37 == r_count_50_io_out ? io_r_55_b : _GEN_10354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10356 = 8'h38 == r_count_50_io_out ? io_r_56_b : _GEN_10355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10357 = 8'h39 == r_count_50_io_out ? io_r_57_b : _GEN_10356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10358 = 8'h3a == r_count_50_io_out ? io_r_58_b : _GEN_10357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10359 = 8'h3b == r_count_50_io_out ? io_r_59_b : _GEN_10358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10360 = 8'h3c == r_count_50_io_out ? io_r_60_b : _GEN_10359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10361 = 8'h3d == r_count_50_io_out ? io_r_61_b : _GEN_10360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10362 = 8'h3e == r_count_50_io_out ? io_r_62_b : _GEN_10361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10363 = 8'h3f == r_count_50_io_out ? io_r_63_b : _GEN_10362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10364 = 8'h40 == r_count_50_io_out ? io_r_64_b : _GEN_10363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10365 = 8'h41 == r_count_50_io_out ? io_r_65_b : _GEN_10364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10366 = 8'h42 == r_count_50_io_out ? io_r_66_b : _GEN_10365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10367 = 8'h43 == r_count_50_io_out ? io_r_67_b : _GEN_10366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10368 = 8'h44 == r_count_50_io_out ? io_r_68_b : _GEN_10367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10369 = 8'h45 == r_count_50_io_out ? io_r_69_b : _GEN_10368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10370 = 8'h46 == r_count_50_io_out ? io_r_70_b : _GEN_10369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10371 = 8'h47 == r_count_50_io_out ? io_r_71_b : _GEN_10370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10372 = 8'h48 == r_count_50_io_out ? io_r_72_b : _GEN_10371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10373 = 8'h49 == r_count_50_io_out ? io_r_73_b : _GEN_10372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10374 = 8'h4a == r_count_50_io_out ? io_r_74_b : _GEN_10373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10375 = 8'h4b == r_count_50_io_out ? io_r_75_b : _GEN_10374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10376 = 8'h4c == r_count_50_io_out ? io_r_76_b : _GEN_10375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10377 = 8'h4d == r_count_50_io_out ? io_r_77_b : _GEN_10376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10378 = 8'h4e == r_count_50_io_out ? io_r_78_b : _GEN_10377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10379 = 8'h4f == r_count_50_io_out ? io_r_79_b : _GEN_10378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10380 = 8'h50 == r_count_50_io_out ? io_r_80_b : _GEN_10379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10381 = 8'h51 == r_count_50_io_out ? io_r_81_b : _GEN_10380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10382 = 8'h52 == r_count_50_io_out ? io_r_82_b : _GEN_10381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10383 = 8'h53 == r_count_50_io_out ? io_r_83_b : _GEN_10382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10384 = 8'h54 == r_count_50_io_out ? io_r_84_b : _GEN_10383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10385 = 8'h55 == r_count_50_io_out ? io_r_85_b : _GEN_10384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10386 = 8'h56 == r_count_50_io_out ? io_r_86_b : _GEN_10385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10387 = 8'h57 == r_count_50_io_out ? io_r_87_b : _GEN_10386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10388 = 8'h58 == r_count_50_io_out ? io_r_88_b : _GEN_10387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10389 = 8'h59 == r_count_50_io_out ? io_r_89_b : _GEN_10388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10390 = 8'h5a == r_count_50_io_out ? io_r_90_b : _GEN_10389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10391 = 8'h5b == r_count_50_io_out ? io_r_91_b : _GEN_10390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10392 = 8'h5c == r_count_50_io_out ? io_r_92_b : _GEN_10391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10393 = 8'h5d == r_count_50_io_out ? io_r_93_b : _GEN_10392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10394 = 8'h5e == r_count_50_io_out ? io_r_94_b : _GEN_10393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10395 = 8'h5f == r_count_50_io_out ? io_r_95_b : _GEN_10394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10396 = 8'h60 == r_count_50_io_out ? io_r_96_b : _GEN_10395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10397 = 8'h61 == r_count_50_io_out ? io_r_97_b : _GEN_10396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10398 = 8'h62 == r_count_50_io_out ? io_r_98_b : _GEN_10397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10399 = 8'h63 == r_count_50_io_out ? io_r_99_b : _GEN_10398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10400 = 8'h64 == r_count_50_io_out ? io_r_100_b : _GEN_10399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10401 = 8'h65 == r_count_50_io_out ? io_r_101_b : _GEN_10400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10402 = 8'h66 == r_count_50_io_out ? io_r_102_b : _GEN_10401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10403 = 8'h67 == r_count_50_io_out ? io_r_103_b : _GEN_10402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10404 = 8'h68 == r_count_50_io_out ? io_r_104_b : _GEN_10403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10405 = 8'h69 == r_count_50_io_out ? io_r_105_b : _GEN_10404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10406 = 8'h6a == r_count_50_io_out ? io_r_106_b : _GEN_10405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10407 = 8'h6b == r_count_50_io_out ? io_r_107_b : _GEN_10406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10408 = 8'h6c == r_count_50_io_out ? io_r_108_b : _GEN_10407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10409 = 8'h6d == r_count_50_io_out ? io_r_109_b : _GEN_10408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10410 = 8'h6e == r_count_50_io_out ? io_r_110_b : _GEN_10409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10411 = 8'h6f == r_count_50_io_out ? io_r_111_b : _GEN_10410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10412 = 8'h70 == r_count_50_io_out ? io_r_112_b : _GEN_10411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10413 = 8'h71 == r_count_50_io_out ? io_r_113_b : _GEN_10412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10414 = 8'h72 == r_count_50_io_out ? io_r_114_b : _GEN_10413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10415 = 8'h73 == r_count_50_io_out ? io_r_115_b : _GEN_10414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10416 = 8'h74 == r_count_50_io_out ? io_r_116_b : _GEN_10415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10417 = 8'h75 == r_count_50_io_out ? io_r_117_b : _GEN_10416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10418 = 8'h76 == r_count_50_io_out ? io_r_118_b : _GEN_10417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10419 = 8'h77 == r_count_50_io_out ? io_r_119_b : _GEN_10418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10420 = 8'h78 == r_count_50_io_out ? io_r_120_b : _GEN_10419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10421 = 8'h79 == r_count_50_io_out ? io_r_121_b : _GEN_10420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10422 = 8'h7a == r_count_50_io_out ? io_r_122_b : _GEN_10421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10423 = 8'h7b == r_count_50_io_out ? io_r_123_b : _GEN_10422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10424 = 8'h7c == r_count_50_io_out ? io_r_124_b : _GEN_10423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10425 = 8'h7d == r_count_50_io_out ? io_r_125_b : _GEN_10424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10426 = 8'h7e == r_count_50_io_out ? io_r_126_b : _GEN_10425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10427 = 8'h7f == r_count_50_io_out ? io_r_127_b : _GEN_10426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10428 = 8'h80 == r_count_50_io_out ? io_r_128_b : _GEN_10427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10429 = 8'h81 == r_count_50_io_out ? io_r_129_b : _GEN_10428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10430 = 8'h82 == r_count_50_io_out ? io_r_130_b : _GEN_10429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10431 = 8'h83 == r_count_50_io_out ? io_r_131_b : _GEN_10430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10432 = 8'h84 == r_count_50_io_out ? io_r_132_b : _GEN_10431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10433 = 8'h85 == r_count_50_io_out ? io_r_133_b : _GEN_10432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10434 = 8'h86 == r_count_50_io_out ? io_r_134_b : _GEN_10433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10435 = 8'h87 == r_count_50_io_out ? io_r_135_b : _GEN_10434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10436 = 8'h88 == r_count_50_io_out ? io_r_136_b : _GEN_10435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10437 = 8'h89 == r_count_50_io_out ? io_r_137_b : _GEN_10436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10438 = 8'h8a == r_count_50_io_out ? io_r_138_b : _GEN_10437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10439 = 8'h8b == r_count_50_io_out ? io_r_139_b : _GEN_10438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10440 = 8'h8c == r_count_50_io_out ? io_r_140_b : _GEN_10439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10441 = 8'h8d == r_count_50_io_out ? io_r_141_b : _GEN_10440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10442 = 8'h8e == r_count_50_io_out ? io_r_142_b : _GEN_10441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10443 = 8'h8f == r_count_50_io_out ? io_r_143_b : _GEN_10442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10444 = 8'h90 == r_count_50_io_out ? io_r_144_b : _GEN_10443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10445 = 8'h91 == r_count_50_io_out ? io_r_145_b : _GEN_10444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10446 = 8'h92 == r_count_50_io_out ? io_r_146_b : _GEN_10445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10447 = 8'h93 == r_count_50_io_out ? io_r_147_b : _GEN_10446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10448 = 8'h94 == r_count_50_io_out ? io_r_148_b : _GEN_10447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10449 = 8'h95 == r_count_50_io_out ? io_r_149_b : _GEN_10448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10450 = 8'h96 == r_count_50_io_out ? io_r_150_b : _GEN_10449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10451 = 8'h97 == r_count_50_io_out ? io_r_151_b : _GEN_10450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10452 = 8'h98 == r_count_50_io_out ? io_r_152_b : _GEN_10451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10453 = 8'h99 == r_count_50_io_out ? io_r_153_b : _GEN_10452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10454 = 8'h9a == r_count_50_io_out ? io_r_154_b : _GEN_10453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10455 = 8'h9b == r_count_50_io_out ? io_r_155_b : _GEN_10454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10456 = 8'h9c == r_count_50_io_out ? io_r_156_b : _GEN_10455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10457 = 8'h9d == r_count_50_io_out ? io_r_157_b : _GEN_10456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10458 = 8'h9e == r_count_50_io_out ? io_r_158_b : _GEN_10457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10459 = 8'h9f == r_count_50_io_out ? io_r_159_b : _GEN_10458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10460 = 8'ha0 == r_count_50_io_out ? io_r_160_b : _GEN_10459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10461 = 8'ha1 == r_count_50_io_out ? io_r_161_b : _GEN_10460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10462 = 8'ha2 == r_count_50_io_out ? io_r_162_b : _GEN_10461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10463 = 8'ha3 == r_count_50_io_out ? io_r_163_b : _GEN_10462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10464 = 8'ha4 == r_count_50_io_out ? io_r_164_b : _GEN_10463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10465 = 8'ha5 == r_count_50_io_out ? io_r_165_b : _GEN_10464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10466 = 8'ha6 == r_count_50_io_out ? io_r_166_b : _GEN_10465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10467 = 8'ha7 == r_count_50_io_out ? io_r_167_b : _GEN_10466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10468 = 8'ha8 == r_count_50_io_out ? io_r_168_b : _GEN_10467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10469 = 8'ha9 == r_count_50_io_out ? io_r_169_b : _GEN_10468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10470 = 8'haa == r_count_50_io_out ? io_r_170_b : _GEN_10469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10471 = 8'hab == r_count_50_io_out ? io_r_171_b : _GEN_10470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10472 = 8'hac == r_count_50_io_out ? io_r_172_b : _GEN_10471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10473 = 8'had == r_count_50_io_out ? io_r_173_b : _GEN_10472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10474 = 8'hae == r_count_50_io_out ? io_r_174_b : _GEN_10473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10475 = 8'haf == r_count_50_io_out ? io_r_175_b : _GEN_10474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10476 = 8'hb0 == r_count_50_io_out ? io_r_176_b : _GEN_10475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10477 = 8'hb1 == r_count_50_io_out ? io_r_177_b : _GEN_10476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10478 = 8'hb2 == r_count_50_io_out ? io_r_178_b : _GEN_10477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10479 = 8'hb3 == r_count_50_io_out ? io_r_179_b : _GEN_10478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10480 = 8'hb4 == r_count_50_io_out ? io_r_180_b : _GEN_10479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10481 = 8'hb5 == r_count_50_io_out ? io_r_181_b : _GEN_10480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10482 = 8'hb6 == r_count_50_io_out ? io_r_182_b : _GEN_10481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10483 = 8'hb7 == r_count_50_io_out ? io_r_183_b : _GEN_10482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10484 = 8'hb8 == r_count_50_io_out ? io_r_184_b : _GEN_10483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10485 = 8'hb9 == r_count_50_io_out ? io_r_185_b : _GEN_10484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10486 = 8'hba == r_count_50_io_out ? io_r_186_b : _GEN_10485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10487 = 8'hbb == r_count_50_io_out ? io_r_187_b : _GEN_10486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10488 = 8'hbc == r_count_50_io_out ? io_r_188_b : _GEN_10487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10489 = 8'hbd == r_count_50_io_out ? io_r_189_b : _GEN_10488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10490 = 8'hbe == r_count_50_io_out ? io_r_190_b : _GEN_10489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10491 = 8'hbf == r_count_50_io_out ? io_r_191_b : _GEN_10490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10492 = 8'hc0 == r_count_50_io_out ? io_r_192_b : _GEN_10491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10493 = 8'hc1 == r_count_50_io_out ? io_r_193_b : _GEN_10492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10494 = 8'hc2 == r_count_50_io_out ? io_r_194_b : _GEN_10493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10495 = 8'hc3 == r_count_50_io_out ? io_r_195_b : _GEN_10494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10496 = 8'hc4 == r_count_50_io_out ? io_r_196_b : _GEN_10495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10497 = 8'hc5 == r_count_50_io_out ? io_r_197_b : _GEN_10496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10498 = 8'hc6 == r_count_50_io_out ? io_r_198_b : _GEN_10497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10501 = 8'h1 == r_count_51_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10502 = 8'h2 == r_count_51_io_out ? io_r_2_b : _GEN_10501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10503 = 8'h3 == r_count_51_io_out ? io_r_3_b : _GEN_10502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10504 = 8'h4 == r_count_51_io_out ? io_r_4_b : _GEN_10503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10505 = 8'h5 == r_count_51_io_out ? io_r_5_b : _GEN_10504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10506 = 8'h6 == r_count_51_io_out ? io_r_6_b : _GEN_10505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10507 = 8'h7 == r_count_51_io_out ? io_r_7_b : _GEN_10506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10508 = 8'h8 == r_count_51_io_out ? io_r_8_b : _GEN_10507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10509 = 8'h9 == r_count_51_io_out ? io_r_9_b : _GEN_10508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10510 = 8'ha == r_count_51_io_out ? io_r_10_b : _GEN_10509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10511 = 8'hb == r_count_51_io_out ? io_r_11_b : _GEN_10510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10512 = 8'hc == r_count_51_io_out ? io_r_12_b : _GEN_10511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10513 = 8'hd == r_count_51_io_out ? io_r_13_b : _GEN_10512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10514 = 8'he == r_count_51_io_out ? io_r_14_b : _GEN_10513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10515 = 8'hf == r_count_51_io_out ? io_r_15_b : _GEN_10514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10516 = 8'h10 == r_count_51_io_out ? io_r_16_b : _GEN_10515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10517 = 8'h11 == r_count_51_io_out ? io_r_17_b : _GEN_10516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10518 = 8'h12 == r_count_51_io_out ? io_r_18_b : _GEN_10517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10519 = 8'h13 == r_count_51_io_out ? io_r_19_b : _GEN_10518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10520 = 8'h14 == r_count_51_io_out ? io_r_20_b : _GEN_10519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10521 = 8'h15 == r_count_51_io_out ? io_r_21_b : _GEN_10520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10522 = 8'h16 == r_count_51_io_out ? io_r_22_b : _GEN_10521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10523 = 8'h17 == r_count_51_io_out ? io_r_23_b : _GEN_10522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10524 = 8'h18 == r_count_51_io_out ? io_r_24_b : _GEN_10523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10525 = 8'h19 == r_count_51_io_out ? io_r_25_b : _GEN_10524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10526 = 8'h1a == r_count_51_io_out ? io_r_26_b : _GEN_10525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10527 = 8'h1b == r_count_51_io_out ? io_r_27_b : _GEN_10526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10528 = 8'h1c == r_count_51_io_out ? io_r_28_b : _GEN_10527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10529 = 8'h1d == r_count_51_io_out ? io_r_29_b : _GEN_10528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10530 = 8'h1e == r_count_51_io_out ? io_r_30_b : _GEN_10529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10531 = 8'h1f == r_count_51_io_out ? io_r_31_b : _GEN_10530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10532 = 8'h20 == r_count_51_io_out ? io_r_32_b : _GEN_10531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10533 = 8'h21 == r_count_51_io_out ? io_r_33_b : _GEN_10532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10534 = 8'h22 == r_count_51_io_out ? io_r_34_b : _GEN_10533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10535 = 8'h23 == r_count_51_io_out ? io_r_35_b : _GEN_10534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10536 = 8'h24 == r_count_51_io_out ? io_r_36_b : _GEN_10535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10537 = 8'h25 == r_count_51_io_out ? io_r_37_b : _GEN_10536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10538 = 8'h26 == r_count_51_io_out ? io_r_38_b : _GEN_10537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10539 = 8'h27 == r_count_51_io_out ? io_r_39_b : _GEN_10538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10540 = 8'h28 == r_count_51_io_out ? io_r_40_b : _GEN_10539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10541 = 8'h29 == r_count_51_io_out ? io_r_41_b : _GEN_10540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10542 = 8'h2a == r_count_51_io_out ? io_r_42_b : _GEN_10541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10543 = 8'h2b == r_count_51_io_out ? io_r_43_b : _GEN_10542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10544 = 8'h2c == r_count_51_io_out ? io_r_44_b : _GEN_10543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10545 = 8'h2d == r_count_51_io_out ? io_r_45_b : _GEN_10544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10546 = 8'h2e == r_count_51_io_out ? io_r_46_b : _GEN_10545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10547 = 8'h2f == r_count_51_io_out ? io_r_47_b : _GEN_10546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10548 = 8'h30 == r_count_51_io_out ? io_r_48_b : _GEN_10547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10549 = 8'h31 == r_count_51_io_out ? io_r_49_b : _GEN_10548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10550 = 8'h32 == r_count_51_io_out ? io_r_50_b : _GEN_10549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10551 = 8'h33 == r_count_51_io_out ? io_r_51_b : _GEN_10550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10552 = 8'h34 == r_count_51_io_out ? io_r_52_b : _GEN_10551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10553 = 8'h35 == r_count_51_io_out ? io_r_53_b : _GEN_10552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10554 = 8'h36 == r_count_51_io_out ? io_r_54_b : _GEN_10553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10555 = 8'h37 == r_count_51_io_out ? io_r_55_b : _GEN_10554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10556 = 8'h38 == r_count_51_io_out ? io_r_56_b : _GEN_10555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10557 = 8'h39 == r_count_51_io_out ? io_r_57_b : _GEN_10556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10558 = 8'h3a == r_count_51_io_out ? io_r_58_b : _GEN_10557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10559 = 8'h3b == r_count_51_io_out ? io_r_59_b : _GEN_10558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10560 = 8'h3c == r_count_51_io_out ? io_r_60_b : _GEN_10559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10561 = 8'h3d == r_count_51_io_out ? io_r_61_b : _GEN_10560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10562 = 8'h3e == r_count_51_io_out ? io_r_62_b : _GEN_10561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10563 = 8'h3f == r_count_51_io_out ? io_r_63_b : _GEN_10562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10564 = 8'h40 == r_count_51_io_out ? io_r_64_b : _GEN_10563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10565 = 8'h41 == r_count_51_io_out ? io_r_65_b : _GEN_10564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10566 = 8'h42 == r_count_51_io_out ? io_r_66_b : _GEN_10565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10567 = 8'h43 == r_count_51_io_out ? io_r_67_b : _GEN_10566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10568 = 8'h44 == r_count_51_io_out ? io_r_68_b : _GEN_10567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10569 = 8'h45 == r_count_51_io_out ? io_r_69_b : _GEN_10568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10570 = 8'h46 == r_count_51_io_out ? io_r_70_b : _GEN_10569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10571 = 8'h47 == r_count_51_io_out ? io_r_71_b : _GEN_10570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10572 = 8'h48 == r_count_51_io_out ? io_r_72_b : _GEN_10571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10573 = 8'h49 == r_count_51_io_out ? io_r_73_b : _GEN_10572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10574 = 8'h4a == r_count_51_io_out ? io_r_74_b : _GEN_10573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10575 = 8'h4b == r_count_51_io_out ? io_r_75_b : _GEN_10574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10576 = 8'h4c == r_count_51_io_out ? io_r_76_b : _GEN_10575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10577 = 8'h4d == r_count_51_io_out ? io_r_77_b : _GEN_10576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10578 = 8'h4e == r_count_51_io_out ? io_r_78_b : _GEN_10577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10579 = 8'h4f == r_count_51_io_out ? io_r_79_b : _GEN_10578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10580 = 8'h50 == r_count_51_io_out ? io_r_80_b : _GEN_10579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10581 = 8'h51 == r_count_51_io_out ? io_r_81_b : _GEN_10580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10582 = 8'h52 == r_count_51_io_out ? io_r_82_b : _GEN_10581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10583 = 8'h53 == r_count_51_io_out ? io_r_83_b : _GEN_10582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10584 = 8'h54 == r_count_51_io_out ? io_r_84_b : _GEN_10583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10585 = 8'h55 == r_count_51_io_out ? io_r_85_b : _GEN_10584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10586 = 8'h56 == r_count_51_io_out ? io_r_86_b : _GEN_10585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10587 = 8'h57 == r_count_51_io_out ? io_r_87_b : _GEN_10586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10588 = 8'h58 == r_count_51_io_out ? io_r_88_b : _GEN_10587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10589 = 8'h59 == r_count_51_io_out ? io_r_89_b : _GEN_10588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10590 = 8'h5a == r_count_51_io_out ? io_r_90_b : _GEN_10589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10591 = 8'h5b == r_count_51_io_out ? io_r_91_b : _GEN_10590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10592 = 8'h5c == r_count_51_io_out ? io_r_92_b : _GEN_10591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10593 = 8'h5d == r_count_51_io_out ? io_r_93_b : _GEN_10592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10594 = 8'h5e == r_count_51_io_out ? io_r_94_b : _GEN_10593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10595 = 8'h5f == r_count_51_io_out ? io_r_95_b : _GEN_10594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10596 = 8'h60 == r_count_51_io_out ? io_r_96_b : _GEN_10595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10597 = 8'h61 == r_count_51_io_out ? io_r_97_b : _GEN_10596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10598 = 8'h62 == r_count_51_io_out ? io_r_98_b : _GEN_10597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10599 = 8'h63 == r_count_51_io_out ? io_r_99_b : _GEN_10598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10600 = 8'h64 == r_count_51_io_out ? io_r_100_b : _GEN_10599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10601 = 8'h65 == r_count_51_io_out ? io_r_101_b : _GEN_10600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10602 = 8'h66 == r_count_51_io_out ? io_r_102_b : _GEN_10601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10603 = 8'h67 == r_count_51_io_out ? io_r_103_b : _GEN_10602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10604 = 8'h68 == r_count_51_io_out ? io_r_104_b : _GEN_10603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10605 = 8'h69 == r_count_51_io_out ? io_r_105_b : _GEN_10604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10606 = 8'h6a == r_count_51_io_out ? io_r_106_b : _GEN_10605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10607 = 8'h6b == r_count_51_io_out ? io_r_107_b : _GEN_10606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10608 = 8'h6c == r_count_51_io_out ? io_r_108_b : _GEN_10607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10609 = 8'h6d == r_count_51_io_out ? io_r_109_b : _GEN_10608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10610 = 8'h6e == r_count_51_io_out ? io_r_110_b : _GEN_10609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10611 = 8'h6f == r_count_51_io_out ? io_r_111_b : _GEN_10610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10612 = 8'h70 == r_count_51_io_out ? io_r_112_b : _GEN_10611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10613 = 8'h71 == r_count_51_io_out ? io_r_113_b : _GEN_10612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10614 = 8'h72 == r_count_51_io_out ? io_r_114_b : _GEN_10613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10615 = 8'h73 == r_count_51_io_out ? io_r_115_b : _GEN_10614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10616 = 8'h74 == r_count_51_io_out ? io_r_116_b : _GEN_10615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10617 = 8'h75 == r_count_51_io_out ? io_r_117_b : _GEN_10616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10618 = 8'h76 == r_count_51_io_out ? io_r_118_b : _GEN_10617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10619 = 8'h77 == r_count_51_io_out ? io_r_119_b : _GEN_10618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10620 = 8'h78 == r_count_51_io_out ? io_r_120_b : _GEN_10619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10621 = 8'h79 == r_count_51_io_out ? io_r_121_b : _GEN_10620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10622 = 8'h7a == r_count_51_io_out ? io_r_122_b : _GEN_10621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10623 = 8'h7b == r_count_51_io_out ? io_r_123_b : _GEN_10622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10624 = 8'h7c == r_count_51_io_out ? io_r_124_b : _GEN_10623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10625 = 8'h7d == r_count_51_io_out ? io_r_125_b : _GEN_10624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10626 = 8'h7e == r_count_51_io_out ? io_r_126_b : _GEN_10625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10627 = 8'h7f == r_count_51_io_out ? io_r_127_b : _GEN_10626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10628 = 8'h80 == r_count_51_io_out ? io_r_128_b : _GEN_10627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10629 = 8'h81 == r_count_51_io_out ? io_r_129_b : _GEN_10628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10630 = 8'h82 == r_count_51_io_out ? io_r_130_b : _GEN_10629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10631 = 8'h83 == r_count_51_io_out ? io_r_131_b : _GEN_10630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10632 = 8'h84 == r_count_51_io_out ? io_r_132_b : _GEN_10631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10633 = 8'h85 == r_count_51_io_out ? io_r_133_b : _GEN_10632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10634 = 8'h86 == r_count_51_io_out ? io_r_134_b : _GEN_10633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10635 = 8'h87 == r_count_51_io_out ? io_r_135_b : _GEN_10634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10636 = 8'h88 == r_count_51_io_out ? io_r_136_b : _GEN_10635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10637 = 8'h89 == r_count_51_io_out ? io_r_137_b : _GEN_10636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10638 = 8'h8a == r_count_51_io_out ? io_r_138_b : _GEN_10637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10639 = 8'h8b == r_count_51_io_out ? io_r_139_b : _GEN_10638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10640 = 8'h8c == r_count_51_io_out ? io_r_140_b : _GEN_10639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10641 = 8'h8d == r_count_51_io_out ? io_r_141_b : _GEN_10640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10642 = 8'h8e == r_count_51_io_out ? io_r_142_b : _GEN_10641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10643 = 8'h8f == r_count_51_io_out ? io_r_143_b : _GEN_10642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10644 = 8'h90 == r_count_51_io_out ? io_r_144_b : _GEN_10643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10645 = 8'h91 == r_count_51_io_out ? io_r_145_b : _GEN_10644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10646 = 8'h92 == r_count_51_io_out ? io_r_146_b : _GEN_10645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10647 = 8'h93 == r_count_51_io_out ? io_r_147_b : _GEN_10646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10648 = 8'h94 == r_count_51_io_out ? io_r_148_b : _GEN_10647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10649 = 8'h95 == r_count_51_io_out ? io_r_149_b : _GEN_10648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10650 = 8'h96 == r_count_51_io_out ? io_r_150_b : _GEN_10649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10651 = 8'h97 == r_count_51_io_out ? io_r_151_b : _GEN_10650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10652 = 8'h98 == r_count_51_io_out ? io_r_152_b : _GEN_10651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10653 = 8'h99 == r_count_51_io_out ? io_r_153_b : _GEN_10652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10654 = 8'h9a == r_count_51_io_out ? io_r_154_b : _GEN_10653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10655 = 8'h9b == r_count_51_io_out ? io_r_155_b : _GEN_10654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10656 = 8'h9c == r_count_51_io_out ? io_r_156_b : _GEN_10655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10657 = 8'h9d == r_count_51_io_out ? io_r_157_b : _GEN_10656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10658 = 8'h9e == r_count_51_io_out ? io_r_158_b : _GEN_10657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10659 = 8'h9f == r_count_51_io_out ? io_r_159_b : _GEN_10658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10660 = 8'ha0 == r_count_51_io_out ? io_r_160_b : _GEN_10659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10661 = 8'ha1 == r_count_51_io_out ? io_r_161_b : _GEN_10660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10662 = 8'ha2 == r_count_51_io_out ? io_r_162_b : _GEN_10661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10663 = 8'ha3 == r_count_51_io_out ? io_r_163_b : _GEN_10662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10664 = 8'ha4 == r_count_51_io_out ? io_r_164_b : _GEN_10663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10665 = 8'ha5 == r_count_51_io_out ? io_r_165_b : _GEN_10664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10666 = 8'ha6 == r_count_51_io_out ? io_r_166_b : _GEN_10665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10667 = 8'ha7 == r_count_51_io_out ? io_r_167_b : _GEN_10666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10668 = 8'ha8 == r_count_51_io_out ? io_r_168_b : _GEN_10667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10669 = 8'ha9 == r_count_51_io_out ? io_r_169_b : _GEN_10668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10670 = 8'haa == r_count_51_io_out ? io_r_170_b : _GEN_10669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10671 = 8'hab == r_count_51_io_out ? io_r_171_b : _GEN_10670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10672 = 8'hac == r_count_51_io_out ? io_r_172_b : _GEN_10671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10673 = 8'had == r_count_51_io_out ? io_r_173_b : _GEN_10672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10674 = 8'hae == r_count_51_io_out ? io_r_174_b : _GEN_10673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10675 = 8'haf == r_count_51_io_out ? io_r_175_b : _GEN_10674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10676 = 8'hb0 == r_count_51_io_out ? io_r_176_b : _GEN_10675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10677 = 8'hb1 == r_count_51_io_out ? io_r_177_b : _GEN_10676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10678 = 8'hb2 == r_count_51_io_out ? io_r_178_b : _GEN_10677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10679 = 8'hb3 == r_count_51_io_out ? io_r_179_b : _GEN_10678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10680 = 8'hb4 == r_count_51_io_out ? io_r_180_b : _GEN_10679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10681 = 8'hb5 == r_count_51_io_out ? io_r_181_b : _GEN_10680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10682 = 8'hb6 == r_count_51_io_out ? io_r_182_b : _GEN_10681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10683 = 8'hb7 == r_count_51_io_out ? io_r_183_b : _GEN_10682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10684 = 8'hb8 == r_count_51_io_out ? io_r_184_b : _GEN_10683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10685 = 8'hb9 == r_count_51_io_out ? io_r_185_b : _GEN_10684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10686 = 8'hba == r_count_51_io_out ? io_r_186_b : _GEN_10685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10687 = 8'hbb == r_count_51_io_out ? io_r_187_b : _GEN_10686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10688 = 8'hbc == r_count_51_io_out ? io_r_188_b : _GEN_10687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10689 = 8'hbd == r_count_51_io_out ? io_r_189_b : _GEN_10688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10690 = 8'hbe == r_count_51_io_out ? io_r_190_b : _GEN_10689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10691 = 8'hbf == r_count_51_io_out ? io_r_191_b : _GEN_10690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10692 = 8'hc0 == r_count_51_io_out ? io_r_192_b : _GEN_10691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10693 = 8'hc1 == r_count_51_io_out ? io_r_193_b : _GEN_10692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10694 = 8'hc2 == r_count_51_io_out ? io_r_194_b : _GEN_10693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10695 = 8'hc3 == r_count_51_io_out ? io_r_195_b : _GEN_10694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10696 = 8'hc4 == r_count_51_io_out ? io_r_196_b : _GEN_10695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10697 = 8'hc5 == r_count_51_io_out ? io_r_197_b : _GEN_10696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10698 = 8'hc6 == r_count_51_io_out ? io_r_198_b : _GEN_10697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10701 = 8'h1 == r_count_52_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10702 = 8'h2 == r_count_52_io_out ? io_r_2_b : _GEN_10701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10703 = 8'h3 == r_count_52_io_out ? io_r_3_b : _GEN_10702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10704 = 8'h4 == r_count_52_io_out ? io_r_4_b : _GEN_10703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10705 = 8'h5 == r_count_52_io_out ? io_r_5_b : _GEN_10704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10706 = 8'h6 == r_count_52_io_out ? io_r_6_b : _GEN_10705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10707 = 8'h7 == r_count_52_io_out ? io_r_7_b : _GEN_10706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10708 = 8'h8 == r_count_52_io_out ? io_r_8_b : _GEN_10707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10709 = 8'h9 == r_count_52_io_out ? io_r_9_b : _GEN_10708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10710 = 8'ha == r_count_52_io_out ? io_r_10_b : _GEN_10709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10711 = 8'hb == r_count_52_io_out ? io_r_11_b : _GEN_10710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10712 = 8'hc == r_count_52_io_out ? io_r_12_b : _GEN_10711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10713 = 8'hd == r_count_52_io_out ? io_r_13_b : _GEN_10712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10714 = 8'he == r_count_52_io_out ? io_r_14_b : _GEN_10713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10715 = 8'hf == r_count_52_io_out ? io_r_15_b : _GEN_10714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10716 = 8'h10 == r_count_52_io_out ? io_r_16_b : _GEN_10715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10717 = 8'h11 == r_count_52_io_out ? io_r_17_b : _GEN_10716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10718 = 8'h12 == r_count_52_io_out ? io_r_18_b : _GEN_10717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10719 = 8'h13 == r_count_52_io_out ? io_r_19_b : _GEN_10718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10720 = 8'h14 == r_count_52_io_out ? io_r_20_b : _GEN_10719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10721 = 8'h15 == r_count_52_io_out ? io_r_21_b : _GEN_10720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10722 = 8'h16 == r_count_52_io_out ? io_r_22_b : _GEN_10721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10723 = 8'h17 == r_count_52_io_out ? io_r_23_b : _GEN_10722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10724 = 8'h18 == r_count_52_io_out ? io_r_24_b : _GEN_10723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10725 = 8'h19 == r_count_52_io_out ? io_r_25_b : _GEN_10724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10726 = 8'h1a == r_count_52_io_out ? io_r_26_b : _GEN_10725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10727 = 8'h1b == r_count_52_io_out ? io_r_27_b : _GEN_10726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10728 = 8'h1c == r_count_52_io_out ? io_r_28_b : _GEN_10727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10729 = 8'h1d == r_count_52_io_out ? io_r_29_b : _GEN_10728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10730 = 8'h1e == r_count_52_io_out ? io_r_30_b : _GEN_10729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10731 = 8'h1f == r_count_52_io_out ? io_r_31_b : _GEN_10730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10732 = 8'h20 == r_count_52_io_out ? io_r_32_b : _GEN_10731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10733 = 8'h21 == r_count_52_io_out ? io_r_33_b : _GEN_10732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10734 = 8'h22 == r_count_52_io_out ? io_r_34_b : _GEN_10733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10735 = 8'h23 == r_count_52_io_out ? io_r_35_b : _GEN_10734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10736 = 8'h24 == r_count_52_io_out ? io_r_36_b : _GEN_10735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10737 = 8'h25 == r_count_52_io_out ? io_r_37_b : _GEN_10736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10738 = 8'h26 == r_count_52_io_out ? io_r_38_b : _GEN_10737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10739 = 8'h27 == r_count_52_io_out ? io_r_39_b : _GEN_10738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10740 = 8'h28 == r_count_52_io_out ? io_r_40_b : _GEN_10739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10741 = 8'h29 == r_count_52_io_out ? io_r_41_b : _GEN_10740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10742 = 8'h2a == r_count_52_io_out ? io_r_42_b : _GEN_10741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10743 = 8'h2b == r_count_52_io_out ? io_r_43_b : _GEN_10742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10744 = 8'h2c == r_count_52_io_out ? io_r_44_b : _GEN_10743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10745 = 8'h2d == r_count_52_io_out ? io_r_45_b : _GEN_10744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10746 = 8'h2e == r_count_52_io_out ? io_r_46_b : _GEN_10745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10747 = 8'h2f == r_count_52_io_out ? io_r_47_b : _GEN_10746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10748 = 8'h30 == r_count_52_io_out ? io_r_48_b : _GEN_10747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10749 = 8'h31 == r_count_52_io_out ? io_r_49_b : _GEN_10748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10750 = 8'h32 == r_count_52_io_out ? io_r_50_b : _GEN_10749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10751 = 8'h33 == r_count_52_io_out ? io_r_51_b : _GEN_10750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10752 = 8'h34 == r_count_52_io_out ? io_r_52_b : _GEN_10751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10753 = 8'h35 == r_count_52_io_out ? io_r_53_b : _GEN_10752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10754 = 8'h36 == r_count_52_io_out ? io_r_54_b : _GEN_10753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10755 = 8'h37 == r_count_52_io_out ? io_r_55_b : _GEN_10754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10756 = 8'h38 == r_count_52_io_out ? io_r_56_b : _GEN_10755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10757 = 8'h39 == r_count_52_io_out ? io_r_57_b : _GEN_10756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10758 = 8'h3a == r_count_52_io_out ? io_r_58_b : _GEN_10757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10759 = 8'h3b == r_count_52_io_out ? io_r_59_b : _GEN_10758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10760 = 8'h3c == r_count_52_io_out ? io_r_60_b : _GEN_10759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10761 = 8'h3d == r_count_52_io_out ? io_r_61_b : _GEN_10760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10762 = 8'h3e == r_count_52_io_out ? io_r_62_b : _GEN_10761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10763 = 8'h3f == r_count_52_io_out ? io_r_63_b : _GEN_10762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10764 = 8'h40 == r_count_52_io_out ? io_r_64_b : _GEN_10763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10765 = 8'h41 == r_count_52_io_out ? io_r_65_b : _GEN_10764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10766 = 8'h42 == r_count_52_io_out ? io_r_66_b : _GEN_10765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10767 = 8'h43 == r_count_52_io_out ? io_r_67_b : _GEN_10766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10768 = 8'h44 == r_count_52_io_out ? io_r_68_b : _GEN_10767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10769 = 8'h45 == r_count_52_io_out ? io_r_69_b : _GEN_10768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10770 = 8'h46 == r_count_52_io_out ? io_r_70_b : _GEN_10769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10771 = 8'h47 == r_count_52_io_out ? io_r_71_b : _GEN_10770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10772 = 8'h48 == r_count_52_io_out ? io_r_72_b : _GEN_10771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10773 = 8'h49 == r_count_52_io_out ? io_r_73_b : _GEN_10772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10774 = 8'h4a == r_count_52_io_out ? io_r_74_b : _GEN_10773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10775 = 8'h4b == r_count_52_io_out ? io_r_75_b : _GEN_10774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10776 = 8'h4c == r_count_52_io_out ? io_r_76_b : _GEN_10775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10777 = 8'h4d == r_count_52_io_out ? io_r_77_b : _GEN_10776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10778 = 8'h4e == r_count_52_io_out ? io_r_78_b : _GEN_10777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10779 = 8'h4f == r_count_52_io_out ? io_r_79_b : _GEN_10778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10780 = 8'h50 == r_count_52_io_out ? io_r_80_b : _GEN_10779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10781 = 8'h51 == r_count_52_io_out ? io_r_81_b : _GEN_10780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10782 = 8'h52 == r_count_52_io_out ? io_r_82_b : _GEN_10781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10783 = 8'h53 == r_count_52_io_out ? io_r_83_b : _GEN_10782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10784 = 8'h54 == r_count_52_io_out ? io_r_84_b : _GEN_10783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10785 = 8'h55 == r_count_52_io_out ? io_r_85_b : _GEN_10784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10786 = 8'h56 == r_count_52_io_out ? io_r_86_b : _GEN_10785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10787 = 8'h57 == r_count_52_io_out ? io_r_87_b : _GEN_10786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10788 = 8'h58 == r_count_52_io_out ? io_r_88_b : _GEN_10787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10789 = 8'h59 == r_count_52_io_out ? io_r_89_b : _GEN_10788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10790 = 8'h5a == r_count_52_io_out ? io_r_90_b : _GEN_10789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10791 = 8'h5b == r_count_52_io_out ? io_r_91_b : _GEN_10790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10792 = 8'h5c == r_count_52_io_out ? io_r_92_b : _GEN_10791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10793 = 8'h5d == r_count_52_io_out ? io_r_93_b : _GEN_10792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10794 = 8'h5e == r_count_52_io_out ? io_r_94_b : _GEN_10793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10795 = 8'h5f == r_count_52_io_out ? io_r_95_b : _GEN_10794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10796 = 8'h60 == r_count_52_io_out ? io_r_96_b : _GEN_10795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10797 = 8'h61 == r_count_52_io_out ? io_r_97_b : _GEN_10796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10798 = 8'h62 == r_count_52_io_out ? io_r_98_b : _GEN_10797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10799 = 8'h63 == r_count_52_io_out ? io_r_99_b : _GEN_10798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10800 = 8'h64 == r_count_52_io_out ? io_r_100_b : _GEN_10799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10801 = 8'h65 == r_count_52_io_out ? io_r_101_b : _GEN_10800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10802 = 8'h66 == r_count_52_io_out ? io_r_102_b : _GEN_10801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10803 = 8'h67 == r_count_52_io_out ? io_r_103_b : _GEN_10802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10804 = 8'h68 == r_count_52_io_out ? io_r_104_b : _GEN_10803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10805 = 8'h69 == r_count_52_io_out ? io_r_105_b : _GEN_10804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10806 = 8'h6a == r_count_52_io_out ? io_r_106_b : _GEN_10805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10807 = 8'h6b == r_count_52_io_out ? io_r_107_b : _GEN_10806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10808 = 8'h6c == r_count_52_io_out ? io_r_108_b : _GEN_10807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10809 = 8'h6d == r_count_52_io_out ? io_r_109_b : _GEN_10808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10810 = 8'h6e == r_count_52_io_out ? io_r_110_b : _GEN_10809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10811 = 8'h6f == r_count_52_io_out ? io_r_111_b : _GEN_10810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10812 = 8'h70 == r_count_52_io_out ? io_r_112_b : _GEN_10811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10813 = 8'h71 == r_count_52_io_out ? io_r_113_b : _GEN_10812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10814 = 8'h72 == r_count_52_io_out ? io_r_114_b : _GEN_10813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10815 = 8'h73 == r_count_52_io_out ? io_r_115_b : _GEN_10814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10816 = 8'h74 == r_count_52_io_out ? io_r_116_b : _GEN_10815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10817 = 8'h75 == r_count_52_io_out ? io_r_117_b : _GEN_10816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10818 = 8'h76 == r_count_52_io_out ? io_r_118_b : _GEN_10817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10819 = 8'h77 == r_count_52_io_out ? io_r_119_b : _GEN_10818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10820 = 8'h78 == r_count_52_io_out ? io_r_120_b : _GEN_10819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10821 = 8'h79 == r_count_52_io_out ? io_r_121_b : _GEN_10820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10822 = 8'h7a == r_count_52_io_out ? io_r_122_b : _GEN_10821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10823 = 8'h7b == r_count_52_io_out ? io_r_123_b : _GEN_10822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10824 = 8'h7c == r_count_52_io_out ? io_r_124_b : _GEN_10823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10825 = 8'h7d == r_count_52_io_out ? io_r_125_b : _GEN_10824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10826 = 8'h7e == r_count_52_io_out ? io_r_126_b : _GEN_10825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10827 = 8'h7f == r_count_52_io_out ? io_r_127_b : _GEN_10826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10828 = 8'h80 == r_count_52_io_out ? io_r_128_b : _GEN_10827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10829 = 8'h81 == r_count_52_io_out ? io_r_129_b : _GEN_10828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10830 = 8'h82 == r_count_52_io_out ? io_r_130_b : _GEN_10829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10831 = 8'h83 == r_count_52_io_out ? io_r_131_b : _GEN_10830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10832 = 8'h84 == r_count_52_io_out ? io_r_132_b : _GEN_10831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10833 = 8'h85 == r_count_52_io_out ? io_r_133_b : _GEN_10832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10834 = 8'h86 == r_count_52_io_out ? io_r_134_b : _GEN_10833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10835 = 8'h87 == r_count_52_io_out ? io_r_135_b : _GEN_10834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10836 = 8'h88 == r_count_52_io_out ? io_r_136_b : _GEN_10835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10837 = 8'h89 == r_count_52_io_out ? io_r_137_b : _GEN_10836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10838 = 8'h8a == r_count_52_io_out ? io_r_138_b : _GEN_10837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10839 = 8'h8b == r_count_52_io_out ? io_r_139_b : _GEN_10838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10840 = 8'h8c == r_count_52_io_out ? io_r_140_b : _GEN_10839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10841 = 8'h8d == r_count_52_io_out ? io_r_141_b : _GEN_10840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10842 = 8'h8e == r_count_52_io_out ? io_r_142_b : _GEN_10841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10843 = 8'h8f == r_count_52_io_out ? io_r_143_b : _GEN_10842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10844 = 8'h90 == r_count_52_io_out ? io_r_144_b : _GEN_10843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10845 = 8'h91 == r_count_52_io_out ? io_r_145_b : _GEN_10844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10846 = 8'h92 == r_count_52_io_out ? io_r_146_b : _GEN_10845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10847 = 8'h93 == r_count_52_io_out ? io_r_147_b : _GEN_10846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10848 = 8'h94 == r_count_52_io_out ? io_r_148_b : _GEN_10847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10849 = 8'h95 == r_count_52_io_out ? io_r_149_b : _GEN_10848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10850 = 8'h96 == r_count_52_io_out ? io_r_150_b : _GEN_10849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10851 = 8'h97 == r_count_52_io_out ? io_r_151_b : _GEN_10850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10852 = 8'h98 == r_count_52_io_out ? io_r_152_b : _GEN_10851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10853 = 8'h99 == r_count_52_io_out ? io_r_153_b : _GEN_10852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10854 = 8'h9a == r_count_52_io_out ? io_r_154_b : _GEN_10853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10855 = 8'h9b == r_count_52_io_out ? io_r_155_b : _GEN_10854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10856 = 8'h9c == r_count_52_io_out ? io_r_156_b : _GEN_10855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10857 = 8'h9d == r_count_52_io_out ? io_r_157_b : _GEN_10856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10858 = 8'h9e == r_count_52_io_out ? io_r_158_b : _GEN_10857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10859 = 8'h9f == r_count_52_io_out ? io_r_159_b : _GEN_10858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10860 = 8'ha0 == r_count_52_io_out ? io_r_160_b : _GEN_10859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10861 = 8'ha1 == r_count_52_io_out ? io_r_161_b : _GEN_10860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10862 = 8'ha2 == r_count_52_io_out ? io_r_162_b : _GEN_10861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10863 = 8'ha3 == r_count_52_io_out ? io_r_163_b : _GEN_10862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10864 = 8'ha4 == r_count_52_io_out ? io_r_164_b : _GEN_10863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10865 = 8'ha5 == r_count_52_io_out ? io_r_165_b : _GEN_10864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10866 = 8'ha6 == r_count_52_io_out ? io_r_166_b : _GEN_10865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10867 = 8'ha7 == r_count_52_io_out ? io_r_167_b : _GEN_10866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10868 = 8'ha8 == r_count_52_io_out ? io_r_168_b : _GEN_10867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10869 = 8'ha9 == r_count_52_io_out ? io_r_169_b : _GEN_10868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10870 = 8'haa == r_count_52_io_out ? io_r_170_b : _GEN_10869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10871 = 8'hab == r_count_52_io_out ? io_r_171_b : _GEN_10870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10872 = 8'hac == r_count_52_io_out ? io_r_172_b : _GEN_10871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10873 = 8'had == r_count_52_io_out ? io_r_173_b : _GEN_10872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10874 = 8'hae == r_count_52_io_out ? io_r_174_b : _GEN_10873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10875 = 8'haf == r_count_52_io_out ? io_r_175_b : _GEN_10874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10876 = 8'hb0 == r_count_52_io_out ? io_r_176_b : _GEN_10875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10877 = 8'hb1 == r_count_52_io_out ? io_r_177_b : _GEN_10876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10878 = 8'hb2 == r_count_52_io_out ? io_r_178_b : _GEN_10877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10879 = 8'hb3 == r_count_52_io_out ? io_r_179_b : _GEN_10878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10880 = 8'hb4 == r_count_52_io_out ? io_r_180_b : _GEN_10879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10881 = 8'hb5 == r_count_52_io_out ? io_r_181_b : _GEN_10880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10882 = 8'hb6 == r_count_52_io_out ? io_r_182_b : _GEN_10881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10883 = 8'hb7 == r_count_52_io_out ? io_r_183_b : _GEN_10882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10884 = 8'hb8 == r_count_52_io_out ? io_r_184_b : _GEN_10883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10885 = 8'hb9 == r_count_52_io_out ? io_r_185_b : _GEN_10884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10886 = 8'hba == r_count_52_io_out ? io_r_186_b : _GEN_10885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10887 = 8'hbb == r_count_52_io_out ? io_r_187_b : _GEN_10886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10888 = 8'hbc == r_count_52_io_out ? io_r_188_b : _GEN_10887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10889 = 8'hbd == r_count_52_io_out ? io_r_189_b : _GEN_10888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10890 = 8'hbe == r_count_52_io_out ? io_r_190_b : _GEN_10889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10891 = 8'hbf == r_count_52_io_out ? io_r_191_b : _GEN_10890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10892 = 8'hc0 == r_count_52_io_out ? io_r_192_b : _GEN_10891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10893 = 8'hc1 == r_count_52_io_out ? io_r_193_b : _GEN_10892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10894 = 8'hc2 == r_count_52_io_out ? io_r_194_b : _GEN_10893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10895 = 8'hc3 == r_count_52_io_out ? io_r_195_b : _GEN_10894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10896 = 8'hc4 == r_count_52_io_out ? io_r_196_b : _GEN_10895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10897 = 8'hc5 == r_count_52_io_out ? io_r_197_b : _GEN_10896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10898 = 8'hc6 == r_count_52_io_out ? io_r_198_b : _GEN_10897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10901 = 8'h1 == r_count_53_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10902 = 8'h2 == r_count_53_io_out ? io_r_2_b : _GEN_10901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10903 = 8'h3 == r_count_53_io_out ? io_r_3_b : _GEN_10902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10904 = 8'h4 == r_count_53_io_out ? io_r_4_b : _GEN_10903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10905 = 8'h5 == r_count_53_io_out ? io_r_5_b : _GEN_10904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10906 = 8'h6 == r_count_53_io_out ? io_r_6_b : _GEN_10905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10907 = 8'h7 == r_count_53_io_out ? io_r_7_b : _GEN_10906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10908 = 8'h8 == r_count_53_io_out ? io_r_8_b : _GEN_10907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10909 = 8'h9 == r_count_53_io_out ? io_r_9_b : _GEN_10908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10910 = 8'ha == r_count_53_io_out ? io_r_10_b : _GEN_10909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10911 = 8'hb == r_count_53_io_out ? io_r_11_b : _GEN_10910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10912 = 8'hc == r_count_53_io_out ? io_r_12_b : _GEN_10911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10913 = 8'hd == r_count_53_io_out ? io_r_13_b : _GEN_10912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10914 = 8'he == r_count_53_io_out ? io_r_14_b : _GEN_10913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10915 = 8'hf == r_count_53_io_out ? io_r_15_b : _GEN_10914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10916 = 8'h10 == r_count_53_io_out ? io_r_16_b : _GEN_10915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10917 = 8'h11 == r_count_53_io_out ? io_r_17_b : _GEN_10916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10918 = 8'h12 == r_count_53_io_out ? io_r_18_b : _GEN_10917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10919 = 8'h13 == r_count_53_io_out ? io_r_19_b : _GEN_10918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10920 = 8'h14 == r_count_53_io_out ? io_r_20_b : _GEN_10919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10921 = 8'h15 == r_count_53_io_out ? io_r_21_b : _GEN_10920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10922 = 8'h16 == r_count_53_io_out ? io_r_22_b : _GEN_10921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10923 = 8'h17 == r_count_53_io_out ? io_r_23_b : _GEN_10922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10924 = 8'h18 == r_count_53_io_out ? io_r_24_b : _GEN_10923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10925 = 8'h19 == r_count_53_io_out ? io_r_25_b : _GEN_10924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10926 = 8'h1a == r_count_53_io_out ? io_r_26_b : _GEN_10925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10927 = 8'h1b == r_count_53_io_out ? io_r_27_b : _GEN_10926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10928 = 8'h1c == r_count_53_io_out ? io_r_28_b : _GEN_10927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10929 = 8'h1d == r_count_53_io_out ? io_r_29_b : _GEN_10928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10930 = 8'h1e == r_count_53_io_out ? io_r_30_b : _GEN_10929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10931 = 8'h1f == r_count_53_io_out ? io_r_31_b : _GEN_10930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10932 = 8'h20 == r_count_53_io_out ? io_r_32_b : _GEN_10931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10933 = 8'h21 == r_count_53_io_out ? io_r_33_b : _GEN_10932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10934 = 8'h22 == r_count_53_io_out ? io_r_34_b : _GEN_10933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10935 = 8'h23 == r_count_53_io_out ? io_r_35_b : _GEN_10934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10936 = 8'h24 == r_count_53_io_out ? io_r_36_b : _GEN_10935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10937 = 8'h25 == r_count_53_io_out ? io_r_37_b : _GEN_10936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10938 = 8'h26 == r_count_53_io_out ? io_r_38_b : _GEN_10937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10939 = 8'h27 == r_count_53_io_out ? io_r_39_b : _GEN_10938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10940 = 8'h28 == r_count_53_io_out ? io_r_40_b : _GEN_10939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10941 = 8'h29 == r_count_53_io_out ? io_r_41_b : _GEN_10940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10942 = 8'h2a == r_count_53_io_out ? io_r_42_b : _GEN_10941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10943 = 8'h2b == r_count_53_io_out ? io_r_43_b : _GEN_10942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10944 = 8'h2c == r_count_53_io_out ? io_r_44_b : _GEN_10943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10945 = 8'h2d == r_count_53_io_out ? io_r_45_b : _GEN_10944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10946 = 8'h2e == r_count_53_io_out ? io_r_46_b : _GEN_10945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10947 = 8'h2f == r_count_53_io_out ? io_r_47_b : _GEN_10946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10948 = 8'h30 == r_count_53_io_out ? io_r_48_b : _GEN_10947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10949 = 8'h31 == r_count_53_io_out ? io_r_49_b : _GEN_10948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10950 = 8'h32 == r_count_53_io_out ? io_r_50_b : _GEN_10949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10951 = 8'h33 == r_count_53_io_out ? io_r_51_b : _GEN_10950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10952 = 8'h34 == r_count_53_io_out ? io_r_52_b : _GEN_10951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10953 = 8'h35 == r_count_53_io_out ? io_r_53_b : _GEN_10952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10954 = 8'h36 == r_count_53_io_out ? io_r_54_b : _GEN_10953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10955 = 8'h37 == r_count_53_io_out ? io_r_55_b : _GEN_10954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10956 = 8'h38 == r_count_53_io_out ? io_r_56_b : _GEN_10955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10957 = 8'h39 == r_count_53_io_out ? io_r_57_b : _GEN_10956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10958 = 8'h3a == r_count_53_io_out ? io_r_58_b : _GEN_10957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10959 = 8'h3b == r_count_53_io_out ? io_r_59_b : _GEN_10958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10960 = 8'h3c == r_count_53_io_out ? io_r_60_b : _GEN_10959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10961 = 8'h3d == r_count_53_io_out ? io_r_61_b : _GEN_10960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10962 = 8'h3e == r_count_53_io_out ? io_r_62_b : _GEN_10961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10963 = 8'h3f == r_count_53_io_out ? io_r_63_b : _GEN_10962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10964 = 8'h40 == r_count_53_io_out ? io_r_64_b : _GEN_10963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10965 = 8'h41 == r_count_53_io_out ? io_r_65_b : _GEN_10964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10966 = 8'h42 == r_count_53_io_out ? io_r_66_b : _GEN_10965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10967 = 8'h43 == r_count_53_io_out ? io_r_67_b : _GEN_10966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10968 = 8'h44 == r_count_53_io_out ? io_r_68_b : _GEN_10967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10969 = 8'h45 == r_count_53_io_out ? io_r_69_b : _GEN_10968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10970 = 8'h46 == r_count_53_io_out ? io_r_70_b : _GEN_10969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10971 = 8'h47 == r_count_53_io_out ? io_r_71_b : _GEN_10970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10972 = 8'h48 == r_count_53_io_out ? io_r_72_b : _GEN_10971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10973 = 8'h49 == r_count_53_io_out ? io_r_73_b : _GEN_10972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10974 = 8'h4a == r_count_53_io_out ? io_r_74_b : _GEN_10973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10975 = 8'h4b == r_count_53_io_out ? io_r_75_b : _GEN_10974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10976 = 8'h4c == r_count_53_io_out ? io_r_76_b : _GEN_10975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10977 = 8'h4d == r_count_53_io_out ? io_r_77_b : _GEN_10976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10978 = 8'h4e == r_count_53_io_out ? io_r_78_b : _GEN_10977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10979 = 8'h4f == r_count_53_io_out ? io_r_79_b : _GEN_10978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10980 = 8'h50 == r_count_53_io_out ? io_r_80_b : _GEN_10979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10981 = 8'h51 == r_count_53_io_out ? io_r_81_b : _GEN_10980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10982 = 8'h52 == r_count_53_io_out ? io_r_82_b : _GEN_10981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10983 = 8'h53 == r_count_53_io_out ? io_r_83_b : _GEN_10982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10984 = 8'h54 == r_count_53_io_out ? io_r_84_b : _GEN_10983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10985 = 8'h55 == r_count_53_io_out ? io_r_85_b : _GEN_10984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10986 = 8'h56 == r_count_53_io_out ? io_r_86_b : _GEN_10985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10987 = 8'h57 == r_count_53_io_out ? io_r_87_b : _GEN_10986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10988 = 8'h58 == r_count_53_io_out ? io_r_88_b : _GEN_10987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10989 = 8'h59 == r_count_53_io_out ? io_r_89_b : _GEN_10988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10990 = 8'h5a == r_count_53_io_out ? io_r_90_b : _GEN_10989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10991 = 8'h5b == r_count_53_io_out ? io_r_91_b : _GEN_10990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10992 = 8'h5c == r_count_53_io_out ? io_r_92_b : _GEN_10991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10993 = 8'h5d == r_count_53_io_out ? io_r_93_b : _GEN_10992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10994 = 8'h5e == r_count_53_io_out ? io_r_94_b : _GEN_10993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10995 = 8'h5f == r_count_53_io_out ? io_r_95_b : _GEN_10994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10996 = 8'h60 == r_count_53_io_out ? io_r_96_b : _GEN_10995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10997 = 8'h61 == r_count_53_io_out ? io_r_97_b : _GEN_10996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10998 = 8'h62 == r_count_53_io_out ? io_r_98_b : _GEN_10997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_10999 = 8'h63 == r_count_53_io_out ? io_r_99_b : _GEN_10998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11000 = 8'h64 == r_count_53_io_out ? io_r_100_b : _GEN_10999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11001 = 8'h65 == r_count_53_io_out ? io_r_101_b : _GEN_11000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11002 = 8'h66 == r_count_53_io_out ? io_r_102_b : _GEN_11001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11003 = 8'h67 == r_count_53_io_out ? io_r_103_b : _GEN_11002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11004 = 8'h68 == r_count_53_io_out ? io_r_104_b : _GEN_11003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11005 = 8'h69 == r_count_53_io_out ? io_r_105_b : _GEN_11004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11006 = 8'h6a == r_count_53_io_out ? io_r_106_b : _GEN_11005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11007 = 8'h6b == r_count_53_io_out ? io_r_107_b : _GEN_11006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11008 = 8'h6c == r_count_53_io_out ? io_r_108_b : _GEN_11007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11009 = 8'h6d == r_count_53_io_out ? io_r_109_b : _GEN_11008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11010 = 8'h6e == r_count_53_io_out ? io_r_110_b : _GEN_11009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11011 = 8'h6f == r_count_53_io_out ? io_r_111_b : _GEN_11010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11012 = 8'h70 == r_count_53_io_out ? io_r_112_b : _GEN_11011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11013 = 8'h71 == r_count_53_io_out ? io_r_113_b : _GEN_11012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11014 = 8'h72 == r_count_53_io_out ? io_r_114_b : _GEN_11013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11015 = 8'h73 == r_count_53_io_out ? io_r_115_b : _GEN_11014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11016 = 8'h74 == r_count_53_io_out ? io_r_116_b : _GEN_11015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11017 = 8'h75 == r_count_53_io_out ? io_r_117_b : _GEN_11016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11018 = 8'h76 == r_count_53_io_out ? io_r_118_b : _GEN_11017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11019 = 8'h77 == r_count_53_io_out ? io_r_119_b : _GEN_11018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11020 = 8'h78 == r_count_53_io_out ? io_r_120_b : _GEN_11019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11021 = 8'h79 == r_count_53_io_out ? io_r_121_b : _GEN_11020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11022 = 8'h7a == r_count_53_io_out ? io_r_122_b : _GEN_11021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11023 = 8'h7b == r_count_53_io_out ? io_r_123_b : _GEN_11022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11024 = 8'h7c == r_count_53_io_out ? io_r_124_b : _GEN_11023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11025 = 8'h7d == r_count_53_io_out ? io_r_125_b : _GEN_11024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11026 = 8'h7e == r_count_53_io_out ? io_r_126_b : _GEN_11025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11027 = 8'h7f == r_count_53_io_out ? io_r_127_b : _GEN_11026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11028 = 8'h80 == r_count_53_io_out ? io_r_128_b : _GEN_11027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11029 = 8'h81 == r_count_53_io_out ? io_r_129_b : _GEN_11028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11030 = 8'h82 == r_count_53_io_out ? io_r_130_b : _GEN_11029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11031 = 8'h83 == r_count_53_io_out ? io_r_131_b : _GEN_11030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11032 = 8'h84 == r_count_53_io_out ? io_r_132_b : _GEN_11031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11033 = 8'h85 == r_count_53_io_out ? io_r_133_b : _GEN_11032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11034 = 8'h86 == r_count_53_io_out ? io_r_134_b : _GEN_11033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11035 = 8'h87 == r_count_53_io_out ? io_r_135_b : _GEN_11034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11036 = 8'h88 == r_count_53_io_out ? io_r_136_b : _GEN_11035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11037 = 8'h89 == r_count_53_io_out ? io_r_137_b : _GEN_11036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11038 = 8'h8a == r_count_53_io_out ? io_r_138_b : _GEN_11037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11039 = 8'h8b == r_count_53_io_out ? io_r_139_b : _GEN_11038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11040 = 8'h8c == r_count_53_io_out ? io_r_140_b : _GEN_11039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11041 = 8'h8d == r_count_53_io_out ? io_r_141_b : _GEN_11040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11042 = 8'h8e == r_count_53_io_out ? io_r_142_b : _GEN_11041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11043 = 8'h8f == r_count_53_io_out ? io_r_143_b : _GEN_11042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11044 = 8'h90 == r_count_53_io_out ? io_r_144_b : _GEN_11043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11045 = 8'h91 == r_count_53_io_out ? io_r_145_b : _GEN_11044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11046 = 8'h92 == r_count_53_io_out ? io_r_146_b : _GEN_11045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11047 = 8'h93 == r_count_53_io_out ? io_r_147_b : _GEN_11046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11048 = 8'h94 == r_count_53_io_out ? io_r_148_b : _GEN_11047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11049 = 8'h95 == r_count_53_io_out ? io_r_149_b : _GEN_11048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11050 = 8'h96 == r_count_53_io_out ? io_r_150_b : _GEN_11049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11051 = 8'h97 == r_count_53_io_out ? io_r_151_b : _GEN_11050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11052 = 8'h98 == r_count_53_io_out ? io_r_152_b : _GEN_11051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11053 = 8'h99 == r_count_53_io_out ? io_r_153_b : _GEN_11052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11054 = 8'h9a == r_count_53_io_out ? io_r_154_b : _GEN_11053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11055 = 8'h9b == r_count_53_io_out ? io_r_155_b : _GEN_11054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11056 = 8'h9c == r_count_53_io_out ? io_r_156_b : _GEN_11055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11057 = 8'h9d == r_count_53_io_out ? io_r_157_b : _GEN_11056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11058 = 8'h9e == r_count_53_io_out ? io_r_158_b : _GEN_11057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11059 = 8'h9f == r_count_53_io_out ? io_r_159_b : _GEN_11058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11060 = 8'ha0 == r_count_53_io_out ? io_r_160_b : _GEN_11059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11061 = 8'ha1 == r_count_53_io_out ? io_r_161_b : _GEN_11060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11062 = 8'ha2 == r_count_53_io_out ? io_r_162_b : _GEN_11061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11063 = 8'ha3 == r_count_53_io_out ? io_r_163_b : _GEN_11062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11064 = 8'ha4 == r_count_53_io_out ? io_r_164_b : _GEN_11063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11065 = 8'ha5 == r_count_53_io_out ? io_r_165_b : _GEN_11064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11066 = 8'ha6 == r_count_53_io_out ? io_r_166_b : _GEN_11065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11067 = 8'ha7 == r_count_53_io_out ? io_r_167_b : _GEN_11066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11068 = 8'ha8 == r_count_53_io_out ? io_r_168_b : _GEN_11067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11069 = 8'ha9 == r_count_53_io_out ? io_r_169_b : _GEN_11068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11070 = 8'haa == r_count_53_io_out ? io_r_170_b : _GEN_11069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11071 = 8'hab == r_count_53_io_out ? io_r_171_b : _GEN_11070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11072 = 8'hac == r_count_53_io_out ? io_r_172_b : _GEN_11071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11073 = 8'had == r_count_53_io_out ? io_r_173_b : _GEN_11072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11074 = 8'hae == r_count_53_io_out ? io_r_174_b : _GEN_11073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11075 = 8'haf == r_count_53_io_out ? io_r_175_b : _GEN_11074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11076 = 8'hb0 == r_count_53_io_out ? io_r_176_b : _GEN_11075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11077 = 8'hb1 == r_count_53_io_out ? io_r_177_b : _GEN_11076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11078 = 8'hb2 == r_count_53_io_out ? io_r_178_b : _GEN_11077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11079 = 8'hb3 == r_count_53_io_out ? io_r_179_b : _GEN_11078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11080 = 8'hb4 == r_count_53_io_out ? io_r_180_b : _GEN_11079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11081 = 8'hb5 == r_count_53_io_out ? io_r_181_b : _GEN_11080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11082 = 8'hb6 == r_count_53_io_out ? io_r_182_b : _GEN_11081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11083 = 8'hb7 == r_count_53_io_out ? io_r_183_b : _GEN_11082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11084 = 8'hb8 == r_count_53_io_out ? io_r_184_b : _GEN_11083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11085 = 8'hb9 == r_count_53_io_out ? io_r_185_b : _GEN_11084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11086 = 8'hba == r_count_53_io_out ? io_r_186_b : _GEN_11085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11087 = 8'hbb == r_count_53_io_out ? io_r_187_b : _GEN_11086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11088 = 8'hbc == r_count_53_io_out ? io_r_188_b : _GEN_11087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11089 = 8'hbd == r_count_53_io_out ? io_r_189_b : _GEN_11088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11090 = 8'hbe == r_count_53_io_out ? io_r_190_b : _GEN_11089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11091 = 8'hbf == r_count_53_io_out ? io_r_191_b : _GEN_11090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11092 = 8'hc0 == r_count_53_io_out ? io_r_192_b : _GEN_11091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11093 = 8'hc1 == r_count_53_io_out ? io_r_193_b : _GEN_11092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11094 = 8'hc2 == r_count_53_io_out ? io_r_194_b : _GEN_11093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11095 = 8'hc3 == r_count_53_io_out ? io_r_195_b : _GEN_11094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11096 = 8'hc4 == r_count_53_io_out ? io_r_196_b : _GEN_11095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11097 = 8'hc5 == r_count_53_io_out ? io_r_197_b : _GEN_11096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11098 = 8'hc6 == r_count_53_io_out ? io_r_198_b : _GEN_11097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11101 = 8'h1 == r_count_54_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11102 = 8'h2 == r_count_54_io_out ? io_r_2_b : _GEN_11101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11103 = 8'h3 == r_count_54_io_out ? io_r_3_b : _GEN_11102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11104 = 8'h4 == r_count_54_io_out ? io_r_4_b : _GEN_11103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11105 = 8'h5 == r_count_54_io_out ? io_r_5_b : _GEN_11104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11106 = 8'h6 == r_count_54_io_out ? io_r_6_b : _GEN_11105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11107 = 8'h7 == r_count_54_io_out ? io_r_7_b : _GEN_11106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11108 = 8'h8 == r_count_54_io_out ? io_r_8_b : _GEN_11107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11109 = 8'h9 == r_count_54_io_out ? io_r_9_b : _GEN_11108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11110 = 8'ha == r_count_54_io_out ? io_r_10_b : _GEN_11109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11111 = 8'hb == r_count_54_io_out ? io_r_11_b : _GEN_11110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11112 = 8'hc == r_count_54_io_out ? io_r_12_b : _GEN_11111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11113 = 8'hd == r_count_54_io_out ? io_r_13_b : _GEN_11112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11114 = 8'he == r_count_54_io_out ? io_r_14_b : _GEN_11113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11115 = 8'hf == r_count_54_io_out ? io_r_15_b : _GEN_11114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11116 = 8'h10 == r_count_54_io_out ? io_r_16_b : _GEN_11115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11117 = 8'h11 == r_count_54_io_out ? io_r_17_b : _GEN_11116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11118 = 8'h12 == r_count_54_io_out ? io_r_18_b : _GEN_11117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11119 = 8'h13 == r_count_54_io_out ? io_r_19_b : _GEN_11118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11120 = 8'h14 == r_count_54_io_out ? io_r_20_b : _GEN_11119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11121 = 8'h15 == r_count_54_io_out ? io_r_21_b : _GEN_11120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11122 = 8'h16 == r_count_54_io_out ? io_r_22_b : _GEN_11121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11123 = 8'h17 == r_count_54_io_out ? io_r_23_b : _GEN_11122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11124 = 8'h18 == r_count_54_io_out ? io_r_24_b : _GEN_11123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11125 = 8'h19 == r_count_54_io_out ? io_r_25_b : _GEN_11124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11126 = 8'h1a == r_count_54_io_out ? io_r_26_b : _GEN_11125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11127 = 8'h1b == r_count_54_io_out ? io_r_27_b : _GEN_11126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11128 = 8'h1c == r_count_54_io_out ? io_r_28_b : _GEN_11127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11129 = 8'h1d == r_count_54_io_out ? io_r_29_b : _GEN_11128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11130 = 8'h1e == r_count_54_io_out ? io_r_30_b : _GEN_11129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11131 = 8'h1f == r_count_54_io_out ? io_r_31_b : _GEN_11130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11132 = 8'h20 == r_count_54_io_out ? io_r_32_b : _GEN_11131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11133 = 8'h21 == r_count_54_io_out ? io_r_33_b : _GEN_11132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11134 = 8'h22 == r_count_54_io_out ? io_r_34_b : _GEN_11133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11135 = 8'h23 == r_count_54_io_out ? io_r_35_b : _GEN_11134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11136 = 8'h24 == r_count_54_io_out ? io_r_36_b : _GEN_11135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11137 = 8'h25 == r_count_54_io_out ? io_r_37_b : _GEN_11136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11138 = 8'h26 == r_count_54_io_out ? io_r_38_b : _GEN_11137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11139 = 8'h27 == r_count_54_io_out ? io_r_39_b : _GEN_11138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11140 = 8'h28 == r_count_54_io_out ? io_r_40_b : _GEN_11139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11141 = 8'h29 == r_count_54_io_out ? io_r_41_b : _GEN_11140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11142 = 8'h2a == r_count_54_io_out ? io_r_42_b : _GEN_11141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11143 = 8'h2b == r_count_54_io_out ? io_r_43_b : _GEN_11142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11144 = 8'h2c == r_count_54_io_out ? io_r_44_b : _GEN_11143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11145 = 8'h2d == r_count_54_io_out ? io_r_45_b : _GEN_11144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11146 = 8'h2e == r_count_54_io_out ? io_r_46_b : _GEN_11145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11147 = 8'h2f == r_count_54_io_out ? io_r_47_b : _GEN_11146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11148 = 8'h30 == r_count_54_io_out ? io_r_48_b : _GEN_11147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11149 = 8'h31 == r_count_54_io_out ? io_r_49_b : _GEN_11148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11150 = 8'h32 == r_count_54_io_out ? io_r_50_b : _GEN_11149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11151 = 8'h33 == r_count_54_io_out ? io_r_51_b : _GEN_11150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11152 = 8'h34 == r_count_54_io_out ? io_r_52_b : _GEN_11151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11153 = 8'h35 == r_count_54_io_out ? io_r_53_b : _GEN_11152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11154 = 8'h36 == r_count_54_io_out ? io_r_54_b : _GEN_11153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11155 = 8'h37 == r_count_54_io_out ? io_r_55_b : _GEN_11154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11156 = 8'h38 == r_count_54_io_out ? io_r_56_b : _GEN_11155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11157 = 8'h39 == r_count_54_io_out ? io_r_57_b : _GEN_11156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11158 = 8'h3a == r_count_54_io_out ? io_r_58_b : _GEN_11157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11159 = 8'h3b == r_count_54_io_out ? io_r_59_b : _GEN_11158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11160 = 8'h3c == r_count_54_io_out ? io_r_60_b : _GEN_11159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11161 = 8'h3d == r_count_54_io_out ? io_r_61_b : _GEN_11160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11162 = 8'h3e == r_count_54_io_out ? io_r_62_b : _GEN_11161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11163 = 8'h3f == r_count_54_io_out ? io_r_63_b : _GEN_11162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11164 = 8'h40 == r_count_54_io_out ? io_r_64_b : _GEN_11163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11165 = 8'h41 == r_count_54_io_out ? io_r_65_b : _GEN_11164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11166 = 8'h42 == r_count_54_io_out ? io_r_66_b : _GEN_11165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11167 = 8'h43 == r_count_54_io_out ? io_r_67_b : _GEN_11166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11168 = 8'h44 == r_count_54_io_out ? io_r_68_b : _GEN_11167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11169 = 8'h45 == r_count_54_io_out ? io_r_69_b : _GEN_11168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11170 = 8'h46 == r_count_54_io_out ? io_r_70_b : _GEN_11169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11171 = 8'h47 == r_count_54_io_out ? io_r_71_b : _GEN_11170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11172 = 8'h48 == r_count_54_io_out ? io_r_72_b : _GEN_11171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11173 = 8'h49 == r_count_54_io_out ? io_r_73_b : _GEN_11172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11174 = 8'h4a == r_count_54_io_out ? io_r_74_b : _GEN_11173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11175 = 8'h4b == r_count_54_io_out ? io_r_75_b : _GEN_11174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11176 = 8'h4c == r_count_54_io_out ? io_r_76_b : _GEN_11175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11177 = 8'h4d == r_count_54_io_out ? io_r_77_b : _GEN_11176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11178 = 8'h4e == r_count_54_io_out ? io_r_78_b : _GEN_11177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11179 = 8'h4f == r_count_54_io_out ? io_r_79_b : _GEN_11178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11180 = 8'h50 == r_count_54_io_out ? io_r_80_b : _GEN_11179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11181 = 8'h51 == r_count_54_io_out ? io_r_81_b : _GEN_11180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11182 = 8'h52 == r_count_54_io_out ? io_r_82_b : _GEN_11181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11183 = 8'h53 == r_count_54_io_out ? io_r_83_b : _GEN_11182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11184 = 8'h54 == r_count_54_io_out ? io_r_84_b : _GEN_11183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11185 = 8'h55 == r_count_54_io_out ? io_r_85_b : _GEN_11184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11186 = 8'h56 == r_count_54_io_out ? io_r_86_b : _GEN_11185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11187 = 8'h57 == r_count_54_io_out ? io_r_87_b : _GEN_11186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11188 = 8'h58 == r_count_54_io_out ? io_r_88_b : _GEN_11187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11189 = 8'h59 == r_count_54_io_out ? io_r_89_b : _GEN_11188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11190 = 8'h5a == r_count_54_io_out ? io_r_90_b : _GEN_11189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11191 = 8'h5b == r_count_54_io_out ? io_r_91_b : _GEN_11190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11192 = 8'h5c == r_count_54_io_out ? io_r_92_b : _GEN_11191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11193 = 8'h5d == r_count_54_io_out ? io_r_93_b : _GEN_11192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11194 = 8'h5e == r_count_54_io_out ? io_r_94_b : _GEN_11193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11195 = 8'h5f == r_count_54_io_out ? io_r_95_b : _GEN_11194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11196 = 8'h60 == r_count_54_io_out ? io_r_96_b : _GEN_11195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11197 = 8'h61 == r_count_54_io_out ? io_r_97_b : _GEN_11196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11198 = 8'h62 == r_count_54_io_out ? io_r_98_b : _GEN_11197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11199 = 8'h63 == r_count_54_io_out ? io_r_99_b : _GEN_11198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11200 = 8'h64 == r_count_54_io_out ? io_r_100_b : _GEN_11199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11201 = 8'h65 == r_count_54_io_out ? io_r_101_b : _GEN_11200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11202 = 8'h66 == r_count_54_io_out ? io_r_102_b : _GEN_11201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11203 = 8'h67 == r_count_54_io_out ? io_r_103_b : _GEN_11202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11204 = 8'h68 == r_count_54_io_out ? io_r_104_b : _GEN_11203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11205 = 8'h69 == r_count_54_io_out ? io_r_105_b : _GEN_11204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11206 = 8'h6a == r_count_54_io_out ? io_r_106_b : _GEN_11205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11207 = 8'h6b == r_count_54_io_out ? io_r_107_b : _GEN_11206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11208 = 8'h6c == r_count_54_io_out ? io_r_108_b : _GEN_11207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11209 = 8'h6d == r_count_54_io_out ? io_r_109_b : _GEN_11208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11210 = 8'h6e == r_count_54_io_out ? io_r_110_b : _GEN_11209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11211 = 8'h6f == r_count_54_io_out ? io_r_111_b : _GEN_11210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11212 = 8'h70 == r_count_54_io_out ? io_r_112_b : _GEN_11211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11213 = 8'h71 == r_count_54_io_out ? io_r_113_b : _GEN_11212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11214 = 8'h72 == r_count_54_io_out ? io_r_114_b : _GEN_11213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11215 = 8'h73 == r_count_54_io_out ? io_r_115_b : _GEN_11214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11216 = 8'h74 == r_count_54_io_out ? io_r_116_b : _GEN_11215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11217 = 8'h75 == r_count_54_io_out ? io_r_117_b : _GEN_11216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11218 = 8'h76 == r_count_54_io_out ? io_r_118_b : _GEN_11217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11219 = 8'h77 == r_count_54_io_out ? io_r_119_b : _GEN_11218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11220 = 8'h78 == r_count_54_io_out ? io_r_120_b : _GEN_11219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11221 = 8'h79 == r_count_54_io_out ? io_r_121_b : _GEN_11220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11222 = 8'h7a == r_count_54_io_out ? io_r_122_b : _GEN_11221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11223 = 8'h7b == r_count_54_io_out ? io_r_123_b : _GEN_11222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11224 = 8'h7c == r_count_54_io_out ? io_r_124_b : _GEN_11223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11225 = 8'h7d == r_count_54_io_out ? io_r_125_b : _GEN_11224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11226 = 8'h7e == r_count_54_io_out ? io_r_126_b : _GEN_11225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11227 = 8'h7f == r_count_54_io_out ? io_r_127_b : _GEN_11226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11228 = 8'h80 == r_count_54_io_out ? io_r_128_b : _GEN_11227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11229 = 8'h81 == r_count_54_io_out ? io_r_129_b : _GEN_11228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11230 = 8'h82 == r_count_54_io_out ? io_r_130_b : _GEN_11229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11231 = 8'h83 == r_count_54_io_out ? io_r_131_b : _GEN_11230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11232 = 8'h84 == r_count_54_io_out ? io_r_132_b : _GEN_11231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11233 = 8'h85 == r_count_54_io_out ? io_r_133_b : _GEN_11232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11234 = 8'h86 == r_count_54_io_out ? io_r_134_b : _GEN_11233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11235 = 8'h87 == r_count_54_io_out ? io_r_135_b : _GEN_11234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11236 = 8'h88 == r_count_54_io_out ? io_r_136_b : _GEN_11235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11237 = 8'h89 == r_count_54_io_out ? io_r_137_b : _GEN_11236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11238 = 8'h8a == r_count_54_io_out ? io_r_138_b : _GEN_11237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11239 = 8'h8b == r_count_54_io_out ? io_r_139_b : _GEN_11238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11240 = 8'h8c == r_count_54_io_out ? io_r_140_b : _GEN_11239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11241 = 8'h8d == r_count_54_io_out ? io_r_141_b : _GEN_11240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11242 = 8'h8e == r_count_54_io_out ? io_r_142_b : _GEN_11241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11243 = 8'h8f == r_count_54_io_out ? io_r_143_b : _GEN_11242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11244 = 8'h90 == r_count_54_io_out ? io_r_144_b : _GEN_11243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11245 = 8'h91 == r_count_54_io_out ? io_r_145_b : _GEN_11244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11246 = 8'h92 == r_count_54_io_out ? io_r_146_b : _GEN_11245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11247 = 8'h93 == r_count_54_io_out ? io_r_147_b : _GEN_11246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11248 = 8'h94 == r_count_54_io_out ? io_r_148_b : _GEN_11247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11249 = 8'h95 == r_count_54_io_out ? io_r_149_b : _GEN_11248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11250 = 8'h96 == r_count_54_io_out ? io_r_150_b : _GEN_11249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11251 = 8'h97 == r_count_54_io_out ? io_r_151_b : _GEN_11250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11252 = 8'h98 == r_count_54_io_out ? io_r_152_b : _GEN_11251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11253 = 8'h99 == r_count_54_io_out ? io_r_153_b : _GEN_11252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11254 = 8'h9a == r_count_54_io_out ? io_r_154_b : _GEN_11253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11255 = 8'h9b == r_count_54_io_out ? io_r_155_b : _GEN_11254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11256 = 8'h9c == r_count_54_io_out ? io_r_156_b : _GEN_11255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11257 = 8'h9d == r_count_54_io_out ? io_r_157_b : _GEN_11256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11258 = 8'h9e == r_count_54_io_out ? io_r_158_b : _GEN_11257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11259 = 8'h9f == r_count_54_io_out ? io_r_159_b : _GEN_11258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11260 = 8'ha0 == r_count_54_io_out ? io_r_160_b : _GEN_11259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11261 = 8'ha1 == r_count_54_io_out ? io_r_161_b : _GEN_11260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11262 = 8'ha2 == r_count_54_io_out ? io_r_162_b : _GEN_11261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11263 = 8'ha3 == r_count_54_io_out ? io_r_163_b : _GEN_11262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11264 = 8'ha4 == r_count_54_io_out ? io_r_164_b : _GEN_11263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11265 = 8'ha5 == r_count_54_io_out ? io_r_165_b : _GEN_11264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11266 = 8'ha6 == r_count_54_io_out ? io_r_166_b : _GEN_11265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11267 = 8'ha7 == r_count_54_io_out ? io_r_167_b : _GEN_11266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11268 = 8'ha8 == r_count_54_io_out ? io_r_168_b : _GEN_11267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11269 = 8'ha9 == r_count_54_io_out ? io_r_169_b : _GEN_11268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11270 = 8'haa == r_count_54_io_out ? io_r_170_b : _GEN_11269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11271 = 8'hab == r_count_54_io_out ? io_r_171_b : _GEN_11270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11272 = 8'hac == r_count_54_io_out ? io_r_172_b : _GEN_11271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11273 = 8'had == r_count_54_io_out ? io_r_173_b : _GEN_11272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11274 = 8'hae == r_count_54_io_out ? io_r_174_b : _GEN_11273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11275 = 8'haf == r_count_54_io_out ? io_r_175_b : _GEN_11274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11276 = 8'hb0 == r_count_54_io_out ? io_r_176_b : _GEN_11275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11277 = 8'hb1 == r_count_54_io_out ? io_r_177_b : _GEN_11276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11278 = 8'hb2 == r_count_54_io_out ? io_r_178_b : _GEN_11277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11279 = 8'hb3 == r_count_54_io_out ? io_r_179_b : _GEN_11278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11280 = 8'hb4 == r_count_54_io_out ? io_r_180_b : _GEN_11279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11281 = 8'hb5 == r_count_54_io_out ? io_r_181_b : _GEN_11280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11282 = 8'hb6 == r_count_54_io_out ? io_r_182_b : _GEN_11281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11283 = 8'hb7 == r_count_54_io_out ? io_r_183_b : _GEN_11282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11284 = 8'hb8 == r_count_54_io_out ? io_r_184_b : _GEN_11283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11285 = 8'hb9 == r_count_54_io_out ? io_r_185_b : _GEN_11284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11286 = 8'hba == r_count_54_io_out ? io_r_186_b : _GEN_11285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11287 = 8'hbb == r_count_54_io_out ? io_r_187_b : _GEN_11286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11288 = 8'hbc == r_count_54_io_out ? io_r_188_b : _GEN_11287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11289 = 8'hbd == r_count_54_io_out ? io_r_189_b : _GEN_11288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11290 = 8'hbe == r_count_54_io_out ? io_r_190_b : _GEN_11289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11291 = 8'hbf == r_count_54_io_out ? io_r_191_b : _GEN_11290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11292 = 8'hc0 == r_count_54_io_out ? io_r_192_b : _GEN_11291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11293 = 8'hc1 == r_count_54_io_out ? io_r_193_b : _GEN_11292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11294 = 8'hc2 == r_count_54_io_out ? io_r_194_b : _GEN_11293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11295 = 8'hc3 == r_count_54_io_out ? io_r_195_b : _GEN_11294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11296 = 8'hc4 == r_count_54_io_out ? io_r_196_b : _GEN_11295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11297 = 8'hc5 == r_count_54_io_out ? io_r_197_b : _GEN_11296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11298 = 8'hc6 == r_count_54_io_out ? io_r_198_b : _GEN_11297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11301 = 8'h1 == r_count_55_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11302 = 8'h2 == r_count_55_io_out ? io_r_2_b : _GEN_11301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11303 = 8'h3 == r_count_55_io_out ? io_r_3_b : _GEN_11302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11304 = 8'h4 == r_count_55_io_out ? io_r_4_b : _GEN_11303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11305 = 8'h5 == r_count_55_io_out ? io_r_5_b : _GEN_11304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11306 = 8'h6 == r_count_55_io_out ? io_r_6_b : _GEN_11305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11307 = 8'h7 == r_count_55_io_out ? io_r_7_b : _GEN_11306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11308 = 8'h8 == r_count_55_io_out ? io_r_8_b : _GEN_11307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11309 = 8'h9 == r_count_55_io_out ? io_r_9_b : _GEN_11308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11310 = 8'ha == r_count_55_io_out ? io_r_10_b : _GEN_11309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11311 = 8'hb == r_count_55_io_out ? io_r_11_b : _GEN_11310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11312 = 8'hc == r_count_55_io_out ? io_r_12_b : _GEN_11311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11313 = 8'hd == r_count_55_io_out ? io_r_13_b : _GEN_11312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11314 = 8'he == r_count_55_io_out ? io_r_14_b : _GEN_11313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11315 = 8'hf == r_count_55_io_out ? io_r_15_b : _GEN_11314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11316 = 8'h10 == r_count_55_io_out ? io_r_16_b : _GEN_11315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11317 = 8'h11 == r_count_55_io_out ? io_r_17_b : _GEN_11316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11318 = 8'h12 == r_count_55_io_out ? io_r_18_b : _GEN_11317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11319 = 8'h13 == r_count_55_io_out ? io_r_19_b : _GEN_11318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11320 = 8'h14 == r_count_55_io_out ? io_r_20_b : _GEN_11319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11321 = 8'h15 == r_count_55_io_out ? io_r_21_b : _GEN_11320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11322 = 8'h16 == r_count_55_io_out ? io_r_22_b : _GEN_11321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11323 = 8'h17 == r_count_55_io_out ? io_r_23_b : _GEN_11322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11324 = 8'h18 == r_count_55_io_out ? io_r_24_b : _GEN_11323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11325 = 8'h19 == r_count_55_io_out ? io_r_25_b : _GEN_11324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11326 = 8'h1a == r_count_55_io_out ? io_r_26_b : _GEN_11325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11327 = 8'h1b == r_count_55_io_out ? io_r_27_b : _GEN_11326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11328 = 8'h1c == r_count_55_io_out ? io_r_28_b : _GEN_11327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11329 = 8'h1d == r_count_55_io_out ? io_r_29_b : _GEN_11328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11330 = 8'h1e == r_count_55_io_out ? io_r_30_b : _GEN_11329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11331 = 8'h1f == r_count_55_io_out ? io_r_31_b : _GEN_11330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11332 = 8'h20 == r_count_55_io_out ? io_r_32_b : _GEN_11331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11333 = 8'h21 == r_count_55_io_out ? io_r_33_b : _GEN_11332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11334 = 8'h22 == r_count_55_io_out ? io_r_34_b : _GEN_11333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11335 = 8'h23 == r_count_55_io_out ? io_r_35_b : _GEN_11334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11336 = 8'h24 == r_count_55_io_out ? io_r_36_b : _GEN_11335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11337 = 8'h25 == r_count_55_io_out ? io_r_37_b : _GEN_11336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11338 = 8'h26 == r_count_55_io_out ? io_r_38_b : _GEN_11337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11339 = 8'h27 == r_count_55_io_out ? io_r_39_b : _GEN_11338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11340 = 8'h28 == r_count_55_io_out ? io_r_40_b : _GEN_11339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11341 = 8'h29 == r_count_55_io_out ? io_r_41_b : _GEN_11340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11342 = 8'h2a == r_count_55_io_out ? io_r_42_b : _GEN_11341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11343 = 8'h2b == r_count_55_io_out ? io_r_43_b : _GEN_11342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11344 = 8'h2c == r_count_55_io_out ? io_r_44_b : _GEN_11343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11345 = 8'h2d == r_count_55_io_out ? io_r_45_b : _GEN_11344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11346 = 8'h2e == r_count_55_io_out ? io_r_46_b : _GEN_11345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11347 = 8'h2f == r_count_55_io_out ? io_r_47_b : _GEN_11346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11348 = 8'h30 == r_count_55_io_out ? io_r_48_b : _GEN_11347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11349 = 8'h31 == r_count_55_io_out ? io_r_49_b : _GEN_11348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11350 = 8'h32 == r_count_55_io_out ? io_r_50_b : _GEN_11349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11351 = 8'h33 == r_count_55_io_out ? io_r_51_b : _GEN_11350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11352 = 8'h34 == r_count_55_io_out ? io_r_52_b : _GEN_11351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11353 = 8'h35 == r_count_55_io_out ? io_r_53_b : _GEN_11352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11354 = 8'h36 == r_count_55_io_out ? io_r_54_b : _GEN_11353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11355 = 8'h37 == r_count_55_io_out ? io_r_55_b : _GEN_11354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11356 = 8'h38 == r_count_55_io_out ? io_r_56_b : _GEN_11355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11357 = 8'h39 == r_count_55_io_out ? io_r_57_b : _GEN_11356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11358 = 8'h3a == r_count_55_io_out ? io_r_58_b : _GEN_11357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11359 = 8'h3b == r_count_55_io_out ? io_r_59_b : _GEN_11358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11360 = 8'h3c == r_count_55_io_out ? io_r_60_b : _GEN_11359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11361 = 8'h3d == r_count_55_io_out ? io_r_61_b : _GEN_11360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11362 = 8'h3e == r_count_55_io_out ? io_r_62_b : _GEN_11361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11363 = 8'h3f == r_count_55_io_out ? io_r_63_b : _GEN_11362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11364 = 8'h40 == r_count_55_io_out ? io_r_64_b : _GEN_11363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11365 = 8'h41 == r_count_55_io_out ? io_r_65_b : _GEN_11364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11366 = 8'h42 == r_count_55_io_out ? io_r_66_b : _GEN_11365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11367 = 8'h43 == r_count_55_io_out ? io_r_67_b : _GEN_11366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11368 = 8'h44 == r_count_55_io_out ? io_r_68_b : _GEN_11367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11369 = 8'h45 == r_count_55_io_out ? io_r_69_b : _GEN_11368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11370 = 8'h46 == r_count_55_io_out ? io_r_70_b : _GEN_11369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11371 = 8'h47 == r_count_55_io_out ? io_r_71_b : _GEN_11370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11372 = 8'h48 == r_count_55_io_out ? io_r_72_b : _GEN_11371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11373 = 8'h49 == r_count_55_io_out ? io_r_73_b : _GEN_11372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11374 = 8'h4a == r_count_55_io_out ? io_r_74_b : _GEN_11373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11375 = 8'h4b == r_count_55_io_out ? io_r_75_b : _GEN_11374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11376 = 8'h4c == r_count_55_io_out ? io_r_76_b : _GEN_11375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11377 = 8'h4d == r_count_55_io_out ? io_r_77_b : _GEN_11376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11378 = 8'h4e == r_count_55_io_out ? io_r_78_b : _GEN_11377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11379 = 8'h4f == r_count_55_io_out ? io_r_79_b : _GEN_11378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11380 = 8'h50 == r_count_55_io_out ? io_r_80_b : _GEN_11379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11381 = 8'h51 == r_count_55_io_out ? io_r_81_b : _GEN_11380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11382 = 8'h52 == r_count_55_io_out ? io_r_82_b : _GEN_11381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11383 = 8'h53 == r_count_55_io_out ? io_r_83_b : _GEN_11382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11384 = 8'h54 == r_count_55_io_out ? io_r_84_b : _GEN_11383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11385 = 8'h55 == r_count_55_io_out ? io_r_85_b : _GEN_11384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11386 = 8'h56 == r_count_55_io_out ? io_r_86_b : _GEN_11385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11387 = 8'h57 == r_count_55_io_out ? io_r_87_b : _GEN_11386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11388 = 8'h58 == r_count_55_io_out ? io_r_88_b : _GEN_11387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11389 = 8'h59 == r_count_55_io_out ? io_r_89_b : _GEN_11388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11390 = 8'h5a == r_count_55_io_out ? io_r_90_b : _GEN_11389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11391 = 8'h5b == r_count_55_io_out ? io_r_91_b : _GEN_11390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11392 = 8'h5c == r_count_55_io_out ? io_r_92_b : _GEN_11391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11393 = 8'h5d == r_count_55_io_out ? io_r_93_b : _GEN_11392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11394 = 8'h5e == r_count_55_io_out ? io_r_94_b : _GEN_11393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11395 = 8'h5f == r_count_55_io_out ? io_r_95_b : _GEN_11394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11396 = 8'h60 == r_count_55_io_out ? io_r_96_b : _GEN_11395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11397 = 8'h61 == r_count_55_io_out ? io_r_97_b : _GEN_11396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11398 = 8'h62 == r_count_55_io_out ? io_r_98_b : _GEN_11397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11399 = 8'h63 == r_count_55_io_out ? io_r_99_b : _GEN_11398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11400 = 8'h64 == r_count_55_io_out ? io_r_100_b : _GEN_11399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11401 = 8'h65 == r_count_55_io_out ? io_r_101_b : _GEN_11400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11402 = 8'h66 == r_count_55_io_out ? io_r_102_b : _GEN_11401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11403 = 8'h67 == r_count_55_io_out ? io_r_103_b : _GEN_11402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11404 = 8'h68 == r_count_55_io_out ? io_r_104_b : _GEN_11403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11405 = 8'h69 == r_count_55_io_out ? io_r_105_b : _GEN_11404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11406 = 8'h6a == r_count_55_io_out ? io_r_106_b : _GEN_11405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11407 = 8'h6b == r_count_55_io_out ? io_r_107_b : _GEN_11406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11408 = 8'h6c == r_count_55_io_out ? io_r_108_b : _GEN_11407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11409 = 8'h6d == r_count_55_io_out ? io_r_109_b : _GEN_11408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11410 = 8'h6e == r_count_55_io_out ? io_r_110_b : _GEN_11409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11411 = 8'h6f == r_count_55_io_out ? io_r_111_b : _GEN_11410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11412 = 8'h70 == r_count_55_io_out ? io_r_112_b : _GEN_11411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11413 = 8'h71 == r_count_55_io_out ? io_r_113_b : _GEN_11412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11414 = 8'h72 == r_count_55_io_out ? io_r_114_b : _GEN_11413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11415 = 8'h73 == r_count_55_io_out ? io_r_115_b : _GEN_11414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11416 = 8'h74 == r_count_55_io_out ? io_r_116_b : _GEN_11415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11417 = 8'h75 == r_count_55_io_out ? io_r_117_b : _GEN_11416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11418 = 8'h76 == r_count_55_io_out ? io_r_118_b : _GEN_11417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11419 = 8'h77 == r_count_55_io_out ? io_r_119_b : _GEN_11418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11420 = 8'h78 == r_count_55_io_out ? io_r_120_b : _GEN_11419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11421 = 8'h79 == r_count_55_io_out ? io_r_121_b : _GEN_11420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11422 = 8'h7a == r_count_55_io_out ? io_r_122_b : _GEN_11421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11423 = 8'h7b == r_count_55_io_out ? io_r_123_b : _GEN_11422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11424 = 8'h7c == r_count_55_io_out ? io_r_124_b : _GEN_11423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11425 = 8'h7d == r_count_55_io_out ? io_r_125_b : _GEN_11424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11426 = 8'h7e == r_count_55_io_out ? io_r_126_b : _GEN_11425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11427 = 8'h7f == r_count_55_io_out ? io_r_127_b : _GEN_11426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11428 = 8'h80 == r_count_55_io_out ? io_r_128_b : _GEN_11427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11429 = 8'h81 == r_count_55_io_out ? io_r_129_b : _GEN_11428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11430 = 8'h82 == r_count_55_io_out ? io_r_130_b : _GEN_11429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11431 = 8'h83 == r_count_55_io_out ? io_r_131_b : _GEN_11430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11432 = 8'h84 == r_count_55_io_out ? io_r_132_b : _GEN_11431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11433 = 8'h85 == r_count_55_io_out ? io_r_133_b : _GEN_11432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11434 = 8'h86 == r_count_55_io_out ? io_r_134_b : _GEN_11433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11435 = 8'h87 == r_count_55_io_out ? io_r_135_b : _GEN_11434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11436 = 8'h88 == r_count_55_io_out ? io_r_136_b : _GEN_11435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11437 = 8'h89 == r_count_55_io_out ? io_r_137_b : _GEN_11436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11438 = 8'h8a == r_count_55_io_out ? io_r_138_b : _GEN_11437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11439 = 8'h8b == r_count_55_io_out ? io_r_139_b : _GEN_11438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11440 = 8'h8c == r_count_55_io_out ? io_r_140_b : _GEN_11439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11441 = 8'h8d == r_count_55_io_out ? io_r_141_b : _GEN_11440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11442 = 8'h8e == r_count_55_io_out ? io_r_142_b : _GEN_11441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11443 = 8'h8f == r_count_55_io_out ? io_r_143_b : _GEN_11442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11444 = 8'h90 == r_count_55_io_out ? io_r_144_b : _GEN_11443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11445 = 8'h91 == r_count_55_io_out ? io_r_145_b : _GEN_11444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11446 = 8'h92 == r_count_55_io_out ? io_r_146_b : _GEN_11445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11447 = 8'h93 == r_count_55_io_out ? io_r_147_b : _GEN_11446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11448 = 8'h94 == r_count_55_io_out ? io_r_148_b : _GEN_11447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11449 = 8'h95 == r_count_55_io_out ? io_r_149_b : _GEN_11448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11450 = 8'h96 == r_count_55_io_out ? io_r_150_b : _GEN_11449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11451 = 8'h97 == r_count_55_io_out ? io_r_151_b : _GEN_11450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11452 = 8'h98 == r_count_55_io_out ? io_r_152_b : _GEN_11451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11453 = 8'h99 == r_count_55_io_out ? io_r_153_b : _GEN_11452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11454 = 8'h9a == r_count_55_io_out ? io_r_154_b : _GEN_11453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11455 = 8'h9b == r_count_55_io_out ? io_r_155_b : _GEN_11454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11456 = 8'h9c == r_count_55_io_out ? io_r_156_b : _GEN_11455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11457 = 8'h9d == r_count_55_io_out ? io_r_157_b : _GEN_11456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11458 = 8'h9e == r_count_55_io_out ? io_r_158_b : _GEN_11457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11459 = 8'h9f == r_count_55_io_out ? io_r_159_b : _GEN_11458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11460 = 8'ha0 == r_count_55_io_out ? io_r_160_b : _GEN_11459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11461 = 8'ha1 == r_count_55_io_out ? io_r_161_b : _GEN_11460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11462 = 8'ha2 == r_count_55_io_out ? io_r_162_b : _GEN_11461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11463 = 8'ha3 == r_count_55_io_out ? io_r_163_b : _GEN_11462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11464 = 8'ha4 == r_count_55_io_out ? io_r_164_b : _GEN_11463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11465 = 8'ha5 == r_count_55_io_out ? io_r_165_b : _GEN_11464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11466 = 8'ha6 == r_count_55_io_out ? io_r_166_b : _GEN_11465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11467 = 8'ha7 == r_count_55_io_out ? io_r_167_b : _GEN_11466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11468 = 8'ha8 == r_count_55_io_out ? io_r_168_b : _GEN_11467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11469 = 8'ha9 == r_count_55_io_out ? io_r_169_b : _GEN_11468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11470 = 8'haa == r_count_55_io_out ? io_r_170_b : _GEN_11469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11471 = 8'hab == r_count_55_io_out ? io_r_171_b : _GEN_11470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11472 = 8'hac == r_count_55_io_out ? io_r_172_b : _GEN_11471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11473 = 8'had == r_count_55_io_out ? io_r_173_b : _GEN_11472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11474 = 8'hae == r_count_55_io_out ? io_r_174_b : _GEN_11473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11475 = 8'haf == r_count_55_io_out ? io_r_175_b : _GEN_11474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11476 = 8'hb0 == r_count_55_io_out ? io_r_176_b : _GEN_11475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11477 = 8'hb1 == r_count_55_io_out ? io_r_177_b : _GEN_11476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11478 = 8'hb2 == r_count_55_io_out ? io_r_178_b : _GEN_11477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11479 = 8'hb3 == r_count_55_io_out ? io_r_179_b : _GEN_11478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11480 = 8'hb4 == r_count_55_io_out ? io_r_180_b : _GEN_11479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11481 = 8'hb5 == r_count_55_io_out ? io_r_181_b : _GEN_11480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11482 = 8'hb6 == r_count_55_io_out ? io_r_182_b : _GEN_11481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11483 = 8'hb7 == r_count_55_io_out ? io_r_183_b : _GEN_11482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11484 = 8'hb8 == r_count_55_io_out ? io_r_184_b : _GEN_11483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11485 = 8'hb9 == r_count_55_io_out ? io_r_185_b : _GEN_11484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11486 = 8'hba == r_count_55_io_out ? io_r_186_b : _GEN_11485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11487 = 8'hbb == r_count_55_io_out ? io_r_187_b : _GEN_11486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11488 = 8'hbc == r_count_55_io_out ? io_r_188_b : _GEN_11487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11489 = 8'hbd == r_count_55_io_out ? io_r_189_b : _GEN_11488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11490 = 8'hbe == r_count_55_io_out ? io_r_190_b : _GEN_11489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11491 = 8'hbf == r_count_55_io_out ? io_r_191_b : _GEN_11490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11492 = 8'hc0 == r_count_55_io_out ? io_r_192_b : _GEN_11491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11493 = 8'hc1 == r_count_55_io_out ? io_r_193_b : _GEN_11492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11494 = 8'hc2 == r_count_55_io_out ? io_r_194_b : _GEN_11493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11495 = 8'hc3 == r_count_55_io_out ? io_r_195_b : _GEN_11494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11496 = 8'hc4 == r_count_55_io_out ? io_r_196_b : _GEN_11495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11497 = 8'hc5 == r_count_55_io_out ? io_r_197_b : _GEN_11496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11498 = 8'hc6 == r_count_55_io_out ? io_r_198_b : _GEN_11497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11501 = 8'h1 == r_count_56_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11502 = 8'h2 == r_count_56_io_out ? io_r_2_b : _GEN_11501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11503 = 8'h3 == r_count_56_io_out ? io_r_3_b : _GEN_11502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11504 = 8'h4 == r_count_56_io_out ? io_r_4_b : _GEN_11503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11505 = 8'h5 == r_count_56_io_out ? io_r_5_b : _GEN_11504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11506 = 8'h6 == r_count_56_io_out ? io_r_6_b : _GEN_11505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11507 = 8'h7 == r_count_56_io_out ? io_r_7_b : _GEN_11506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11508 = 8'h8 == r_count_56_io_out ? io_r_8_b : _GEN_11507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11509 = 8'h9 == r_count_56_io_out ? io_r_9_b : _GEN_11508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11510 = 8'ha == r_count_56_io_out ? io_r_10_b : _GEN_11509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11511 = 8'hb == r_count_56_io_out ? io_r_11_b : _GEN_11510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11512 = 8'hc == r_count_56_io_out ? io_r_12_b : _GEN_11511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11513 = 8'hd == r_count_56_io_out ? io_r_13_b : _GEN_11512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11514 = 8'he == r_count_56_io_out ? io_r_14_b : _GEN_11513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11515 = 8'hf == r_count_56_io_out ? io_r_15_b : _GEN_11514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11516 = 8'h10 == r_count_56_io_out ? io_r_16_b : _GEN_11515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11517 = 8'h11 == r_count_56_io_out ? io_r_17_b : _GEN_11516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11518 = 8'h12 == r_count_56_io_out ? io_r_18_b : _GEN_11517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11519 = 8'h13 == r_count_56_io_out ? io_r_19_b : _GEN_11518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11520 = 8'h14 == r_count_56_io_out ? io_r_20_b : _GEN_11519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11521 = 8'h15 == r_count_56_io_out ? io_r_21_b : _GEN_11520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11522 = 8'h16 == r_count_56_io_out ? io_r_22_b : _GEN_11521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11523 = 8'h17 == r_count_56_io_out ? io_r_23_b : _GEN_11522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11524 = 8'h18 == r_count_56_io_out ? io_r_24_b : _GEN_11523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11525 = 8'h19 == r_count_56_io_out ? io_r_25_b : _GEN_11524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11526 = 8'h1a == r_count_56_io_out ? io_r_26_b : _GEN_11525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11527 = 8'h1b == r_count_56_io_out ? io_r_27_b : _GEN_11526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11528 = 8'h1c == r_count_56_io_out ? io_r_28_b : _GEN_11527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11529 = 8'h1d == r_count_56_io_out ? io_r_29_b : _GEN_11528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11530 = 8'h1e == r_count_56_io_out ? io_r_30_b : _GEN_11529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11531 = 8'h1f == r_count_56_io_out ? io_r_31_b : _GEN_11530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11532 = 8'h20 == r_count_56_io_out ? io_r_32_b : _GEN_11531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11533 = 8'h21 == r_count_56_io_out ? io_r_33_b : _GEN_11532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11534 = 8'h22 == r_count_56_io_out ? io_r_34_b : _GEN_11533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11535 = 8'h23 == r_count_56_io_out ? io_r_35_b : _GEN_11534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11536 = 8'h24 == r_count_56_io_out ? io_r_36_b : _GEN_11535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11537 = 8'h25 == r_count_56_io_out ? io_r_37_b : _GEN_11536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11538 = 8'h26 == r_count_56_io_out ? io_r_38_b : _GEN_11537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11539 = 8'h27 == r_count_56_io_out ? io_r_39_b : _GEN_11538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11540 = 8'h28 == r_count_56_io_out ? io_r_40_b : _GEN_11539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11541 = 8'h29 == r_count_56_io_out ? io_r_41_b : _GEN_11540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11542 = 8'h2a == r_count_56_io_out ? io_r_42_b : _GEN_11541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11543 = 8'h2b == r_count_56_io_out ? io_r_43_b : _GEN_11542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11544 = 8'h2c == r_count_56_io_out ? io_r_44_b : _GEN_11543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11545 = 8'h2d == r_count_56_io_out ? io_r_45_b : _GEN_11544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11546 = 8'h2e == r_count_56_io_out ? io_r_46_b : _GEN_11545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11547 = 8'h2f == r_count_56_io_out ? io_r_47_b : _GEN_11546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11548 = 8'h30 == r_count_56_io_out ? io_r_48_b : _GEN_11547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11549 = 8'h31 == r_count_56_io_out ? io_r_49_b : _GEN_11548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11550 = 8'h32 == r_count_56_io_out ? io_r_50_b : _GEN_11549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11551 = 8'h33 == r_count_56_io_out ? io_r_51_b : _GEN_11550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11552 = 8'h34 == r_count_56_io_out ? io_r_52_b : _GEN_11551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11553 = 8'h35 == r_count_56_io_out ? io_r_53_b : _GEN_11552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11554 = 8'h36 == r_count_56_io_out ? io_r_54_b : _GEN_11553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11555 = 8'h37 == r_count_56_io_out ? io_r_55_b : _GEN_11554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11556 = 8'h38 == r_count_56_io_out ? io_r_56_b : _GEN_11555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11557 = 8'h39 == r_count_56_io_out ? io_r_57_b : _GEN_11556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11558 = 8'h3a == r_count_56_io_out ? io_r_58_b : _GEN_11557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11559 = 8'h3b == r_count_56_io_out ? io_r_59_b : _GEN_11558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11560 = 8'h3c == r_count_56_io_out ? io_r_60_b : _GEN_11559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11561 = 8'h3d == r_count_56_io_out ? io_r_61_b : _GEN_11560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11562 = 8'h3e == r_count_56_io_out ? io_r_62_b : _GEN_11561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11563 = 8'h3f == r_count_56_io_out ? io_r_63_b : _GEN_11562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11564 = 8'h40 == r_count_56_io_out ? io_r_64_b : _GEN_11563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11565 = 8'h41 == r_count_56_io_out ? io_r_65_b : _GEN_11564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11566 = 8'h42 == r_count_56_io_out ? io_r_66_b : _GEN_11565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11567 = 8'h43 == r_count_56_io_out ? io_r_67_b : _GEN_11566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11568 = 8'h44 == r_count_56_io_out ? io_r_68_b : _GEN_11567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11569 = 8'h45 == r_count_56_io_out ? io_r_69_b : _GEN_11568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11570 = 8'h46 == r_count_56_io_out ? io_r_70_b : _GEN_11569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11571 = 8'h47 == r_count_56_io_out ? io_r_71_b : _GEN_11570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11572 = 8'h48 == r_count_56_io_out ? io_r_72_b : _GEN_11571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11573 = 8'h49 == r_count_56_io_out ? io_r_73_b : _GEN_11572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11574 = 8'h4a == r_count_56_io_out ? io_r_74_b : _GEN_11573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11575 = 8'h4b == r_count_56_io_out ? io_r_75_b : _GEN_11574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11576 = 8'h4c == r_count_56_io_out ? io_r_76_b : _GEN_11575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11577 = 8'h4d == r_count_56_io_out ? io_r_77_b : _GEN_11576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11578 = 8'h4e == r_count_56_io_out ? io_r_78_b : _GEN_11577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11579 = 8'h4f == r_count_56_io_out ? io_r_79_b : _GEN_11578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11580 = 8'h50 == r_count_56_io_out ? io_r_80_b : _GEN_11579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11581 = 8'h51 == r_count_56_io_out ? io_r_81_b : _GEN_11580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11582 = 8'h52 == r_count_56_io_out ? io_r_82_b : _GEN_11581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11583 = 8'h53 == r_count_56_io_out ? io_r_83_b : _GEN_11582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11584 = 8'h54 == r_count_56_io_out ? io_r_84_b : _GEN_11583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11585 = 8'h55 == r_count_56_io_out ? io_r_85_b : _GEN_11584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11586 = 8'h56 == r_count_56_io_out ? io_r_86_b : _GEN_11585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11587 = 8'h57 == r_count_56_io_out ? io_r_87_b : _GEN_11586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11588 = 8'h58 == r_count_56_io_out ? io_r_88_b : _GEN_11587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11589 = 8'h59 == r_count_56_io_out ? io_r_89_b : _GEN_11588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11590 = 8'h5a == r_count_56_io_out ? io_r_90_b : _GEN_11589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11591 = 8'h5b == r_count_56_io_out ? io_r_91_b : _GEN_11590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11592 = 8'h5c == r_count_56_io_out ? io_r_92_b : _GEN_11591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11593 = 8'h5d == r_count_56_io_out ? io_r_93_b : _GEN_11592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11594 = 8'h5e == r_count_56_io_out ? io_r_94_b : _GEN_11593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11595 = 8'h5f == r_count_56_io_out ? io_r_95_b : _GEN_11594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11596 = 8'h60 == r_count_56_io_out ? io_r_96_b : _GEN_11595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11597 = 8'h61 == r_count_56_io_out ? io_r_97_b : _GEN_11596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11598 = 8'h62 == r_count_56_io_out ? io_r_98_b : _GEN_11597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11599 = 8'h63 == r_count_56_io_out ? io_r_99_b : _GEN_11598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11600 = 8'h64 == r_count_56_io_out ? io_r_100_b : _GEN_11599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11601 = 8'h65 == r_count_56_io_out ? io_r_101_b : _GEN_11600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11602 = 8'h66 == r_count_56_io_out ? io_r_102_b : _GEN_11601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11603 = 8'h67 == r_count_56_io_out ? io_r_103_b : _GEN_11602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11604 = 8'h68 == r_count_56_io_out ? io_r_104_b : _GEN_11603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11605 = 8'h69 == r_count_56_io_out ? io_r_105_b : _GEN_11604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11606 = 8'h6a == r_count_56_io_out ? io_r_106_b : _GEN_11605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11607 = 8'h6b == r_count_56_io_out ? io_r_107_b : _GEN_11606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11608 = 8'h6c == r_count_56_io_out ? io_r_108_b : _GEN_11607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11609 = 8'h6d == r_count_56_io_out ? io_r_109_b : _GEN_11608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11610 = 8'h6e == r_count_56_io_out ? io_r_110_b : _GEN_11609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11611 = 8'h6f == r_count_56_io_out ? io_r_111_b : _GEN_11610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11612 = 8'h70 == r_count_56_io_out ? io_r_112_b : _GEN_11611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11613 = 8'h71 == r_count_56_io_out ? io_r_113_b : _GEN_11612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11614 = 8'h72 == r_count_56_io_out ? io_r_114_b : _GEN_11613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11615 = 8'h73 == r_count_56_io_out ? io_r_115_b : _GEN_11614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11616 = 8'h74 == r_count_56_io_out ? io_r_116_b : _GEN_11615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11617 = 8'h75 == r_count_56_io_out ? io_r_117_b : _GEN_11616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11618 = 8'h76 == r_count_56_io_out ? io_r_118_b : _GEN_11617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11619 = 8'h77 == r_count_56_io_out ? io_r_119_b : _GEN_11618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11620 = 8'h78 == r_count_56_io_out ? io_r_120_b : _GEN_11619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11621 = 8'h79 == r_count_56_io_out ? io_r_121_b : _GEN_11620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11622 = 8'h7a == r_count_56_io_out ? io_r_122_b : _GEN_11621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11623 = 8'h7b == r_count_56_io_out ? io_r_123_b : _GEN_11622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11624 = 8'h7c == r_count_56_io_out ? io_r_124_b : _GEN_11623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11625 = 8'h7d == r_count_56_io_out ? io_r_125_b : _GEN_11624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11626 = 8'h7e == r_count_56_io_out ? io_r_126_b : _GEN_11625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11627 = 8'h7f == r_count_56_io_out ? io_r_127_b : _GEN_11626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11628 = 8'h80 == r_count_56_io_out ? io_r_128_b : _GEN_11627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11629 = 8'h81 == r_count_56_io_out ? io_r_129_b : _GEN_11628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11630 = 8'h82 == r_count_56_io_out ? io_r_130_b : _GEN_11629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11631 = 8'h83 == r_count_56_io_out ? io_r_131_b : _GEN_11630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11632 = 8'h84 == r_count_56_io_out ? io_r_132_b : _GEN_11631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11633 = 8'h85 == r_count_56_io_out ? io_r_133_b : _GEN_11632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11634 = 8'h86 == r_count_56_io_out ? io_r_134_b : _GEN_11633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11635 = 8'h87 == r_count_56_io_out ? io_r_135_b : _GEN_11634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11636 = 8'h88 == r_count_56_io_out ? io_r_136_b : _GEN_11635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11637 = 8'h89 == r_count_56_io_out ? io_r_137_b : _GEN_11636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11638 = 8'h8a == r_count_56_io_out ? io_r_138_b : _GEN_11637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11639 = 8'h8b == r_count_56_io_out ? io_r_139_b : _GEN_11638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11640 = 8'h8c == r_count_56_io_out ? io_r_140_b : _GEN_11639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11641 = 8'h8d == r_count_56_io_out ? io_r_141_b : _GEN_11640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11642 = 8'h8e == r_count_56_io_out ? io_r_142_b : _GEN_11641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11643 = 8'h8f == r_count_56_io_out ? io_r_143_b : _GEN_11642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11644 = 8'h90 == r_count_56_io_out ? io_r_144_b : _GEN_11643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11645 = 8'h91 == r_count_56_io_out ? io_r_145_b : _GEN_11644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11646 = 8'h92 == r_count_56_io_out ? io_r_146_b : _GEN_11645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11647 = 8'h93 == r_count_56_io_out ? io_r_147_b : _GEN_11646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11648 = 8'h94 == r_count_56_io_out ? io_r_148_b : _GEN_11647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11649 = 8'h95 == r_count_56_io_out ? io_r_149_b : _GEN_11648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11650 = 8'h96 == r_count_56_io_out ? io_r_150_b : _GEN_11649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11651 = 8'h97 == r_count_56_io_out ? io_r_151_b : _GEN_11650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11652 = 8'h98 == r_count_56_io_out ? io_r_152_b : _GEN_11651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11653 = 8'h99 == r_count_56_io_out ? io_r_153_b : _GEN_11652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11654 = 8'h9a == r_count_56_io_out ? io_r_154_b : _GEN_11653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11655 = 8'h9b == r_count_56_io_out ? io_r_155_b : _GEN_11654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11656 = 8'h9c == r_count_56_io_out ? io_r_156_b : _GEN_11655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11657 = 8'h9d == r_count_56_io_out ? io_r_157_b : _GEN_11656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11658 = 8'h9e == r_count_56_io_out ? io_r_158_b : _GEN_11657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11659 = 8'h9f == r_count_56_io_out ? io_r_159_b : _GEN_11658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11660 = 8'ha0 == r_count_56_io_out ? io_r_160_b : _GEN_11659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11661 = 8'ha1 == r_count_56_io_out ? io_r_161_b : _GEN_11660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11662 = 8'ha2 == r_count_56_io_out ? io_r_162_b : _GEN_11661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11663 = 8'ha3 == r_count_56_io_out ? io_r_163_b : _GEN_11662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11664 = 8'ha4 == r_count_56_io_out ? io_r_164_b : _GEN_11663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11665 = 8'ha5 == r_count_56_io_out ? io_r_165_b : _GEN_11664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11666 = 8'ha6 == r_count_56_io_out ? io_r_166_b : _GEN_11665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11667 = 8'ha7 == r_count_56_io_out ? io_r_167_b : _GEN_11666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11668 = 8'ha8 == r_count_56_io_out ? io_r_168_b : _GEN_11667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11669 = 8'ha9 == r_count_56_io_out ? io_r_169_b : _GEN_11668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11670 = 8'haa == r_count_56_io_out ? io_r_170_b : _GEN_11669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11671 = 8'hab == r_count_56_io_out ? io_r_171_b : _GEN_11670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11672 = 8'hac == r_count_56_io_out ? io_r_172_b : _GEN_11671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11673 = 8'had == r_count_56_io_out ? io_r_173_b : _GEN_11672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11674 = 8'hae == r_count_56_io_out ? io_r_174_b : _GEN_11673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11675 = 8'haf == r_count_56_io_out ? io_r_175_b : _GEN_11674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11676 = 8'hb0 == r_count_56_io_out ? io_r_176_b : _GEN_11675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11677 = 8'hb1 == r_count_56_io_out ? io_r_177_b : _GEN_11676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11678 = 8'hb2 == r_count_56_io_out ? io_r_178_b : _GEN_11677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11679 = 8'hb3 == r_count_56_io_out ? io_r_179_b : _GEN_11678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11680 = 8'hb4 == r_count_56_io_out ? io_r_180_b : _GEN_11679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11681 = 8'hb5 == r_count_56_io_out ? io_r_181_b : _GEN_11680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11682 = 8'hb6 == r_count_56_io_out ? io_r_182_b : _GEN_11681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11683 = 8'hb7 == r_count_56_io_out ? io_r_183_b : _GEN_11682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11684 = 8'hb8 == r_count_56_io_out ? io_r_184_b : _GEN_11683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11685 = 8'hb9 == r_count_56_io_out ? io_r_185_b : _GEN_11684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11686 = 8'hba == r_count_56_io_out ? io_r_186_b : _GEN_11685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11687 = 8'hbb == r_count_56_io_out ? io_r_187_b : _GEN_11686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11688 = 8'hbc == r_count_56_io_out ? io_r_188_b : _GEN_11687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11689 = 8'hbd == r_count_56_io_out ? io_r_189_b : _GEN_11688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11690 = 8'hbe == r_count_56_io_out ? io_r_190_b : _GEN_11689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11691 = 8'hbf == r_count_56_io_out ? io_r_191_b : _GEN_11690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11692 = 8'hc0 == r_count_56_io_out ? io_r_192_b : _GEN_11691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11693 = 8'hc1 == r_count_56_io_out ? io_r_193_b : _GEN_11692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11694 = 8'hc2 == r_count_56_io_out ? io_r_194_b : _GEN_11693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11695 = 8'hc3 == r_count_56_io_out ? io_r_195_b : _GEN_11694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11696 = 8'hc4 == r_count_56_io_out ? io_r_196_b : _GEN_11695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11697 = 8'hc5 == r_count_56_io_out ? io_r_197_b : _GEN_11696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11698 = 8'hc6 == r_count_56_io_out ? io_r_198_b : _GEN_11697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11701 = 8'h1 == r_count_57_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11702 = 8'h2 == r_count_57_io_out ? io_r_2_b : _GEN_11701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11703 = 8'h3 == r_count_57_io_out ? io_r_3_b : _GEN_11702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11704 = 8'h4 == r_count_57_io_out ? io_r_4_b : _GEN_11703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11705 = 8'h5 == r_count_57_io_out ? io_r_5_b : _GEN_11704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11706 = 8'h6 == r_count_57_io_out ? io_r_6_b : _GEN_11705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11707 = 8'h7 == r_count_57_io_out ? io_r_7_b : _GEN_11706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11708 = 8'h8 == r_count_57_io_out ? io_r_8_b : _GEN_11707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11709 = 8'h9 == r_count_57_io_out ? io_r_9_b : _GEN_11708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11710 = 8'ha == r_count_57_io_out ? io_r_10_b : _GEN_11709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11711 = 8'hb == r_count_57_io_out ? io_r_11_b : _GEN_11710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11712 = 8'hc == r_count_57_io_out ? io_r_12_b : _GEN_11711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11713 = 8'hd == r_count_57_io_out ? io_r_13_b : _GEN_11712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11714 = 8'he == r_count_57_io_out ? io_r_14_b : _GEN_11713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11715 = 8'hf == r_count_57_io_out ? io_r_15_b : _GEN_11714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11716 = 8'h10 == r_count_57_io_out ? io_r_16_b : _GEN_11715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11717 = 8'h11 == r_count_57_io_out ? io_r_17_b : _GEN_11716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11718 = 8'h12 == r_count_57_io_out ? io_r_18_b : _GEN_11717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11719 = 8'h13 == r_count_57_io_out ? io_r_19_b : _GEN_11718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11720 = 8'h14 == r_count_57_io_out ? io_r_20_b : _GEN_11719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11721 = 8'h15 == r_count_57_io_out ? io_r_21_b : _GEN_11720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11722 = 8'h16 == r_count_57_io_out ? io_r_22_b : _GEN_11721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11723 = 8'h17 == r_count_57_io_out ? io_r_23_b : _GEN_11722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11724 = 8'h18 == r_count_57_io_out ? io_r_24_b : _GEN_11723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11725 = 8'h19 == r_count_57_io_out ? io_r_25_b : _GEN_11724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11726 = 8'h1a == r_count_57_io_out ? io_r_26_b : _GEN_11725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11727 = 8'h1b == r_count_57_io_out ? io_r_27_b : _GEN_11726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11728 = 8'h1c == r_count_57_io_out ? io_r_28_b : _GEN_11727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11729 = 8'h1d == r_count_57_io_out ? io_r_29_b : _GEN_11728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11730 = 8'h1e == r_count_57_io_out ? io_r_30_b : _GEN_11729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11731 = 8'h1f == r_count_57_io_out ? io_r_31_b : _GEN_11730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11732 = 8'h20 == r_count_57_io_out ? io_r_32_b : _GEN_11731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11733 = 8'h21 == r_count_57_io_out ? io_r_33_b : _GEN_11732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11734 = 8'h22 == r_count_57_io_out ? io_r_34_b : _GEN_11733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11735 = 8'h23 == r_count_57_io_out ? io_r_35_b : _GEN_11734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11736 = 8'h24 == r_count_57_io_out ? io_r_36_b : _GEN_11735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11737 = 8'h25 == r_count_57_io_out ? io_r_37_b : _GEN_11736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11738 = 8'h26 == r_count_57_io_out ? io_r_38_b : _GEN_11737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11739 = 8'h27 == r_count_57_io_out ? io_r_39_b : _GEN_11738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11740 = 8'h28 == r_count_57_io_out ? io_r_40_b : _GEN_11739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11741 = 8'h29 == r_count_57_io_out ? io_r_41_b : _GEN_11740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11742 = 8'h2a == r_count_57_io_out ? io_r_42_b : _GEN_11741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11743 = 8'h2b == r_count_57_io_out ? io_r_43_b : _GEN_11742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11744 = 8'h2c == r_count_57_io_out ? io_r_44_b : _GEN_11743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11745 = 8'h2d == r_count_57_io_out ? io_r_45_b : _GEN_11744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11746 = 8'h2e == r_count_57_io_out ? io_r_46_b : _GEN_11745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11747 = 8'h2f == r_count_57_io_out ? io_r_47_b : _GEN_11746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11748 = 8'h30 == r_count_57_io_out ? io_r_48_b : _GEN_11747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11749 = 8'h31 == r_count_57_io_out ? io_r_49_b : _GEN_11748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11750 = 8'h32 == r_count_57_io_out ? io_r_50_b : _GEN_11749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11751 = 8'h33 == r_count_57_io_out ? io_r_51_b : _GEN_11750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11752 = 8'h34 == r_count_57_io_out ? io_r_52_b : _GEN_11751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11753 = 8'h35 == r_count_57_io_out ? io_r_53_b : _GEN_11752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11754 = 8'h36 == r_count_57_io_out ? io_r_54_b : _GEN_11753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11755 = 8'h37 == r_count_57_io_out ? io_r_55_b : _GEN_11754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11756 = 8'h38 == r_count_57_io_out ? io_r_56_b : _GEN_11755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11757 = 8'h39 == r_count_57_io_out ? io_r_57_b : _GEN_11756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11758 = 8'h3a == r_count_57_io_out ? io_r_58_b : _GEN_11757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11759 = 8'h3b == r_count_57_io_out ? io_r_59_b : _GEN_11758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11760 = 8'h3c == r_count_57_io_out ? io_r_60_b : _GEN_11759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11761 = 8'h3d == r_count_57_io_out ? io_r_61_b : _GEN_11760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11762 = 8'h3e == r_count_57_io_out ? io_r_62_b : _GEN_11761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11763 = 8'h3f == r_count_57_io_out ? io_r_63_b : _GEN_11762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11764 = 8'h40 == r_count_57_io_out ? io_r_64_b : _GEN_11763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11765 = 8'h41 == r_count_57_io_out ? io_r_65_b : _GEN_11764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11766 = 8'h42 == r_count_57_io_out ? io_r_66_b : _GEN_11765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11767 = 8'h43 == r_count_57_io_out ? io_r_67_b : _GEN_11766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11768 = 8'h44 == r_count_57_io_out ? io_r_68_b : _GEN_11767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11769 = 8'h45 == r_count_57_io_out ? io_r_69_b : _GEN_11768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11770 = 8'h46 == r_count_57_io_out ? io_r_70_b : _GEN_11769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11771 = 8'h47 == r_count_57_io_out ? io_r_71_b : _GEN_11770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11772 = 8'h48 == r_count_57_io_out ? io_r_72_b : _GEN_11771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11773 = 8'h49 == r_count_57_io_out ? io_r_73_b : _GEN_11772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11774 = 8'h4a == r_count_57_io_out ? io_r_74_b : _GEN_11773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11775 = 8'h4b == r_count_57_io_out ? io_r_75_b : _GEN_11774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11776 = 8'h4c == r_count_57_io_out ? io_r_76_b : _GEN_11775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11777 = 8'h4d == r_count_57_io_out ? io_r_77_b : _GEN_11776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11778 = 8'h4e == r_count_57_io_out ? io_r_78_b : _GEN_11777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11779 = 8'h4f == r_count_57_io_out ? io_r_79_b : _GEN_11778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11780 = 8'h50 == r_count_57_io_out ? io_r_80_b : _GEN_11779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11781 = 8'h51 == r_count_57_io_out ? io_r_81_b : _GEN_11780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11782 = 8'h52 == r_count_57_io_out ? io_r_82_b : _GEN_11781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11783 = 8'h53 == r_count_57_io_out ? io_r_83_b : _GEN_11782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11784 = 8'h54 == r_count_57_io_out ? io_r_84_b : _GEN_11783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11785 = 8'h55 == r_count_57_io_out ? io_r_85_b : _GEN_11784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11786 = 8'h56 == r_count_57_io_out ? io_r_86_b : _GEN_11785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11787 = 8'h57 == r_count_57_io_out ? io_r_87_b : _GEN_11786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11788 = 8'h58 == r_count_57_io_out ? io_r_88_b : _GEN_11787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11789 = 8'h59 == r_count_57_io_out ? io_r_89_b : _GEN_11788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11790 = 8'h5a == r_count_57_io_out ? io_r_90_b : _GEN_11789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11791 = 8'h5b == r_count_57_io_out ? io_r_91_b : _GEN_11790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11792 = 8'h5c == r_count_57_io_out ? io_r_92_b : _GEN_11791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11793 = 8'h5d == r_count_57_io_out ? io_r_93_b : _GEN_11792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11794 = 8'h5e == r_count_57_io_out ? io_r_94_b : _GEN_11793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11795 = 8'h5f == r_count_57_io_out ? io_r_95_b : _GEN_11794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11796 = 8'h60 == r_count_57_io_out ? io_r_96_b : _GEN_11795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11797 = 8'h61 == r_count_57_io_out ? io_r_97_b : _GEN_11796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11798 = 8'h62 == r_count_57_io_out ? io_r_98_b : _GEN_11797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11799 = 8'h63 == r_count_57_io_out ? io_r_99_b : _GEN_11798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11800 = 8'h64 == r_count_57_io_out ? io_r_100_b : _GEN_11799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11801 = 8'h65 == r_count_57_io_out ? io_r_101_b : _GEN_11800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11802 = 8'h66 == r_count_57_io_out ? io_r_102_b : _GEN_11801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11803 = 8'h67 == r_count_57_io_out ? io_r_103_b : _GEN_11802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11804 = 8'h68 == r_count_57_io_out ? io_r_104_b : _GEN_11803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11805 = 8'h69 == r_count_57_io_out ? io_r_105_b : _GEN_11804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11806 = 8'h6a == r_count_57_io_out ? io_r_106_b : _GEN_11805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11807 = 8'h6b == r_count_57_io_out ? io_r_107_b : _GEN_11806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11808 = 8'h6c == r_count_57_io_out ? io_r_108_b : _GEN_11807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11809 = 8'h6d == r_count_57_io_out ? io_r_109_b : _GEN_11808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11810 = 8'h6e == r_count_57_io_out ? io_r_110_b : _GEN_11809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11811 = 8'h6f == r_count_57_io_out ? io_r_111_b : _GEN_11810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11812 = 8'h70 == r_count_57_io_out ? io_r_112_b : _GEN_11811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11813 = 8'h71 == r_count_57_io_out ? io_r_113_b : _GEN_11812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11814 = 8'h72 == r_count_57_io_out ? io_r_114_b : _GEN_11813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11815 = 8'h73 == r_count_57_io_out ? io_r_115_b : _GEN_11814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11816 = 8'h74 == r_count_57_io_out ? io_r_116_b : _GEN_11815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11817 = 8'h75 == r_count_57_io_out ? io_r_117_b : _GEN_11816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11818 = 8'h76 == r_count_57_io_out ? io_r_118_b : _GEN_11817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11819 = 8'h77 == r_count_57_io_out ? io_r_119_b : _GEN_11818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11820 = 8'h78 == r_count_57_io_out ? io_r_120_b : _GEN_11819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11821 = 8'h79 == r_count_57_io_out ? io_r_121_b : _GEN_11820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11822 = 8'h7a == r_count_57_io_out ? io_r_122_b : _GEN_11821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11823 = 8'h7b == r_count_57_io_out ? io_r_123_b : _GEN_11822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11824 = 8'h7c == r_count_57_io_out ? io_r_124_b : _GEN_11823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11825 = 8'h7d == r_count_57_io_out ? io_r_125_b : _GEN_11824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11826 = 8'h7e == r_count_57_io_out ? io_r_126_b : _GEN_11825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11827 = 8'h7f == r_count_57_io_out ? io_r_127_b : _GEN_11826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11828 = 8'h80 == r_count_57_io_out ? io_r_128_b : _GEN_11827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11829 = 8'h81 == r_count_57_io_out ? io_r_129_b : _GEN_11828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11830 = 8'h82 == r_count_57_io_out ? io_r_130_b : _GEN_11829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11831 = 8'h83 == r_count_57_io_out ? io_r_131_b : _GEN_11830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11832 = 8'h84 == r_count_57_io_out ? io_r_132_b : _GEN_11831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11833 = 8'h85 == r_count_57_io_out ? io_r_133_b : _GEN_11832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11834 = 8'h86 == r_count_57_io_out ? io_r_134_b : _GEN_11833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11835 = 8'h87 == r_count_57_io_out ? io_r_135_b : _GEN_11834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11836 = 8'h88 == r_count_57_io_out ? io_r_136_b : _GEN_11835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11837 = 8'h89 == r_count_57_io_out ? io_r_137_b : _GEN_11836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11838 = 8'h8a == r_count_57_io_out ? io_r_138_b : _GEN_11837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11839 = 8'h8b == r_count_57_io_out ? io_r_139_b : _GEN_11838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11840 = 8'h8c == r_count_57_io_out ? io_r_140_b : _GEN_11839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11841 = 8'h8d == r_count_57_io_out ? io_r_141_b : _GEN_11840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11842 = 8'h8e == r_count_57_io_out ? io_r_142_b : _GEN_11841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11843 = 8'h8f == r_count_57_io_out ? io_r_143_b : _GEN_11842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11844 = 8'h90 == r_count_57_io_out ? io_r_144_b : _GEN_11843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11845 = 8'h91 == r_count_57_io_out ? io_r_145_b : _GEN_11844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11846 = 8'h92 == r_count_57_io_out ? io_r_146_b : _GEN_11845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11847 = 8'h93 == r_count_57_io_out ? io_r_147_b : _GEN_11846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11848 = 8'h94 == r_count_57_io_out ? io_r_148_b : _GEN_11847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11849 = 8'h95 == r_count_57_io_out ? io_r_149_b : _GEN_11848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11850 = 8'h96 == r_count_57_io_out ? io_r_150_b : _GEN_11849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11851 = 8'h97 == r_count_57_io_out ? io_r_151_b : _GEN_11850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11852 = 8'h98 == r_count_57_io_out ? io_r_152_b : _GEN_11851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11853 = 8'h99 == r_count_57_io_out ? io_r_153_b : _GEN_11852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11854 = 8'h9a == r_count_57_io_out ? io_r_154_b : _GEN_11853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11855 = 8'h9b == r_count_57_io_out ? io_r_155_b : _GEN_11854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11856 = 8'h9c == r_count_57_io_out ? io_r_156_b : _GEN_11855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11857 = 8'h9d == r_count_57_io_out ? io_r_157_b : _GEN_11856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11858 = 8'h9e == r_count_57_io_out ? io_r_158_b : _GEN_11857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11859 = 8'h9f == r_count_57_io_out ? io_r_159_b : _GEN_11858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11860 = 8'ha0 == r_count_57_io_out ? io_r_160_b : _GEN_11859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11861 = 8'ha1 == r_count_57_io_out ? io_r_161_b : _GEN_11860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11862 = 8'ha2 == r_count_57_io_out ? io_r_162_b : _GEN_11861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11863 = 8'ha3 == r_count_57_io_out ? io_r_163_b : _GEN_11862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11864 = 8'ha4 == r_count_57_io_out ? io_r_164_b : _GEN_11863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11865 = 8'ha5 == r_count_57_io_out ? io_r_165_b : _GEN_11864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11866 = 8'ha6 == r_count_57_io_out ? io_r_166_b : _GEN_11865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11867 = 8'ha7 == r_count_57_io_out ? io_r_167_b : _GEN_11866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11868 = 8'ha8 == r_count_57_io_out ? io_r_168_b : _GEN_11867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11869 = 8'ha9 == r_count_57_io_out ? io_r_169_b : _GEN_11868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11870 = 8'haa == r_count_57_io_out ? io_r_170_b : _GEN_11869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11871 = 8'hab == r_count_57_io_out ? io_r_171_b : _GEN_11870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11872 = 8'hac == r_count_57_io_out ? io_r_172_b : _GEN_11871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11873 = 8'had == r_count_57_io_out ? io_r_173_b : _GEN_11872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11874 = 8'hae == r_count_57_io_out ? io_r_174_b : _GEN_11873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11875 = 8'haf == r_count_57_io_out ? io_r_175_b : _GEN_11874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11876 = 8'hb0 == r_count_57_io_out ? io_r_176_b : _GEN_11875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11877 = 8'hb1 == r_count_57_io_out ? io_r_177_b : _GEN_11876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11878 = 8'hb2 == r_count_57_io_out ? io_r_178_b : _GEN_11877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11879 = 8'hb3 == r_count_57_io_out ? io_r_179_b : _GEN_11878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11880 = 8'hb4 == r_count_57_io_out ? io_r_180_b : _GEN_11879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11881 = 8'hb5 == r_count_57_io_out ? io_r_181_b : _GEN_11880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11882 = 8'hb6 == r_count_57_io_out ? io_r_182_b : _GEN_11881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11883 = 8'hb7 == r_count_57_io_out ? io_r_183_b : _GEN_11882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11884 = 8'hb8 == r_count_57_io_out ? io_r_184_b : _GEN_11883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11885 = 8'hb9 == r_count_57_io_out ? io_r_185_b : _GEN_11884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11886 = 8'hba == r_count_57_io_out ? io_r_186_b : _GEN_11885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11887 = 8'hbb == r_count_57_io_out ? io_r_187_b : _GEN_11886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11888 = 8'hbc == r_count_57_io_out ? io_r_188_b : _GEN_11887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11889 = 8'hbd == r_count_57_io_out ? io_r_189_b : _GEN_11888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11890 = 8'hbe == r_count_57_io_out ? io_r_190_b : _GEN_11889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11891 = 8'hbf == r_count_57_io_out ? io_r_191_b : _GEN_11890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11892 = 8'hc0 == r_count_57_io_out ? io_r_192_b : _GEN_11891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11893 = 8'hc1 == r_count_57_io_out ? io_r_193_b : _GEN_11892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11894 = 8'hc2 == r_count_57_io_out ? io_r_194_b : _GEN_11893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11895 = 8'hc3 == r_count_57_io_out ? io_r_195_b : _GEN_11894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11896 = 8'hc4 == r_count_57_io_out ? io_r_196_b : _GEN_11895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11897 = 8'hc5 == r_count_57_io_out ? io_r_197_b : _GEN_11896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11898 = 8'hc6 == r_count_57_io_out ? io_r_198_b : _GEN_11897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11901 = 8'h1 == r_count_58_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11902 = 8'h2 == r_count_58_io_out ? io_r_2_b : _GEN_11901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11903 = 8'h3 == r_count_58_io_out ? io_r_3_b : _GEN_11902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11904 = 8'h4 == r_count_58_io_out ? io_r_4_b : _GEN_11903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11905 = 8'h5 == r_count_58_io_out ? io_r_5_b : _GEN_11904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11906 = 8'h6 == r_count_58_io_out ? io_r_6_b : _GEN_11905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11907 = 8'h7 == r_count_58_io_out ? io_r_7_b : _GEN_11906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11908 = 8'h8 == r_count_58_io_out ? io_r_8_b : _GEN_11907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11909 = 8'h9 == r_count_58_io_out ? io_r_9_b : _GEN_11908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11910 = 8'ha == r_count_58_io_out ? io_r_10_b : _GEN_11909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11911 = 8'hb == r_count_58_io_out ? io_r_11_b : _GEN_11910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11912 = 8'hc == r_count_58_io_out ? io_r_12_b : _GEN_11911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11913 = 8'hd == r_count_58_io_out ? io_r_13_b : _GEN_11912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11914 = 8'he == r_count_58_io_out ? io_r_14_b : _GEN_11913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11915 = 8'hf == r_count_58_io_out ? io_r_15_b : _GEN_11914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11916 = 8'h10 == r_count_58_io_out ? io_r_16_b : _GEN_11915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11917 = 8'h11 == r_count_58_io_out ? io_r_17_b : _GEN_11916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11918 = 8'h12 == r_count_58_io_out ? io_r_18_b : _GEN_11917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11919 = 8'h13 == r_count_58_io_out ? io_r_19_b : _GEN_11918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11920 = 8'h14 == r_count_58_io_out ? io_r_20_b : _GEN_11919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11921 = 8'h15 == r_count_58_io_out ? io_r_21_b : _GEN_11920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11922 = 8'h16 == r_count_58_io_out ? io_r_22_b : _GEN_11921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11923 = 8'h17 == r_count_58_io_out ? io_r_23_b : _GEN_11922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11924 = 8'h18 == r_count_58_io_out ? io_r_24_b : _GEN_11923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11925 = 8'h19 == r_count_58_io_out ? io_r_25_b : _GEN_11924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11926 = 8'h1a == r_count_58_io_out ? io_r_26_b : _GEN_11925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11927 = 8'h1b == r_count_58_io_out ? io_r_27_b : _GEN_11926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11928 = 8'h1c == r_count_58_io_out ? io_r_28_b : _GEN_11927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11929 = 8'h1d == r_count_58_io_out ? io_r_29_b : _GEN_11928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11930 = 8'h1e == r_count_58_io_out ? io_r_30_b : _GEN_11929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11931 = 8'h1f == r_count_58_io_out ? io_r_31_b : _GEN_11930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11932 = 8'h20 == r_count_58_io_out ? io_r_32_b : _GEN_11931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11933 = 8'h21 == r_count_58_io_out ? io_r_33_b : _GEN_11932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11934 = 8'h22 == r_count_58_io_out ? io_r_34_b : _GEN_11933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11935 = 8'h23 == r_count_58_io_out ? io_r_35_b : _GEN_11934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11936 = 8'h24 == r_count_58_io_out ? io_r_36_b : _GEN_11935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11937 = 8'h25 == r_count_58_io_out ? io_r_37_b : _GEN_11936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11938 = 8'h26 == r_count_58_io_out ? io_r_38_b : _GEN_11937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11939 = 8'h27 == r_count_58_io_out ? io_r_39_b : _GEN_11938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11940 = 8'h28 == r_count_58_io_out ? io_r_40_b : _GEN_11939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11941 = 8'h29 == r_count_58_io_out ? io_r_41_b : _GEN_11940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11942 = 8'h2a == r_count_58_io_out ? io_r_42_b : _GEN_11941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11943 = 8'h2b == r_count_58_io_out ? io_r_43_b : _GEN_11942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11944 = 8'h2c == r_count_58_io_out ? io_r_44_b : _GEN_11943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11945 = 8'h2d == r_count_58_io_out ? io_r_45_b : _GEN_11944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11946 = 8'h2e == r_count_58_io_out ? io_r_46_b : _GEN_11945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11947 = 8'h2f == r_count_58_io_out ? io_r_47_b : _GEN_11946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11948 = 8'h30 == r_count_58_io_out ? io_r_48_b : _GEN_11947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11949 = 8'h31 == r_count_58_io_out ? io_r_49_b : _GEN_11948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11950 = 8'h32 == r_count_58_io_out ? io_r_50_b : _GEN_11949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11951 = 8'h33 == r_count_58_io_out ? io_r_51_b : _GEN_11950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11952 = 8'h34 == r_count_58_io_out ? io_r_52_b : _GEN_11951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11953 = 8'h35 == r_count_58_io_out ? io_r_53_b : _GEN_11952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11954 = 8'h36 == r_count_58_io_out ? io_r_54_b : _GEN_11953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11955 = 8'h37 == r_count_58_io_out ? io_r_55_b : _GEN_11954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11956 = 8'h38 == r_count_58_io_out ? io_r_56_b : _GEN_11955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11957 = 8'h39 == r_count_58_io_out ? io_r_57_b : _GEN_11956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11958 = 8'h3a == r_count_58_io_out ? io_r_58_b : _GEN_11957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11959 = 8'h3b == r_count_58_io_out ? io_r_59_b : _GEN_11958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11960 = 8'h3c == r_count_58_io_out ? io_r_60_b : _GEN_11959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11961 = 8'h3d == r_count_58_io_out ? io_r_61_b : _GEN_11960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11962 = 8'h3e == r_count_58_io_out ? io_r_62_b : _GEN_11961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11963 = 8'h3f == r_count_58_io_out ? io_r_63_b : _GEN_11962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11964 = 8'h40 == r_count_58_io_out ? io_r_64_b : _GEN_11963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11965 = 8'h41 == r_count_58_io_out ? io_r_65_b : _GEN_11964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11966 = 8'h42 == r_count_58_io_out ? io_r_66_b : _GEN_11965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11967 = 8'h43 == r_count_58_io_out ? io_r_67_b : _GEN_11966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11968 = 8'h44 == r_count_58_io_out ? io_r_68_b : _GEN_11967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11969 = 8'h45 == r_count_58_io_out ? io_r_69_b : _GEN_11968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11970 = 8'h46 == r_count_58_io_out ? io_r_70_b : _GEN_11969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11971 = 8'h47 == r_count_58_io_out ? io_r_71_b : _GEN_11970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11972 = 8'h48 == r_count_58_io_out ? io_r_72_b : _GEN_11971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11973 = 8'h49 == r_count_58_io_out ? io_r_73_b : _GEN_11972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11974 = 8'h4a == r_count_58_io_out ? io_r_74_b : _GEN_11973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11975 = 8'h4b == r_count_58_io_out ? io_r_75_b : _GEN_11974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11976 = 8'h4c == r_count_58_io_out ? io_r_76_b : _GEN_11975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11977 = 8'h4d == r_count_58_io_out ? io_r_77_b : _GEN_11976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11978 = 8'h4e == r_count_58_io_out ? io_r_78_b : _GEN_11977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11979 = 8'h4f == r_count_58_io_out ? io_r_79_b : _GEN_11978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11980 = 8'h50 == r_count_58_io_out ? io_r_80_b : _GEN_11979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11981 = 8'h51 == r_count_58_io_out ? io_r_81_b : _GEN_11980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11982 = 8'h52 == r_count_58_io_out ? io_r_82_b : _GEN_11981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11983 = 8'h53 == r_count_58_io_out ? io_r_83_b : _GEN_11982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11984 = 8'h54 == r_count_58_io_out ? io_r_84_b : _GEN_11983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11985 = 8'h55 == r_count_58_io_out ? io_r_85_b : _GEN_11984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11986 = 8'h56 == r_count_58_io_out ? io_r_86_b : _GEN_11985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11987 = 8'h57 == r_count_58_io_out ? io_r_87_b : _GEN_11986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11988 = 8'h58 == r_count_58_io_out ? io_r_88_b : _GEN_11987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11989 = 8'h59 == r_count_58_io_out ? io_r_89_b : _GEN_11988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11990 = 8'h5a == r_count_58_io_out ? io_r_90_b : _GEN_11989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11991 = 8'h5b == r_count_58_io_out ? io_r_91_b : _GEN_11990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11992 = 8'h5c == r_count_58_io_out ? io_r_92_b : _GEN_11991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11993 = 8'h5d == r_count_58_io_out ? io_r_93_b : _GEN_11992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11994 = 8'h5e == r_count_58_io_out ? io_r_94_b : _GEN_11993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11995 = 8'h5f == r_count_58_io_out ? io_r_95_b : _GEN_11994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11996 = 8'h60 == r_count_58_io_out ? io_r_96_b : _GEN_11995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11997 = 8'h61 == r_count_58_io_out ? io_r_97_b : _GEN_11996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11998 = 8'h62 == r_count_58_io_out ? io_r_98_b : _GEN_11997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_11999 = 8'h63 == r_count_58_io_out ? io_r_99_b : _GEN_11998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12000 = 8'h64 == r_count_58_io_out ? io_r_100_b : _GEN_11999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12001 = 8'h65 == r_count_58_io_out ? io_r_101_b : _GEN_12000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12002 = 8'h66 == r_count_58_io_out ? io_r_102_b : _GEN_12001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12003 = 8'h67 == r_count_58_io_out ? io_r_103_b : _GEN_12002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12004 = 8'h68 == r_count_58_io_out ? io_r_104_b : _GEN_12003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12005 = 8'h69 == r_count_58_io_out ? io_r_105_b : _GEN_12004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12006 = 8'h6a == r_count_58_io_out ? io_r_106_b : _GEN_12005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12007 = 8'h6b == r_count_58_io_out ? io_r_107_b : _GEN_12006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12008 = 8'h6c == r_count_58_io_out ? io_r_108_b : _GEN_12007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12009 = 8'h6d == r_count_58_io_out ? io_r_109_b : _GEN_12008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12010 = 8'h6e == r_count_58_io_out ? io_r_110_b : _GEN_12009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12011 = 8'h6f == r_count_58_io_out ? io_r_111_b : _GEN_12010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12012 = 8'h70 == r_count_58_io_out ? io_r_112_b : _GEN_12011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12013 = 8'h71 == r_count_58_io_out ? io_r_113_b : _GEN_12012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12014 = 8'h72 == r_count_58_io_out ? io_r_114_b : _GEN_12013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12015 = 8'h73 == r_count_58_io_out ? io_r_115_b : _GEN_12014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12016 = 8'h74 == r_count_58_io_out ? io_r_116_b : _GEN_12015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12017 = 8'h75 == r_count_58_io_out ? io_r_117_b : _GEN_12016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12018 = 8'h76 == r_count_58_io_out ? io_r_118_b : _GEN_12017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12019 = 8'h77 == r_count_58_io_out ? io_r_119_b : _GEN_12018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12020 = 8'h78 == r_count_58_io_out ? io_r_120_b : _GEN_12019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12021 = 8'h79 == r_count_58_io_out ? io_r_121_b : _GEN_12020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12022 = 8'h7a == r_count_58_io_out ? io_r_122_b : _GEN_12021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12023 = 8'h7b == r_count_58_io_out ? io_r_123_b : _GEN_12022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12024 = 8'h7c == r_count_58_io_out ? io_r_124_b : _GEN_12023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12025 = 8'h7d == r_count_58_io_out ? io_r_125_b : _GEN_12024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12026 = 8'h7e == r_count_58_io_out ? io_r_126_b : _GEN_12025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12027 = 8'h7f == r_count_58_io_out ? io_r_127_b : _GEN_12026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12028 = 8'h80 == r_count_58_io_out ? io_r_128_b : _GEN_12027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12029 = 8'h81 == r_count_58_io_out ? io_r_129_b : _GEN_12028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12030 = 8'h82 == r_count_58_io_out ? io_r_130_b : _GEN_12029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12031 = 8'h83 == r_count_58_io_out ? io_r_131_b : _GEN_12030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12032 = 8'h84 == r_count_58_io_out ? io_r_132_b : _GEN_12031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12033 = 8'h85 == r_count_58_io_out ? io_r_133_b : _GEN_12032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12034 = 8'h86 == r_count_58_io_out ? io_r_134_b : _GEN_12033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12035 = 8'h87 == r_count_58_io_out ? io_r_135_b : _GEN_12034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12036 = 8'h88 == r_count_58_io_out ? io_r_136_b : _GEN_12035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12037 = 8'h89 == r_count_58_io_out ? io_r_137_b : _GEN_12036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12038 = 8'h8a == r_count_58_io_out ? io_r_138_b : _GEN_12037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12039 = 8'h8b == r_count_58_io_out ? io_r_139_b : _GEN_12038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12040 = 8'h8c == r_count_58_io_out ? io_r_140_b : _GEN_12039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12041 = 8'h8d == r_count_58_io_out ? io_r_141_b : _GEN_12040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12042 = 8'h8e == r_count_58_io_out ? io_r_142_b : _GEN_12041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12043 = 8'h8f == r_count_58_io_out ? io_r_143_b : _GEN_12042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12044 = 8'h90 == r_count_58_io_out ? io_r_144_b : _GEN_12043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12045 = 8'h91 == r_count_58_io_out ? io_r_145_b : _GEN_12044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12046 = 8'h92 == r_count_58_io_out ? io_r_146_b : _GEN_12045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12047 = 8'h93 == r_count_58_io_out ? io_r_147_b : _GEN_12046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12048 = 8'h94 == r_count_58_io_out ? io_r_148_b : _GEN_12047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12049 = 8'h95 == r_count_58_io_out ? io_r_149_b : _GEN_12048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12050 = 8'h96 == r_count_58_io_out ? io_r_150_b : _GEN_12049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12051 = 8'h97 == r_count_58_io_out ? io_r_151_b : _GEN_12050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12052 = 8'h98 == r_count_58_io_out ? io_r_152_b : _GEN_12051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12053 = 8'h99 == r_count_58_io_out ? io_r_153_b : _GEN_12052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12054 = 8'h9a == r_count_58_io_out ? io_r_154_b : _GEN_12053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12055 = 8'h9b == r_count_58_io_out ? io_r_155_b : _GEN_12054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12056 = 8'h9c == r_count_58_io_out ? io_r_156_b : _GEN_12055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12057 = 8'h9d == r_count_58_io_out ? io_r_157_b : _GEN_12056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12058 = 8'h9e == r_count_58_io_out ? io_r_158_b : _GEN_12057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12059 = 8'h9f == r_count_58_io_out ? io_r_159_b : _GEN_12058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12060 = 8'ha0 == r_count_58_io_out ? io_r_160_b : _GEN_12059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12061 = 8'ha1 == r_count_58_io_out ? io_r_161_b : _GEN_12060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12062 = 8'ha2 == r_count_58_io_out ? io_r_162_b : _GEN_12061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12063 = 8'ha3 == r_count_58_io_out ? io_r_163_b : _GEN_12062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12064 = 8'ha4 == r_count_58_io_out ? io_r_164_b : _GEN_12063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12065 = 8'ha5 == r_count_58_io_out ? io_r_165_b : _GEN_12064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12066 = 8'ha6 == r_count_58_io_out ? io_r_166_b : _GEN_12065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12067 = 8'ha7 == r_count_58_io_out ? io_r_167_b : _GEN_12066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12068 = 8'ha8 == r_count_58_io_out ? io_r_168_b : _GEN_12067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12069 = 8'ha9 == r_count_58_io_out ? io_r_169_b : _GEN_12068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12070 = 8'haa == r_count_58_io_out ? io_r_170_b : _GEN_12069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12071 = 8'hab == r_count_58_io_out ? io_r_171_b : _GEN_12070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12072 = 8'hac == r_count_58_io_out ? io_r_172_b : _GEN_12071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12073 = 8'had == r_count_58_io_out ? io_r_173_b : _GEN_12072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12074 = 8'hae == r_count_58_io_out ? io_r_174_b : _GEN_12073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12075 = 8'haf == r_count_58_io_out ? io_r_175_b : _GEN_12074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12076 = 8'hb0 == r_count_58_io_out ? io_r_176_b : _GEN_12075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12077 = 8'hb1 == r_count_58_io_out ? io_r_177_b : _GEN_12076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12078 = 8'hb2 == r_count_58_io_out ? io_r_178_b : _GEN_12077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12079 = 8'hb3 == r_count_58_io_out ? io_r_179_b : _GEN_12078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12080 = 8'hb4 == r_count_58_io_out ? io_r_180_b : _GEN_12079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12081 = 8'hb5 == r_count_58_io_out ? io_r_181_b : _GEN_12080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12082 = 8'hb6 == r_count_58_io_out ? io_r_182_b : _GEN_12081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12083 = 8'hb7 == r_count_58_io_out ? io_r_183_b : _GEN_12082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12084 = 8'hb8 == r_count_58_io_out ? io_r_184_b : _GEN_12083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12085 = 8'hb9 == r_count_58_io_out ? io_r_185_b : _GEN_12084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12086 = 8'hba == r_count_58_io_out ? io_r_186_b : _GEN_12085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12087 = 8'hbb == r_count_58_io_out ? io_r_187_b : _GEN_12086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12088 = 8'hbc == r_count_58_io_out ? io_r_188_b : _GEN_12087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12089 = 8'hbd == r_count_58_io_out ? io_r_189_b : _GEN_12088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12090 = 8'hbe == r_count_58_io_out ? io_r_190_b : _GEN_12089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12091 = 8'hbf == r_count_58_io_out ? io_r_191_b : _GEN_12090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12092 = 8'hc0 == r_count_58_io_out ? io_r_192_b : _GEN_12091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12093 = 8'hc1 == r_count_58_io_out ? io_r_193_b : _GEN_12092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12094 = 8'hc2 == r_count_58_io_out ? io_r_194_b : _GEN_12093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12095 = 8'hc3 == r_count_58_io_out ? io_r_195_b : _GEN_12094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12096 = 8'hc4 == r_count_58_io_out ? io_r_196_b : _GEN_12095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12097 = 8'hc5 == r_count_58_io_out ? io_r_197_b : _GEN_12096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12098 = 8'hc6 == r_count_58_io_out ? io_r_198_b : _GEN_12097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12101 = 8'h1 == r_count_59_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12102 = 8'h2 == r_count_59_io_out ? io_r_2_b : _GEN_12101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12103 = 8'h3 == r_count_59_io_out ? io_r_3_b : _GEN_12102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12104 = 8'h4 == r_count_59_io_out ? io_r_4_b : _GEN_12103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12105 = 8'h5 == r_count_59_io_out ? io_r_5_b : _GEN_12104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12106 = 8'h6 == r_count_59_io_out ? io_r_6_b : _GEN_12105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12107 = 8'h7 == r_count_59_io_out ? io_r_7_b : _GEN_12106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12108 = 8'h8 == r_count_59_io_out ? io_r_8_b : _GEN_12107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12109 = 8'h9 == r_count_59_io_out ? io_r_9_b : _GEN_12108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12110 = 8'ha == r_count_59_io_out ? io_r_10_b : _GEN_12109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12111 = 8'hb == r_count_59_io_out ? io_r_11_b : _GEN_12110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12112 = 8'hc == r_count_59_io_out ? io_r_12_b : _GEN_12111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12113 = 8'hd == r_count_59_io_out ? io_r_13_b : _GEN_12112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12114 = 8'he == r_count_59_io_out ? io_r_14_b : _GEN_12113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12115 = 8'hf == r_count_59_io_out ? io_r_15_b : _GEN_12114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12116 = 8'h10 == r_count_59_io_out ? io_r_16_b : _GEN_12115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12117 = 8'h11 == r_count_59_io_out ? io_r_17_b : _GEN_12116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12118 = 8'h12 == r_count_59_io_out ? io_r_18_b : _GEN_12117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12119 = 8'h13 == r_count_59_io_out ? io_r_19_b : _GEN_12118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12120 = 8'h14 == r_count_59_io_out ? io_r_20_b : _GEN_12119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12121 = 8'h15 == r_count_59_io_out ? io_r_21_b : _GEN_12120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12122 = 8'h16 == r_count_59_io_out ? io_r_22_b : _GEN_12121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12123 = 8'h17 == r_count_59_io_out ? io_r_23_b : _GEN_12122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12124 = 8'h18 == r_count_59_io_out ? io_r_24_b : _GEN_12123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12125 = 8'h19 == r_count_59_io_out ? io_r_25_b : _GEN_12124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12126 = 8'h1a == r_count_59_io_out ? io_r_26_b : _GEN_12125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12127 = 8'h1b == r_count_59_io_out ? io_r_27_b : _GEN_12126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12128 = 8'h1c == r_count_59_io_out ? io_r_28_b : _GEN_12127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12129 = 8'h1d == r_count_59_io_out ? io_r_29_b : _GEN_12128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12130 = 8'h1e == r_count_59_io_out ? io_r_30_b : _GEN_12129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12131 = 8'h1f == r_count_59_io_out ? io_r_31_b : _GEN_12130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12132 = 8'h20 == r_count_59_io_out ? io_r_32_b : _GEN_12131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12133 = 8'h21 == r_count_59_io_out ? io_r_33_b : _GEN_12132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12134 = 8'h22 == r_count_59_io_out ? io_r_34_b : _GEN_12133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12135 = 8'h23 == r_count_59_io_out ? io_r_35_b : _GEN_12134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12136 = 8'h24 == r_count_59_io_out ? io_r_36_b : _GEN_12135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12137 = 8'h25 == r_count_59_io_out ? io_r_37_b : _GEN_12136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12138 = 8'h26 == r_count_59_io_out ? io_r_38_b : _GEN_12137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12139 = 8'h27 == r_count_59_io_out ? io_r_39_b : _GEN_12138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12140 = 8'h28 == r_count_59_io_out ? io_r_40_b : _GEN_12139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12141 = 8'h29 == r_count_59_io_out ? io_r_41_b : _GEN_12140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12142 = 8'h2a == r_count_59_io_out ? io_r_42_b : _GEN_12141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12143 = 8'h2b == r_count_59_io_out ? io_r_43_b : _GEN_12142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12144 = 8'h2c == r_count_59_io_out ? io_r_44_b : _GEN_12143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12145 = 8'h2d == r_count_59_io_out ? io_r_45_b : _GEN_12144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12146 = 8'h2e == r_count_59_io_out ? io_r_46_b : _GEN_12145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12147 = 8'h2f == r_count_59_io_out ? io_r_47_b : _GEN_12146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12148 = 8'h30 == r_count_59_io_out ? io_r_48_b : _GEN_12147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12149 = 8'h31 == r_count_59_io_out ? io_r_49_b : _GEN_12148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12150 = 8'h32 == r_count_59_io_out ? io_r_50_b : _GEN_12149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12151 = 8'h33 == r_count_59_io_out ? io_r_51_b : _GEN_12150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12152 = 8'h34 == r_count_59_io_out ? io_r_52_b : _GEN_12151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12153 = 8'h35 == r_count_59_io_out ? io_r_53_b : _GEN_12152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12154 = 8'h36 == r_count_59_io_out ? io_r_54_b : _GEN_12153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12155 = 8'h37 == r_count_59_io_out ? io_r_55_b : _GEN_12154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12156 = 8'h38 == r_count_59_io_out ? io_r_56_b : _GEN_12155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12157 = 8'h39 == r_count_59_io_out ? io_r_57_b : _GEN_12156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12158 = 8'h3a == r_count_59_io_out ? io_r_58_b : _GEN_12157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12159 = 8'h3b == r_count_59_io_out ? io_r_59_b : _GEN_12158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12160 = 8'h3c == r_count_59_io_out ? io_r_60_b : _GEN_12159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12161 = 8'h3d == r_count_59_io_out ? io_r_61_b : _GEN_12160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12162 = 8'h3e == r_count_59_io_out ? io_r_62_b : _GEN_12161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12163 = 8'h3f == r_count_59_io_out ? io_r_63_b : _GEN_12162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12164 = 8'h40 == r_count_59_io_out ? io_r_64_b : _GEN_12163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12165 = 8'h41 == r_count_59_io_out ? io_r_65_b : _GEN_12164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12166 = 8'h42 == r_count_59_io_out ? io_r_66_b : _GEN_12165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12167 = 8'h43 == r_count_59_io_out ? io_r_67_b : _GEN_12166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12168 = 8'h44 == r_count_59_io_out ? io_r_68_b : _GEN_12167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12169 = 8'h45 == r_count_59_io_out ? io_r_69_b : _GEN_12168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12170 = 8'h46 == r_count_59_io_out ? io_r_70_b : _GEN_12169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12171 = 8'h47 == r_count_59_io_out ? io_r_71_b : _GEN_12170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12172 = 8'h48 == r_count_59_io_out ? io_r_72_b : _GEN_12171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12173 = 8'h49 == r_count_59_io_out ? io_r_73_b : _GEN_12172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12174 = 8'h4a == r_count_59_io_out ? io_r_74_b : _GEN_12173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12175 = 8'h4b == r_count_59_io_out ? io_r_75_b : _GEN_12174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12176 = 8'h4c == r_count_59_io_out ? io_r_76_b : _GEN_12175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12177 = 8'h4d == r_count_59_io_out ? io_r_77_b : _GEN_12176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12178 = 8'h4e == r_count_59_io_out ? io_r_78_b : _GEN_12177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12179 = 8'h4f == r_count_59_io_out ? io_r_79_b : _GEN_12178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12180 = 8'h50 == r_count_59_io_out ? io_r_80_b : _GEN_12179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12181 = 8'h51 == r_count_59_io_out ? io_r_81_b : _GEN_12180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12182 = 8'h52 == r_count_59_io_out ? io_r_82_b : _GEN_12181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12183 = 8'h53 == r_count_59_io_out ? io_r_83_b : _GEN_12182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12184 = 8'h54 == r_count_59_io_out ? io_r_84_b : _GEN_12183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12185 = 8'h55 == r_count_59_io_out ? io_r_85_b : _GEN_12184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12186 = 8'h56 == r_count_59_io_out ? io_r_86_b : _GEN_12185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12187 = 8'h57 == r_count_59_io_out ? io_r_87_b : _GEN_12186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12188 = 8'h58 == r_count_59_io_out ? io_r_88_b : _GEN_12187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12189 = 8'h59 == r_count_59_io_out ? io_r_89_b : _GEN_12188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12190 = 8'h5a == r_count_59_io_out ? io_r_90_b : _GEN_12189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12191 = 8'h5b == r_count_59_io_out ? io_r_91_b : _GEN_12190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12192 = 8'h5c == r_count_59_io_out ? io_r_92_b : _GEN_12191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12193 = 8'h5d == r_count_59_io_out ? io_r_93_b : _GEN_12192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12194 = 8'h5e == r_count_59_io_out ? io_r_94_b : _GEN_12193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12195 = 8'h5f == r_count_59_io_out ? io_r_95_b : _GEN_12194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12196 = 8'h60 == r_count_59_io_out ? io_r_96_b : _GEN_12195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12197 = 8'h61 == r_count_59_io_out ? io_r_97_b : _GEN_12196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12198 = 8'h62 == r_count_59_io_out ? io_r_98_b : _GEN_12197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12199 = 8'h63 == r_count_59_io_out ? io_r_99_b : _GEN_12198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12200 = 8'h64 == r_count_59_io_out ? io_r_100_b : _GEN_12199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12201 = 8'h65 == r_count_59_io_out ? io_r_101_b : _GEN_12200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12202 = 8'h66 == r_count_59_io_out ? io_r_102_b : _GEN_12201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12203 = 8'h67 == r_count_59_io_out ? io_r_103_b : _GEN_12202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12204 = 8'h68 == r_count_59_io_out ? io_r_104_b : _GEN_12203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12205 = 8'h69 == r_count_59_io_out ? io_r_105_b : _GEN_12204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12206 = 8'h6a == r_count_59_io_out ? io_r_106_b : _GEN_12205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12207 = 8'h6b == r_count_59_io_out ? io_r_107_b : _GEN_12206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12208 = 8'h6c == r_count_59_io_out ? io_r_108_b : _GEN_12207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12209 = 8'h6d == r_count_59_io_out ? io_r_109_b : _GEN_12208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12210 = 8'h6e == r_count_59_io_out ? io_r_110_b : _GEN_12209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12211 = 8'h6f == r_count_59_io_out ? io_r_111_b : _GEN_12210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12212 = 8'h70 == r_count_59_io_out ? io_r_112_b : _GEN_12211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12213 = 8'h71 == r_count_59_io_out ? io_r_113_b : _GEN_12212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12214 = 8'h72 == r_count_59_io_out ? io_r_114_b : _GEN_12213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12215 = 8'h73 == r_count_59_io_out ? io_r_115_b : _GEN_12214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12216 = 8'h74 == r_count_59_io_out ? io_r_116_b : _GEN_12215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12217 = 8'h75 == r_count_59_io_out ? io_r_117_b : _GEN_12216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12218 = 8'h76 == r_count_59_io_out ? io_r_118_b : _GEN_12217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12219 = 8'h77 == r_count_59_io_out ? io_r_119_b : _GEN_12218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12220 = 8'h78 == r_count_59_io_out ? io_r_120_b : _GEN_12219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12221 = 8'h79 == r_count_59_io_out ? io_r_121_b : _GEN_12220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12222 = 8'h7a == r_count_59_io_out ? io_r_122_b : _GEN_12221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12223 = 8'h7b == r_count_59_io_out ? io_r_123_b : _GEN_12222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12224 = 8'h7c == r_count_59_io_out ? io_r_124_b : _GEN_12223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12225 = 8'h7d == r_count_59_io_out ? io_r_125_b : _GEN_12224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12226 = 8'h7e == r_count_59_io_out ? io_r_126_b : _GEN_12225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12227 = 8'h7f == r_count_59_io_out ? io_r_127_b : _GEN_12226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12228 = 8'h80 == r_count_59_io_out ? io_r_128_b : _GEN_12227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12229 = 8'h81 == r_count_59_io_out ? io_r_129_b : _GEN_12228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12230 = 8'h82 == r_count_59_io_out ? io_r_130_b : _GEN_12229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12231 = 8'h83 == r_count_59_io_out ? io_r_131_b : _GEN_12230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12232 = 8'h84 == r_count_59_io_out ? io_r_132_b : _GEN_12231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12233 = 8'h85 == r_count_59_io_out ? io_r_133_b : _GEN_12232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12234 = 8'h86 == r_count_59_io_out ? io_r_134_b : _GEN_12233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12235 = 8'h87 == r_count_59_io_out ? io_r_135_b : _GEN_12234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12236 = 8'h88 == r_count_59_io_out ? io_r_136_b : _GEN_12235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12237 = 8'h89 == r_count_59_io_out ? io_r_137_b : _GEN_12236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12238 = 8'h8a == r_count_59_io_out ? io_r_138_b : _GEN_12237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12239 = 8'h8b == r_count_59_io_out ? io_r_139_b : _GEN_12238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12240 = 8'h8c == r_count_59_io_out ? io_r_140_b : _GEN_12239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12241 = 8'h8d == r_count_59_io_out ? io_r_141_b : _GEN_12240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12242 = 8'h8e == r_count_59_io_out ? io_r_142_b : _GEN_12241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12243 = 8'h8f == r_count_59_io_out ? io_r_143_b : _GEN_12242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12244 = 8'h90 == r_count_59_io_out ? io_r_144_b : _GEN_12243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12245 = 8'h91 == r_count_59_io_out ? io_r_145_b : _GEN_12244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12246 = 8'h92 == r_count_59_io_out ? io_r_146_b : _GEN_12245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12247 = 8'h93 == r_count_59_io_out ? io_r_147_b : _GEN_12246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12248 = 8'h94 == r_count_59_io_out ? io_r_148_b : _GEN_12247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12249 = 8'h95 == r_count_59_io_out ? io_r_149_b : _GEN_12248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12250 = 8'h96 == r_count_59_io_out ? io_r_150_b : _GEN_12249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12251 = 8'h97 == r_count_59_io_out ? io_r_151_b : _GEN_12250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12252 = 8'h98 == r_count_59_io_out ? io_r_152_b : _GEN_12251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12253 = 8'h99 == r_count_59_io_out ? io_r_153_b : _GEN_12252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12254 = 8'h9a == r_count_59_io_out ? io_r_154_b : _GEN_12253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12255 = 8'h9b == r_count_59_io_out ? io_r_155_b : _GEN_12254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12256 = 8'h9c == r_count_59_io_out ? io_r_156_b : _GEN_12255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12257 = 8'h9d == r_count_59_io_out ? io_r_157_b : _GEN_12256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12258 = 8'h9e == r_count_59_io_out ? io_r_158_b : _GEN_12257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12259 = 8'h9f == r_count_59_io_out ? io_r_159_b : _GEN_12258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12260 = 8'ha0 == r_count_59_io_out ? io_r_160_b : _GEN_12259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12261 = 8'ha1 == r_count_59_io_out ? io_r_161_b : _GEN_12260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12262 = 8'ha2 == r_count_59_io_out ? io_r_162_b : _GEN_12261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12263 = 8'ha3 == r_count_59_io_out ? io_r_163_b : _GEN_12262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12264 = 8'ha4 == r_count_59_io_out ? io_r_164_b : _GEN_12263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12265 = 8'ha5 == r_count_59_io_out ? io_r_165_b : _GEN_12264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12266 = 8'ha6 == r_count_59_io_out ? io_r_166_b : _GEN_12265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12267 = 8'ha7 == r_count_59_io_out ? io_r_167_b : _GEN_12266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12268 = 8'ha8 == r_count_59_io_out ? io_r_168_b : _GEN_12267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12269 = 8'ha9 == r_count_59_io_out ? io_r_169_b : _GEN_12268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12270 = 8'haa == r_count_59_io_out ? io_r_170_b : _GEN_12269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12271 = 8'hab == r_count_59_io_out ? io_r_171_b : _GEN_12270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12272 = 8'hac == r_count_59_io_out ? io_r_172_b : _GEN_12271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12273 = 8'had == r_count_59_io_out ? io_r_173_b : _GEN_12272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12274 = 8'hae == r_count_59_io_out ? io_r_174_b : _GEN_12273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12275 = 8'haf == r_count_59_io_out ? io_r_175_b : _GEN_12274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12276 = 8'hb0 == r_count_59_io_out ? io_r_176_b : _GEN_12275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12277 = 8'hb1 == r_count_59_io_out ? io_r_177_b : _GEN_12276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12278 = 8'hb2 == r_count_59_io_out ? io_r_178_b : _GEN_12277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12279 = 8'hb3 == r_count_59_io_out ? io_r_179_b : _GEN_12278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12280 = 8'hb4 == r_count_59_io_out ? io_r_180_b : _GEN_12279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12281 = 8'hb5 == r_count_59_io_out ? io_r_181_b : _GEN_12280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12282 = 8'hb6 == r_count_59_io_out ? io_r_182_b : _GEN_12281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12283 = 8'hb7 == r_count_59_io_out ? io_r_183_b : _GEN_12282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12284 = 8'hb8 == r_count_59_io_out ? io_r_184_b : _GEN_12283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12285 = 8'hb9 == r_count_59_io_out ? io_r_185_b : _GEN_12284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12286 = 8'hba == r_count_59_io_out ? io_r_186_b : _GEN_12285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12287 = 8'hbb == r_count_59_io_out ? io_r_187_b : _GEN_12286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12288 = 8'hbc == r_count_59_io_out ? io_r_188_b : _GEN_12287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12289 = 8'hbd == r_count_59_io_out ? io_r_189_b : _GEN_12288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12290 = 8'hbe == r_count_59_io_out ? io_r_190_b : _GEN_12289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12291 = 8'hbf == r_count_59_io_out ? io_r_191_b : _GEN_12290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12292 = 8'hc0 == r_count_59_io_out ? io_r_192_b : _GEN_12291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12293 = 8'hc1 == r_count_59_io_out ? io_r_193_b : _GEN_12292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12294 = 8'hc2 == r_count_59_io_out ? io_r_194_b : _GEN_12293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12295 = 8'hc3 == r_count_59_io_out ? io_r_195_b : _GEN_12294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12296 = 8'hc4 == r_count_59_io_out ? io_r_196_b : _GEN_12295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12297 = 8'hc5 == r_count_59_io_out ? io_r_197_b : _GEN_12296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12298 = 8'hc6 == r_count_59_io_out ? io_r_198_b : _GEN_12297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12301 = 8'h1 == r_count_60_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12302 = 8'h2 == r_count_60_io_out ? io_r_2_b : _GEN_12301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12303 = 8'h3 == r_count_60_io_out ? io_r_3_b : _GEN_12302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12304 = 8'h4 == r_count_60_io_out ? io_r_4_b : _GEN_12303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12305 = 8'h5 == r_count_60_io_out ? io_r_5_b : _GEN_12304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12306 = 8'h6 == r_count_60_io_out ? io_r_6_b : _GEN_12305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12307 = 8'h7 == r_count_60_io_out ? io_r_7_b : _GEN_12306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12308 = 8'h8 == r_count_60_io_out ? io_r_8_b : _GEN_12307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12309 = 8'h9 == r_count_60_io_out ? io_r_9_b : _GEN_12308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12310 = 8'ha == r_count_60_io_out ? io_r_10_b : _GEN_12309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12311 = 8'hb == r_count_60_io_out ? io_r_11_b : _GEN_12310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12312 = 8'hc == r_count_60_io_out ? io_r_12_b : _GEN_12311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12313 = 8'hd == r_count_60_io_out ? io_r_13_b : _GEN_12312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12314 = 8'he == r_count_60_io_out ? io_r_14_b : _GEN_12313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12315 = 8'hf == r_count_60_io_out ? io_r_15_b : _GEN_12314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12316 = 8'h10 == r_count_60_io_out ? io_r_16_b : _GEN_12315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12317 = 8'h11 == r_count_60_io_out ? io_r_17_b : _GEN_12316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12318 = 8'h12 == r_count_60_io_out ? io_r_18_b : _GEN_12317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12319 = 8'h13 == r_count_60_io_out ? io_r_19_b : _GEN_12318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12320 = 8'h14 == r_count_60_io_out ? io_r_20_b : _GEN_12319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12321 = 8'h15 == r_count_60_io_out ? io_r_21_b : _GEN_12320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12322 = 8'h16 == r_count_60_io_out ? io_r_22_b : _GEN_12321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12323 = 8'h17 == r_count_60_io_out ? io_r_23_b : _GEN_12322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12324 = 8'h18 == r_count_60_io_out ? io_r_24_b : _GEN_12323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12325 = 8'h19 == r_count_60_io_out ? io_r_25_b : _GEN_12324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12326 = 8'h1a == r_count_60_io_out ? io_r_26_b : _GEN_12325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12327 = 8'h1b == r_count_60_io_out ? io_r_27_b : _GEN_12326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12328 = 8'h1c == r_count_60_io_out ? io_r_28_b : _GEN_12327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12329 = 8'h1d == r_count_60_io_out ? io_r_29_b : _GEN_12328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12330 = 8'h1e == r_count_60_io_out ? io_r_30_b : _GEN_12329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12331 = 8'h1f == r_count_60_io_out ? io_r_31_b : _GEN_12330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12332 = 8'h20 == r_count_60_io_out ? io_r_32_b : _GEN_12331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12333 = 8'h21 == r_count_60_io_out ? io_r_33_b : _GEN_12332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12334 = 8'h22 == r_count_60_io_out ? io_r_34_b : _GEN_12333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12335 = 8'h23 == r_count_60_io_out ? io_r_35_b : _GEN_12334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12336 = 8'h24 == r_count_60_io_out ? io_r_36_b : _GEN_12335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12337 = 8'h25 == r_count_60_io_out ? io_r_37_b : _GEN_12336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12338 = 8'h26 == r_count_60_io_out ? io_r_38_b : _GEN_12337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12339 = 8'h27 == r_count_60_io_out ? io_r_39_b : _GEN_12338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12340 = 8'h28 == r_count_60_io_out ? io_r_40_b : _GEN_12339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12341 = 8'h29 == r_count_60_io_out ? io_r_41_b : _GEN_12340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12342 = 8'h2a == r_count_60_io_out ? io_r_42_b : _GEN_12341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12343 = 8'h2b == r_count_60_io_out ? io_r_43_b : _GEN_12342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12344 = 8'h2c == r_count_60_io_out ? io_r_44_b : _GEN_12343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12345 = 8'h2d == r_count_60_io_out ? io_r_45_b : _GEN_12344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12346 = 8'h2e == r_count_60_io_out ? io_r_46_b : _GEN_12345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12347 = 8'h2f == r_count_60_io_out ? io_r_47_b : _GEN_12346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12348 = 8'h30 == r_count_60_io_out ? io_r_48_b : _GEN_12347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12349 = 8'h31 == r_count_60_io_out ? io_r_49_b : _GEN_12348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12350 = 8'h32 == r_count_60_io_out ? io_r_50_b : _GEN_12349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12351 = 8'h33 == r_count_60_io_out ? io_r_51_b : _GEN_12350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12352 = 8'h34 == r_count_60_io_out ? io_r_52_b : _GEN_12351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12353 = 8'h35 == r_count_60_io_out ? io_r_53_b : _GEN_12352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12354 = 8'h36 == r_count_60_io_out ? io_r_54_b : _GEN_12353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12355 = 8'h37 == r_count_60_io_out ? io_r_55_b : _GEN_12354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12356 = 8'h38 == r_count_60_io_out ? io_r_56_b : _GEN_12355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12357 = 8'h39 == r_count_60_io_out ? io_r_57_b : _GEN_12356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12358 = 8'h3a == r_count_60_io_out ? io_r_58_b : _GEN_12357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12359 = 8'h3b == r_count_60_io_out ? io_r_59_b : _GEN_12358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12360 = 8'h3c == r_count_60_io_out ? io_r_60_b : _GEN_12359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12361 = 8'h3d == r_count_60_io_out ? io_r_61_b : _GEN_12360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12362 = 8'h3e == r_count_60_io_out ? io_r_62_b : _GEN_12361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12363 = 8'h3f == r_count_60_io_out ? io_r_63_b : _GEN_12362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12364 = 8'h40 == r_count_60_io_out ? io_r_64_b : _GEN_12363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12365 = 8'h41 == r_count_60_io_out ? io_r_65_b : _GEN_12364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12366 = 8'h42 == r_count_60_io_out ? io_r_66_b : _GEN_12365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12367 = 8'h43 == r_count_60_io_out ? io_r_67_b : _GEN_12366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12368 = 8'h44 == r_count_60_io_out ? io_r_68_b : _GEN_12367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12369 = 8'h45 == r_count_60_io_out ? io_r_69_b : _GEN_12368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12370 = 8'h46 == r_count_60_io_out ? io_r_70_b : _GEN_12369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12371 = 8'h47 == r_count_60_io_out ? io_r_71_b : _GEN_12370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12372 = 8'h48 == r_count_60_io_out ? io_r_72_b : _GEN_12371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12373 = 8'h49 == r_count_60_io_out ? io_r_73_b : _GEN_12372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12374 = 8'h4a == r_count_60_io_out ? io_r_74_b : _GEN_12373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12375 = 8'h4b == r_count_60_io_out ? io_r_75_b : _GEN_12374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12376 = 8'h4c == r_count_60_io_out ? io_r_76_b : _GEN_12375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12377 = 8'h4d == r_count_60_io_out ? io_r_77_b : _GEN_12376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12378 = 8'h4e == r_count_60_io_out ? io_r_78_b : _GEN_12377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12379 = 8'h4f == r_count_60_io_out ? io_r_79_b : _GEN_12378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12380 = 8'h50 == r_count_60_io_out ? io_r_80_b : _GEN_12379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12381 = 8'h51 == r_count_60_io_out ? io_r_81_b : _GEN_12380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12382 = 8'h52 == r_count_60_io_out ? io_r_82_b : _GEN_12381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12383 = 8'h53 == r_count_60_io_out ? io_r_83_b : _GEN_12382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12384 = 8'h54 == r_count_60_io_out ? io_r_84_b : _GEN_12383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12385 = 8'h55 == r_count_60_io_out ? io_r_85_b : _GEN_12384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12386 = 8'h56 == r_count_60_io_out ? io_r_86_b : _GEN_12385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12387 = 8'h57 == r_count_60_io_out ? io_r_87_b : _GEN_12386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12388 = 8'h58 == r_count_60_io_out ? io_r_88_b : _GEN_12387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12389 = 8'h59 == r_count_60_io_out ? io_r_89_b : _GEN_12388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12390 = 8'h5a == r_count_60_io_out ? io_r_90_b : _GEN_12389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12391 = 8'h5b == r_count_60_io_out ? io_r_91_b : _GEN_12390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12392 = 8'h5c == r_count_60_io_out ? io_r_92_b : _GEN_12391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12393 = 8'h5d == r_count_60_io_out ? io_r_93_b : _GEN_12392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12394 = 8'h5e == r_count_60_io_out ? io_r_94_b : _GEN_12393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12395 = 8'h5f == r_count_60_io_out ? io_r_95_b : _GEN_12394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12396 = 8'h60 == r_count_60_io_out ? io_r_96_b : _GEN_12395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12397 = 8'h61 == r_count_60_io_out ? io_r_97_b : _GEN_12396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12398 = 8'h62 == r_count_60_io_out ? io_r_98_b : _GEN_12397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12399 = 8'h63 == r_count_60_io_out ? io_r_99_b : _GEN_12398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12400 = 8'h64 == r_count_60_io_out ? io_r_100_b : _GEN_12399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12401 = 8'h65 == r_count_60_io_out ? io_r_101_b : _GEN_12400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12402 = 8'h66 == r_count_60_io_out ? io_r_102_b : _GEN_12401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12403 = 8'h67 == r_count_60_io_out ? io_r_103_b : _GEN_12402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12404 = 8'h68 == r_count_60_io_out ? io_r_104_b : _GEN_12403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12405 = 8'h69 == r_count_60_io_out ? io_r_105_b : _GEN_12404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12406 = 8'h6a == r_count_60_io_out ? io_r_106_b : _GEN_12405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12407 = 8'h6b == r_count_60_io_out ? io_r_107_b : _GEN_12406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12408 = 8'h6c == r_count_60_io_out ? io_r_108_b : _GEN_12407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12409 = 8'h6d == r_count_60_io_out ? io_r_109_b : _GEN_12408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12410 = 8'h6e == r_count_60_io_out ? io_r_110_b : _GEN_12409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12411 = 8'h6f == r_count_60_io_out ? io_r_111_b : _GEN_12410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12412 = 8'h70 == r_count_60_io_out ? io_r_112_b : _GEN_12411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12413 = 8'h71 == r_count_60_io_out ? io_r_113_b : _GEN_12412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12414 = 8'h72 == r_count_60_io_out ? io_r_114_b : _GEN_12413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12415 = 8'h73 == r_count_60_io_out ? io_r_115_b : _GEN_12414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12416 = 8'h74 == r_count_60_io_out ? io_r_116_b : _GEN_12415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12417 = 8'h75 == r_count_60_io_out ? io_r_117_b : _GEN_12416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12418 = 8'h76 == r_count_60_io_out ? io_r_118_b : _GEN_12417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12419 = 8'h77 == r_count_60_io_out ? io_r_119_b : _GEN_12418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12420 = 8'h78 == r_count_60_io_out ? io_r_120_b : _GEN_12419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12421 = 8'h79 == r_count_60_io_out ? io_r_121_b : _GEN_12420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12422 = 8'h7a == r_count_60_io_out ? io_r_122_b : _GEN_12421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12423 = 8'h7b == r_count_60_io_out ? io_r_123_b : _GEN_12422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12424 = 8'h7c == r_count_60_io_out ? io_r_124_b : _GEN_12423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12425 = 8'h7d == r_count_60_io_out ? io_r_125_b : _GEN_12424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12426 = 8'h7e == r_count_60_io_out ? io_r_126_b : _GEN_12425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12427 = 8'h7f == r_count_60_io_out ? io_r_127_b : _GEN_12426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12428 = 8'h80 == r_count_60_io_out ? io_r_128_b : _GEN_12427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12429 = 8'h81 == r_count_60_io_out ? io_r_129_b : _GEN_12428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12430 = 8'h82 == r_count_60_io_out ? io_r_130_b : _GEN_12429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12431 = 8'h83 == r_count_60_io_out ? io_r_131_b : _GEN_12430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12432 = 8'h84 == r_count_60_io_out ? io_r_132_b : _GEN_12431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12433 = 8'h85 == r_count_60_io_out ? io_r_133_b : _GEN_12432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12434 = 8'h86 == r_count_60_io_out ? io_r_134_b : _GEN_12433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12435 = 8'h87 == r_count_60_io_out ? io_r_135_b : _GEN_12434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12436 = 8'h88 == r_count_60_io_out ? io_r_136_b : _GEN_12435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12437 = 8'h89 == r_count_60_io_out ? io_r_137_b : _GEN_12436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12438 = 8'h8a == r_count_60_io_out ? io_r_138_b : _GEN_12437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12439 = 8'h8b == r_count_60_io_out ? io_r_139_b : _GEN_12438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12440 = 8'h8c == r_count_60_io_out ? io_r_140_b : _GEN_12439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12441 = 8'h8d == r_count_60_io_out ? io_r_141_b : _GEN_12440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12442 = 8'h8e == r_count_60_io_out ? io_r_142_b : _GEN_12441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12443 = 8'h8f == r_count_60_io_out ? io_r_143_b : _GEN_12442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12444 = 8'h90 == r_count_60_io_out ? io_r_144_b : _GEN_12443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12445 = 8'h91 == r_count_60_io_out ? io_r_145_b : _GEN_12444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12446 = 8'h92 == r_count_60_io_out ? io_r_146_b : _GEN_12445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12447 = 8'h93 == r_count_60_io_out ? io_r_147_b : _GEN_12446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12448 = 8'h94 == r_count_60_io_out ? io_r_148_b : _GEN_12447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12449 = 8'h95 == r_count_60_io_out ? io_r_149_b : _GEN_12448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12450 = 8'h96 == r_count_60_io_out ? io_r_150_b : _GEN_12449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12451 = 8'h97 == r_count_60_io_out ? io_r_151_b : _GEN_12450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12452 = 8'h98 == r_count_60_io_out ? io_r_152_b : _GEN_12451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12453 = 8'h99 == r_count_60_io_out ? io_r_153_b : _GEN_12452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12454 = 8'h9a == r_count_60_io_out ? io_r_154_b : _GEN_12453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12455 = 8'h9b == r_count_60_io_out ? io_r_155_b : _GEN_12454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12456 = 8'h9c == r_count_60_io_out ? io_r_156_b : _GEN_12455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12457 = 8'h9d == r_count_60_io_out ? io_r_157_b : _GEN_12456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12458 = 8'h9e == r_count_60_io_out ? io_r_158_b : _GEN_12457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12459 = 8'h9f == r_count_60_io_out ? io_r_159_b : _GEN_12458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12460 = 8'ha0 == r_count_60_io_out ? io_r_160_b : _GEN_12459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12461 = 8'ha1 == r_count_60_io_out ? io_r_161_b : _GEN_12460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12462 = 8'ha2 == r_count_60_io_out ? io_r_162_b : _GEN_12461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12463 = 8'ha3 == r_count_60_io_out ? io_r_163_b : _GEN_12462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12464 = 8'ha4 == r_count_60_io_out ? io_r_164_b : _GEN_12463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12465 = 8'ha5 == r_count_60_io_out ? io_r_165_b : _GEN_12464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12466 = 8'ha6 == r_count_60_io_out ? io_r_166_b : _GEN_12465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12467 = 8'ha7 == r_count_60_io_out ? io_r_167_b : _GEN_12466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12468 = 8'ha8 == r_count_60_io_out ? io_r_168_b : _GEN_12467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12469 = 8'ha9 == r_count_60_io_out ? io_r_169_b : _GEN_12468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12470 = 8'haa == r_count_60_io_out ? io_r_170_b : _GEN_12469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12471 = 8'hab == r_count_60_io_out ? io_r_171_b : _GEN_12470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12472 = 8'hac == r_count_60_io_out ? io_r_172_b : _GEN_12471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12473 = 8'had == r_count_60_io_out ? io_r_173_b : _GEN_12472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12474 = 8'hae == r_count_60_io_out ? io_r_174_b : _GEN_12473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12475 = 8'haf == r_count_60_io_out ? io_r_175_b : _GEN_12474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12476 = 8'hb0 == r_count_60_io_out ? io_r_176_b : _GEN_12475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12477 = 8'hb1 == r_count_60_io_out ? io_r_177_b : _GEN_12476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12478 = 8'hb2 == r_count_60_io_out ? io_r_178_b : _GEN_12477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12479 = 8'hb3 == r_count_60_io_out ? io_r_179_b : _GEN_12478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12480 = 8'hb4 == r_count_60_io_out ? io_r_180_b : _GEN_12479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12481 = 8'hb5 == r_count_60_io_out ? io_r_181_b : _GEN_12480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12482 = 8'hb6 == r_count_60_io_out ? io_r_182_b : _GEN_12481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12483 = 8'hb7 == r_count_60_io_out ? io_r_183_b : _GEN_12482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12484 = 8'hb8 == r_count_60_io_out ? io_r_184_b : _GEN_12483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12485 = 8'hb9 == r_count_60_io_out ? io_r_185_b : _GEN_12484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12486 = 8'hba == r_count_60_io_out ? io_r_186_b : _GEN_12485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12487 = 8'hbb == r_count_60_io_out ? io_r_187_b : _GEN_12486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12488 = 8'hbc == r_count_60_io_out ? io_r_188_b : _GEN_12487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12489 = 8'hbd == r_count_60_io_out ? io_r_189_b : _GEN_12488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12490 = 8'hbe == r_count_60_io_out ? io_r_190_b : _GEN_12489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12491 = 8'hbf == r_count_60_io_out ? io_r_191_b : _GEN_12490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12492 = 8'hc0 == r_count_60_io_out ? io_r_192_b : _GEN_12491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12493 = 8'hc1 == r_count_60_io_out ? io_r_193_b : _GEN_12492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12494 = 8'hc2 == r_count_60_io_out ? io_r_194_b : _GEN_12493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12495 = 8'hc3 == r_count_60_io_out ? io_r_195_b : _GEN_12494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12496 = 8'hc4 == r_count_60_io_out ? io_r_196_b : _GEN_12495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12497 = 8'hc5 == r_count_60_io_out ? io_r_197_b : _GEN_12496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12498 = 8'hc6 == r_count_60_io_out ? io_r_198_b : _GEN_12497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12501 = 8'h1 == r_count_61_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12502 = 8'h2 == r_count_61_io_out ? io_r_2_b : _GEN_12501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12503 = 8'h3 == r_count_61_io_out ? io_r_3_b : _GEN_12502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12504 = 8'h4 == r_count_61_io_out ? io_r_4_b : _GEN_12503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12505 = 8'h5 == r_count_61_io_out ? io_r_5_b : _GEN_12504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12506 = 8'h6 == r_count_61_io_out ? io_r_6_b : _GEN_12505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12507 = 8'h7 == r_count_61_io_out ? io_r_7_b : _GEN_12506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12508 = 8'h8 == r_count_61_io_out ? io_r_8_b : _GEN_12507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12509 = 8'h9 == r_count_61_io_out ? io_r_9_b : _GEN_12508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12510 = 8'ha == r_count_61_io_out ? io_r_10_b : _GEN_12509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12511 = 8'hb == r_count_61_io_out ? io_r_11_b : _GEN_12510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12512 = 8'hc == r_count_61_io_out ? io_r_12_b : _GEN_12511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12513 = 8'hd == r_count_61_io_out ? io_r_13_b : _GEN_12512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12514 = 8'he == r_count_61_io_out ? io_r_14_b : _GEN_12513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12515 = 8'hf == r_count_61_io_out ? io_r_15_b : _GEN_12514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12516 = 8'h10 == r_count_61_io_out ? io_r_16_b : _GEN_12515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12517 = 8'h11 == r_count_61_io_out ? io_r_17_b : _GEN_12516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12518 = 8'h12 == r_count_61_io_out ? io_r_18_b : _GEN_12517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12519 = 8'h13 == r_count_61_io_out ? io_r_19_b : _GEN_12518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12520 = 8'h14 == r_count_61_io_out ? io_r_20_b : _GEN_12519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12521 = 8'h15 == r_count_61_io_out ? io_r_21_b : _GEN_12520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12522 = 8'h16 == r_count_61_io_out ? io_r_22_b : _GEN_12521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12523 = 8'h17 == r_count_61_io_out ? io_r_23_b : _GEN_12522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12524 = 8'h18 == r_count_61_io_out ? io_r_24_b : _GEN_12523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12525 = 8'h19 == r_count_61_io_out ? io_r_25_b : _GEN_12524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12526 = 8'h1a == r_count_61_io_out ? io_r_26_b : _GEN_12525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12527 = 8'h1b == r_count_61_io_out ? io_r_27_b : _GEN_12526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12528 = 8'h1c == r_count_61_io_out ? io_r_28_b : _GEN_12527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12529 = 8'h1d == r_count_61_io_out ? io_r_29_b : _GEN_12528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12530 = 8'h1e == r_count_61_io_out ? io_r_30_b : _GEN_12529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12531 = 8'h1f == r_count_61_io_out ? io_r_31_b : _GEN_12530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12532 = 8'h20 == r_count_61_io_out ? io_r_32_b : _GEN_12531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12533 = 8'h21 == r_count_61_io_out ? io_r_33_b : _GEN_12532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12534 = 8'h22 == r_count_61_io_out ? io_r_34_b : _GEN_12533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12535 = 8'h23 == r_count_61_io_out ? io_r_35_b : _GEN_12534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12536 = 8'h24 == r_count_61_io_out ? io_r_36_b : _GEN_12535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12537 = 8'h25 == r_count_61_io_out ? io_r_37_b : _GEN_12536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12538 = 8'h26 == r_count_61_io_out ? io_r_38_b : _GEN_12537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12539 = 8'h27 == r_count_61_io_out ? io_r_39_b : _GEN_12538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12540 = 8'h28 == r_count_61_io_out ? io_r_40_b : _GEN_12539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12541 = 8'h29 == r_count_61_io_out ? io_r_41_b : _GEN_12540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12542 = 8'h2a == r_count_61_io_out ? io_r_42_b : _GEN_12541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12543 = 8'h2b == r_count_61_io_out ? io_r_43_b : _GEN_12542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12544 = 8'h2c == r_count_61_io_out ? io_r_44_b : _GEN_12543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12545 = 8'h2d == r_count_61_io_out ? io_r_45_b : _GEN_12544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12546 = 8'h2e == r_count_61_io_out ? io_r_46_b : _GEN_12545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12547 = 8'h2f == r_count_61_io_out ? io_r_47_b : _GEN_12546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12548 = 8'h30 == r_count_61_io_out ? io_r_48_b : _GEN_12547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12549 = 8'h31 == r_count_61_io_out ? io_r_49_b : _GEN_12548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12550 = 8'h32 == r_count_61_io_out ? io_r_50_b : _GEN_12549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12551 = 8'h33 == r_count_61_io_out ? io_r_51_b : _GEN_12550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12552 = 8'h34 == r_count_61_io_out ? io_r_52_b : _GEN_12551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12553 = 8'h35 == r_count_61_io_out ? io_r_53_b : _GEN_12552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12554 = 8'h36 == r_count_61_io_out ? io_r_54_b : _GEN_12553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12555 = 8'h37 == r_count_61_io_out ? io_r_55_b : _GEN_12554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12556 = 8'h38 == r_count_61_io_out ? io_r_56_b : _GEN_12555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12557 = 8'h39 == r_count_61_io_out ? io_r_57_b : _GEN_12556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12558 = 8'h3a == r_count_61_io_out ? io_r_58_b : _GEN_12557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12559 = 8'h3b == r_count_61_io_out ? io_r_59_b : _GEN_12558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12560 = 8'h3c == r_count_61_io_out ? io_r_60_b : _GEN_12559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12561 = 8'h3d == r_count_61_io_out ? io_r_61_b : _GEN_12560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12562 = 8'h3e == r_count_61_io_out ? io_r_62_b : _GEN_12561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12563 = 8'h3f == r_count_61_io_out ? io_r_63_b : _GEN_12562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12564 = 8'h40 == r_count_61_io_out ? io_r_64_b : _GEN_12563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12565 = 8'h41 == r_count_61_io_out ? io_r_65_b : _GEN_12564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12566 = 8'h42 == r_count_61_io_out ? io_r_66_b : _GEN_12565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12567 = 8'h43 == r_count_61_io_out ? io_r_67_b : _GEN_12566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12568 = 8'h44 == r_count_61_io_out ? io_r_68_b : _GEN_12567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12569 = 8'h45 == r_count_61_io_out ? io_r_69_b : _GEN_12568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12570 = 8'h46 == r_count_61_io_out ? io_r_70_b : _GEN_12569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12571 = 8'h47 == r_count_61_io_out ? io_r_71_b : _GEN_12570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12572 = 8'h48 == r_count_61_io_out ? io_r_72_b : _GEN_12571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12573 = 8'h49 == r_count_61_io_out ? io_r_73_b : _GEN_12572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12574 = 8'h4a == r_count_61_io_out ? io_r_74_b : _GEN_12573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12575 = 8'h4b == r_count_61_io_out ? io_r_75_b : _GEN_12574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12576 = 8'h4c == r_count_61_io_out ? io_r_76_b : _GEN_12575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12577 = 8'h4d == r_count_61_io_out ? io_r_77_b : _GEN_12576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12578 = 8'h4e == r_count_61_io_out ? io_r_78_b : _GEN_12577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12579 = 8'h4f == r_count_61_io_out ? io_r_79_b : _GEN_12578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12580 = 8'h50 == r_count_61_io_out ? io_r_80_b : _GEN_12579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12581 = 8'h51 == r_count_61_io_out ? io_r_81_b : _GEN_12580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12582 = 8'h52 == r_count_61_io_out ? io_r_82_b : _GEN_12581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12583 = 8'h53 == r_count_61_io_out ? io_r_83_b : _GEN_12582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12584 = 8'h54 == r_count_61_io_out ? io_r_84_b : _GEN_12583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12585 = 8'h55 == r_count_61_io_out ? io_r_85_b : _GEN_12584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12586 = 8'h56 == r_count_61_io_out ? io_r_86_b : _GEN_12585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12587 = 8'h57 == r_count_61_io_out ? io_r_87_b : _GEN_12586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12588 = 8'h58 == r_count_61_io_out ? io_r_88_b : _GEN_12587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12589 = 8'h59 == r_count_61_io_out ? io_r_89_b : _GEN_12588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12590 = 8'h5a == r_count_61_io_out ? io_r_90_b : _GEN_12589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12591 = 8'h5b == r_count_61_io_out ? io_r_91_b : _GEN_12590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12592 = 8'h5c == r_count_61_io_out ? io_r_92_b : _GEN_12591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12593 = 8'h5d == r_count_61_io_out ? io_r_93_b : _GEN_12592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12594 = 8'h5e == r_count_61_io_out ? io_r_94_b : _GEN_12593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12595 = 8'h5f == r_count_61_io_out ? io_r_95_b : _GEN_12594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12596 = 8'h60 == r_count_61_io_out ? io_r_96_b : _GEN_12595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12597 = 8'h61 == r_count_61_io_out ? io_r_97_b : _GEN_12596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12598 = 8'h62 == r_count_61_io_out ? io_r_98_b : _GEN_12597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12599 = 8'h63 == r_count_61_io_out ? io_r_99_b : _GEN_12598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12600 = 8'h64 == r_count_61_io_out ? io_r_100_b : _GEN_12599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12601 = 8'h65 == r_count_61_io_out ? io_r_101_b : _GEN_12600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12602 = 8'h66 == r_count_61_io_out ? io_r_102_b : _GEN_12601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12603 = 8'h67 == r_count_61_io_out ? io_r_103_b : _GEN_12602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12604 = 8'h68 == r_count_61_io_out ? io_r_104_b : _GEN_12603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12605 = 8'h69 == r_count_61_io_out ? io_r_105_b : _GEN_12604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12606 = 8'h6a == r_count_61_io_out ? io_r_106_b : _GEN_12605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12607 = 8'h6b == r_count_61_io_out ? io_r_107_b : _GEN_12606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12608 = 8'h6c == r_count_61_io_out ? io_r_108_b : _GEN_12607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12609 = 8'h6d == r_count_61_io_out ? io_r_109_b : _GEN_12608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12610 = 8'h6e == r_count_61_io_out ? io_r_110_b : _GEN_12609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12611 = 8'h6f == r_count_61_io_out ? io_r_111_b : _GEN_12610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12612 = 8'h70 == r_count_61_io_out ? io_r_112_b : _GEN_12611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12613 = 8'h71 == r_count_61_io_out ? io_r_113_b : _GEN_12612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12614 = 8'h72 == r_count_61_io_out ? io_r_114_b : _GEN_12613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12615 = 8'h73 == r_count_61_io_out ? io_r_115_b : _GEN_12614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12616 = 8'h74 == r_count_61_io_out ? io_r_116_b : _GEN_12615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12617 = 8'h75 == r_count_61_io_out ? io_r_117_b : _GEN_12616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12618 = 8'h76 == r_count_61_io_out ? io_r_118_b : _GEN_12617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12619 = 8'h77 == r_count_61_io_out ? io_r_119_b : _GEN_12618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12620 = 8'h78 == r_count_61_io_out ? io_r_120_b : _GEN_12619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12621 = 8'h79 == r_count_61_io_out ? io_r_121_b : _GEN_12620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12622 = 8'h7a == r_count_61_io_out ? io_r_122_b : _GEN_12621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12623 = 8'h7b == r_count_61_io_out ? io_r_123_b : _GEN_12622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12624 = 8'h7c == r_count_61_io_out ? io_r_124_b : _GEN_12623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12625 = 8'h7d == r_count_61_io_out ? io_r_125_b : _GEN_12624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12626 = 8'h7e == r_count_61_io_out ? io_r_126_b : _GEN_12625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12627 = 8'h7f == r_count_61_io_out ? io_r_127_b : _GEN_12626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12628 = 8'h80 == r_count_61_io_out ? io_r_128_b : _GEN_12627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12629 = 8'h81 == r_count_61_io_out ? io_r_129_b : _GEN_12628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12630 = 8'h82 == r_count_61_io_out ? io_r_130_b : _GEN_12629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12631 = 8'h83 == r_count_61_io_out ? io_r_131_b : _GEN_12630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12632 = 8'h84 == r_count_61_io_out ? io_r_132_b : _GEN_12631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12633 = 8'h85 == r_count_61_io_out ? io_r_133_b : _GEN_12632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12634 = 8'h86 == r_count_61_io_out ? io_r_134_b : _GEN_12633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12635 = 8'h87 == r_count_61_io_out ? io_r_135_b : _GEN_12634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12636 = 8'h88 == r_count_61_io_out ? io_r_136_b : _GEN_12635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12637 = 8'h89 == r_count_61_io_out ? io_r_137_b : _GEN_12636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12638 = 8'h8a == r_count_61_io_out ? io_r_138_b : _GEN_12637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12639 = 8'h8b == r_count_61_io_out ? io_r_139_b : _GEN_12638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12640 = 8'h8c == r_count_61_io_out ? io_r_140_b : _GEN_12639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12641 = 8'h8d == r_count_61_io_out ? io_r_141_b : _GEN_12640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12642 = 8'h8e == r_count_61_io_out ? io_r_142_b : _GEN_12641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12643 = 8'h8f == r_count_61_io_out ? io_r_143_b : _GEN_12642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12644 = 8'h90 == r_count_61_io_out ? io_r_144_b : _GEN_12643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12645 = 8'h91 == r_count_61_io_out ? io_r_145_b : _GEN_12644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12646 = 8'h92 == r_count_61_io_out ? io_r_146_b : _GEN_12645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12647 = 8'h93 == r_count_61_io_out ? io_r_147_b : _GEN_12646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12648 = 8'h94 == r_count_61_io_out ? io_r_148_b : _GEN_12647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12649 = 8'h95 == r_count_61_io_out ? io_r_149_b : _GEN_12648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12650 = 8'h96 == r_count_61_io_out ? io_r_150_b : _GEN_12649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12651 = 8'h97 == r_count_61_io_out ? io_r_151_b : _GEN_12650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12652 = 8'h98 == r_count_61_io_out ? io_r_152_b : _GEN_12651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12653 = 8'h99 == r_count_61_io_out ? io_r_153_b : _GEN_12652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12654 = 8'h9a == r_count_61_io_out ? io_r_154_b : _GEN_12653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12655 = 8'h9b == r_count_61_io_out ? io_r_155_b : _GEN_12654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12656 = 8'h9c == r_count_61_io_out ? io_r_156_b : _GEN_12655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12657 = 8'h9d == r_count_61_io_out ? io_r_157_b : _GEN_12656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12658 = 8'h9e == r_count_61_io_out ? io_r_158_b : _GEN_12657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12659 = 8'h9f == r_count_61_io_out ? io_r_159_b : _GEN_12658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12660 = 8'ha0 == r_count_61_io_out ? io_r_160_b : _GEN_12659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12661 = 8'ha1 == r_count_61_io_out ? io_r_161_b : _GEN_12660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12662 = 8'ha2 == r_count_61_io_out ? io_r_162_b : _GEN_12661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12663 = 8'ha3 == r_count_61_io_out ? io_r_163_b : _GEN_12662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12664 = 8'ha4 == r_count_61_io_out ? io_r_164_b : _GEN_12663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12665 = 8'ha5 == r_count_61_io_out ? io_r_165_b : _GEN_12664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12666 = 8'ha6 == r_count_61_io_out ? io_r_166_b : _GEN_12665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12667 = 8'ha7 == r_count_61_io_out ? io_r_167_b : _GEN_12666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12668 = 8'ha8 == r_count_61_io_out ? io_r_168_b : _GEN_12667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12669 = 8'ha9 == r_count_61_io_out ? io_r_169_b : _GEN_12668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12670 = 8'haa == r_count_61_io_out ? io_r_170_b : _GEN_12669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12671 = 8'hab == r_count_61_io_out ? io_r_171_b : _GEN_12670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12672 = 8'hac == r_count_61_io_out ? io_r_172_b : _GEN_12671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12673 = 8'had == r_count_61_io_out ? io_r_173_b : _GEN_12672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12674 = 8'hae == r_count_61_io_out ? io_r_174_b : _GEN_12673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12675 = 8'haf == r_count_61_io_out ? io_r_175_b : _GEN_12674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12676 = 8'hb0 == r_count_61_io_out ? io_r_176_b : _GEN_12675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12677 = 8'hb1 == r_count_61_io_out ? io_r_177_b : _GEN_12676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12678 = 8'hb2 == r_count_61_io_out ? io_r_178_b : _GEN_12677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12679 = 8'hb3 == r_count_61_io_out ? io_r_179_b : _GEN_12678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12680 = 8'hb4 == r_count_61_io_out ? io_r_180_b : _GEN_12679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12681 = 8'hb5 == r_count_61_io_out ? io_r_181_b : _GEN_12680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12682 = 8'hb6 == r_count_61_io_out ? io_r_182_b : _GEN_12681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12683 = 8'hb7 == r_count_61_io_out ? io_r_183_b : _GEN_12682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12684 = 8'hb8 == r_count_61_io_out ? io_r_184_b : _GEN_12683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12685 = 8'hb9 == r_count_61_io_out ? io_r_185_b : _GEN_12684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12686 = 8'hba == r_count_61_io_out ? io_r_186_b : _GEN_12685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12687 = 8'hbb == r_count_61_io_out ? io_r_187_b : _GEN_12686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12688 = 8'hbc == r_count_61_io_out ? io_r_188_b : _GEN_12687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12689 = 8'hbd == r_count_61_io_out ? io_r_189_b : _GEN_12688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12690 = 8'hbe == r_count_61_io_out ? io_r_190_b : _GEN_12689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12691 = 8'hbf == r_count_61_io_out ? io_r_191_b : _GEN_12690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12692 = 8'hc0 == r_count_61_io_out ? io_r_192_b : _GEN_12691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12693 = 8'hc1 == r_count_61_io_out ? io_r_193_b : _GEN_12692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12694 = 8'hc2 == r_count_61_io_out ? io_r_194_b : _GEN_12693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12695 = 8'hc3 == r_count_61_io_out ? io_r_195_b : _GEN_12694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12696 = 8'hc4 == r_count_61_io_out ? io_r_196_b : _GEN_12695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12697 = 8'hc5 == r_count_61_io_out ? io_r_197_b : _GEN_12696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12698 = 8'hc6 == r_count_61_io_out ? io_r_198_b : _GEN_12697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12701 = 8'h1 == r_count_62_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12702 = 8'h2 == r_count_62_io_out ? io_r_2_b : _GEN_12701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12703 = 8'h3 == r_count_62_io_out ? io_r_3_b : _GEN_12702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12704 = 8'h4 == r_count_62_io_out ? io_r_4_b : _GEN_12703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12705 = 8'h5 == r_count_62_io_out ? io_r_5_b : _GEN_12704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12706 = 8'h6 == r_count_62_io_out ? io_r_6_b : _GEN_12705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12707 = 8'h7 == r_count_62_io_out ? io_r_7_b : _GEN_12706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12708 = 8'h8 == r_count_62_io_out ? io_r_8_b : _GEN_12707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12709 = 8'h9 == r_count_62_io_out ? io_r_9_b : _GEN_12708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12710 = 8'ha == r_count_62_io_out ? io_r_10_b : _GEN_12709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12711 = 8'hb == r_count_62_io_out ? io_r_11_b : _GEN_12710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12712 = 8'hc == r_count_62_io_out ? io_r_12_b : _GEN_12711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12713 = 8'hd == r_count_62_io_out ? io_r_13_b : _GEN_12712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12714 = 8'he == r_count_62_io_out ? io_r_14_b : _GEN_12713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12715 = 8'hf == r_count_62_io_out ? io_r_15_b : _GEN_12714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12716 = 8'h10 == r_count_62_io_out ? io_r_16_b : _GEN_12715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12717 = 8'h11 == r_count_62_io_out ? io_r_17_b : _GEN_12716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12718 = 8'h12 == r_count_62_io_out ? io_r_18_b : _GEN_12717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12719 = 8'h13 == r_count_62_io_out ? io_r_19_b : _GEN_12718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12720 = 8'h14 == r_count_62_io_out ? io_r_20_b : _GEN_12719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12721 = 8'h15 == r_count_62_io_out ? io_r_21_b : _GEN_12720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12722 = 8'h16 == r_count_62_io_out ? io_r_22_b : _GEN_12721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12723 = 8'h17 == r_count_62_io_out ? io_r_23_b : _GEN_12722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12724 = 8'h18 == r_count_62_io_out ? io_r_24_b : _GEN_12723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12725 = 8'h19 == r_count_62_io_out ? io_r_25_b : _GEN_12724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12726 = 8'h1a == r_count_62_io_out ? io_r_26_b : _GEN_12725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12727 = 8'h1b == r_count_62_io_out ? io_r_27_b : _GEN_12726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12728 = 8'h1c == r_count_62_io_out ? io_r_28_b : _GEN_12727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12729 = 8'h1d == r_count_62_io_out ? io_r_29_b : _GEN_12728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12730 = 8'h1e == r_count_62_io_out ? io_r_30_b : _GEN_12729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12731 = 8'h1f == r_count_62_io_out ? io_r_31_b : _GEN_12730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12732 = 8'h20 == r_count_62_io_out ? io_r_32_b : _GEN_12731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12733 = 8'h21 == r_count_62_io_out ? io_r_33_b : _GEN_12732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12734 = 8'h22 == r_count_62_io_out ? io_r_34_b : _GEN_12733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12735 = 8'h23 == r_count_62_io_out ? io_r_35_b : _GEN_12734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12736 = 8'h24 == r_count_62_io_out ? io_r_36_b : _GEN_12735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12737 = 8'h25 == r_count_62_io_out ? io_r_37_b : _GEN_12736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12738 = 8'h26 == r_count_62_io_out ? io_r_38_b : _GEN_12737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12739 = 8'h27 == r_count_62_io_out ? io_r_39_b : _GEN_12738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12740 = 8'h28 == r_count_62_io_out ? io_r_40_b : _GEN_12739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12741 = 8'h29 == r_count_62_io_out ? io_r_41_b : _GEN_12740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12742 = 8'h2a == r_count_62_io_out ? io_r_42_b : _GEN_12741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12743 = 8'h2b == r_count_62_io_out ? io_r_43_b : _GEN_12742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12744 = 8'h2c == r_count_62_io_out ? io_r_44_b : _GEN_12743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12745 = 8'h2d == r_count_62_io_out ? io_r_45_b : _GEN_12744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12746 = 8'h2e == r_count_62_io_out ? io_r_46_b : _GEN_12745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12747 = 8'h2f == r_count_62_io_out ? io_r_47_b : _GEN_12746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12748 = 8'h30 == r_count_62_io_out ? io_r_48_b : _GEN_12747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12749 = 8'h31 == r_count_62_io_out ? io_r_49_b : _GEN_12748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12750 = 8'h32 == r_count_62_io_out ? io_r_50_b : _GEN_12749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12751 = 8'h33 == r_count_62_io_out ? io_r_51_b : _GEN_12750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12752 = 8'h34 == r_count_62_io_out ? io_r_52_b : _GEN_12751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12753 = 8'h35 == r_count_62_io_out ? io_r_53_b : _GEN_12752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12754 = 8'h36 == r_count_62_io_out ? io_r_54_b : _GEN_12753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12755 = 8'h37 == r_count_62_io_out ? io_r_55_b : _GEN_12754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12756 = 8'h38 == r_count_62_io_out ? io_r_56_b : _GEN_12755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12757 = 8'h39 == r_count_62_io_out ? io_r_57_b : _GEN_12756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12758 = 8'h3a == r_count_62_io_out ? io_r_58_b : _GEN_12757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12759 = 8'h3b == r_count_62_io_out ? io_r_59_b : _GEN_12758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12760 = 8'h3c == r_count_62_io_out ? io_r_60_b : _GEN_12759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12761 = 8'h3d == r_count_62_io_out ? io_r_61_b : _GEN_12760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12762 = 8'h3e == r_count_62_io_out ? io_r_62_b : _GEN_12761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12763 = 8'h3f == r_count_62_io_out ? io_r_63_b : _GEN_12762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12764 = 8'h40 == r_count_62_io_out ? io_r_64_b : _GEN_12763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12765 = 8'h41 == r_count_62_io_out ? io_r_65_b : _GEN_12764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12766 = 8'h42 == r_count_62_io_out ? io_r_66_b : _GEN_12765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12767 = 8'h43 == r_count_62_io_out ? io_r_67_b : _GEN_12766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12768 = 8'h44 == r_count_62_io_out ? io_r_68_b : _GEN_12767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12769 = 8'h45 == r_count_62_io_out ? io_r_69_b : _GEN_12768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12770 = 8'h46 == r_count_62_io_out ? io_r_70_b : _GEN_12769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12771 = 8'h47 == r_count_62_io_out ? io_r_71_b : _GEN_12770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12772 = 8'h48 == r_count_62_io_out ? io_r_72_b : _GEN_12771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12773 = 8'h49 == r_count_62_io_out ? io_r_73_b : _GEN_12772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12774 = 8'h4a == r_count_62_io_out ? io_r_74_b : _GEN_12773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12775 = 8'h4b == r_count_62_io_out ? io_r_75_b : _GEN_12774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12776 = 8'h4c == r_count_62_io_out ? io_r_76_b : _GEN_12775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12777 = 8'h4d == r_count_62_io_out ? io_r_77_b : _GEN_12776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12778 = 8'h4e == r_count_62_io_out ? io_r_78_b : _GEN_12777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12779 = 8'h4f == r_count_62_io_out ? io_r_79_b : _GEN_12778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12780 = 8'h50 == r_count_62_io_out ? io_r_80_b : _GEN_12779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12781 = 8'h51 == r_count_62_io_out ? io_r_81_b : _GEN_12780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12782 = 8'h52 == r_count_62_io_out ? io_r_82_b : _GEN_12781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12783 = 8'h53 == r_count_62_io_out ? io_r_83_b : _GEN_12782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12784 = 8'h54 == r_count_62_io_out ? io_r_84_b : _GEN_12783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12785 = 8'h55 == r_count_62_io_out ? io_r_85_b : _GEN_12784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12786 = 8'h56 == r_count_62_io_out ? io_r_86_b : _GEN_12785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12787 = 8'h57 == r_count_62_io_out ? io_r_87_b : _GEN_12786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12788 = 8'h58 == r_count_62_io_out ? io_r_88_b : _GEN_12787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12789 = 8'h59 == r_count_62_io_out ? io_r_89_b : _GEN_12788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12790 = 8'h5a == r_count_62_io_out ? io_r_90_b : _GEN_12789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12791 = 8'h5b == r_count_62_io_out ? io_r_91_b : _GEN_12790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12792 = 8'h5c == r_count_62_io_out ? io_r_92_b : _GEN_12791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12793 = 8'h5d == r_count_62_io_out ? io_r_93_b : _GEN_12792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12794 = 8'h5e == r_count_62_io_out ? io_r_94_b : _GEN_12793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12795 = 8'h5f == r_count_62_io_out ? io_r_95_b : _GEN_12794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12796 = 8'h60 == r_count_62_io_out ? io_r_96_b : _GEN_12795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12797 = 8'h61 == r_count_62_io_out ? io_r_97_b : _GEN_12796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12798 = 8'h62 == r_count_62_io_out ? io_r_98_b : _GEN_12797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12799 = 8'h63 == r_count_62_io_out ? io_r_99_b : _GEN_12798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12800 = 8'h64 == r_count_62_io_out ? io_r_100_b : _GEN_12799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12801 = 8'h65 == r_count_62_io_out ? io_r_101_b : _GEN_12800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12802 = 8'h66 == r_count_62_io_out ? io_r_102_b : _GEN_12801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12803 = 8'h67 == r_count_62_io_out ? io_r_103_b : _GEN_12802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12804 = 8'h68 == r_count_62_io_out ? io_r_104_b : _GEN_12803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12805 = 8'h69 == r_count_62_io_out ? io_r_105_b : _GEN_12804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12806 = 8'h6a == r_count_62_io_out ? io_r_106_b : _GEN_12805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12807 = 8'h6b == r_count_62_io_out ? io_r_107_b : _GEN_12806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12808 = 8'h6c == r_count_62_io_out ? io_r_108_b : _GEN_12807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12809 = 8'h6d == r_count_62_io_out ? io_r_109_b : _GEN_12808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12810 = 8'h6e == r_count_62_io_out ? io_r_110_b : _GEN_12809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12811 = 8'h6f == r_count_62_io_out ? io_r_111_b : _GEN_12810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12812 = 8'h70 == r_count_62_io_out ? io_r_112_b : _GEN_12811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12813 = 8'h71 == r_count_62_io_out ? io_r_113_b : _GEN_12812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12814 = 8'h72 == r_count_62_io_out ? io_r_114_b : _GEN_12813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12815 = 8'h73 == r_count_62_io_out ? io_r_115_b : _GEN_12814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12816 = 8'h74 == r_count_62_io_out ? io_r_116_b : _GEN_12815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12817 = 8'h75 == r_count_62_io_out ? io_r_117_b : _GEN_12816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12818 = 8'h76 == r_count_62_io_out ? io_r_118_b : _GEN_12817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12819 = 8'h77 == r_count_62_io_out ? io_r_119_b : _GEN_12818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12820 = 8'h78 == r_count_62_io_out ? io_r_120_b : _GEN_12819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12821 = 8'h79 == r_count_62_io_out ? io_r_121_b : _GEN_12820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12822 = 8'h7a == r_count_62_io_out ? io_r_122_b : _GEN_12821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12823 = 8'h7b == r_count_62_io_out ? io_r_123_b : _GEN_12822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12824 = 8'h7c == r_count_62_io_out ? io_r_124_b : _GEN_12823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12825 = 8'h7d == r_count_62_io_out ? io_r_125_b : _GEN_12824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12826 = 8'h7e == r_count_62_io_out ? io_r_126_b : _GEN_12825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12827 = 8'h7f == r_count_62_io_out ? io_r_127_b : _GEN_12826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12828 = 8'h80 == r_count_62_io_out ? io_r_128_b : _GEN_12827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12829 = 8'h81 == r_count_62_io_out ? io_r_129_b : _GEN_12828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12830 = 8'h82 == r_count_62_io_out ? io_r_130_b : _GEN_12829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12831 = 8'h83 == r_count_62_io_out ? io_r_131_b : _GEN_12830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12832 = 8'h84 == r_count_62_io_out ? io_r_132_b : _GEN_12831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12833 = 8'h85 == r_count_62_io_out ? io_r_133_b : _GEN_12832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12834 = 8'h86 == r_count_62_io_out ? io_r_134_b : _GEN_12833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12835 = 8'h87 == r_count_62_io_out ? io_r_135_b : _GEN_12834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12836 = 8'h88 == r_count_62_io_out ? io_r_136_b : _GEN_12835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12837 = 8'h89 == r_count_62_io_out ? io_r_137_b : _GEN_12836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12838 = 8'h8a == r_count_62_io_out ? io_r_138_b : _GEN_12837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12839 = 8'h8b == r_count_62_io_out ? io_r_139_b : _GEN_12838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12840 = 8'h8c == r_count_62_io_out ? io_r_140_b : _GEN_12839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12841 = 8'h8d == r_count_62_io_out ? io_r_141_b : _GEN_12840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12842 = 8'h8e == r_count_62_io_out ? io_r_142_b : _GEN_12841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12843 = 8'h8f == r_count_62_io_out ? io_r_143_b : _GEN_12842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12844 = 8'h90 == r_count_62_io_out ? io_r_144_b : _GEN_12843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12845 = 8'h91 == r_count_62_io_out ? io_r_145_b : _GEN_12844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12846 = 8'h92 == r_count_62_io_out ? io_r_146_b : _GEN_12845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12847 = 8'h93 == r_count_62_io_out ? io_r_147_b : _GEN_12846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12848 = 8'h94 == r_count_62_io_out ? io_r_148_b : _GEN_12847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12849 = 8'h95 == r_count_62_io_out ? io_r_149_b : _GEN_12848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12850 = 8'h96 == r_count_62_io_out ? io_r_150_b : _GEN_12849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12851 = 8'h97 == r_count_62_io_out ? io_r_151_b : _GEN_12850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12852 = 8'h98 == r_count_62_io_out ? io_r_152_b : _GEN_12851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12853 = 8'h99 == r_count_62_io_out ? io_r_153_b : _GEN_12852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12854 = 8'h9a == r_count_62_io_out ? io_r_154_b : _GEN_12853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12855 = 8'h9b == r_count_62_io_out ? io_r_155_b : _GEN_12854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12856 = 8'h9c == r_count_62_io_out ? io_r_156_b : _GEN_12855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12857 = 8'h9d == r_count_62_io_out ? io_r_157_b : _GEN_12856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12858 = 8'h9e == r_count_62_io_out ? io_r_158_b : _GEN_12857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12859 = 8'h9f == r_count_62_io_out ? io_r_159_b : _GEN_12858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12860 = 8'ha0 == r_count_62_io_out ? io_r_160_b : _GEN_12859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12861 = 8'ha1 == r_count_62_io_out ? io_r_161_b : _GEN_12860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12862 = 8'ha2 == r_count_62_io_out ? io_r_162_b : _GEN_12861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12863 = 8'ha3 == r_count_62_io_out ? io_r_163_b : _GEN_12862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12864 = 8'ha4 == r_count_62_io_out ? io_r_164_b : _GEN_12863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12865 = 8'ha5 == r_count_62_io_out ? io_r_165_b : _GEN_12864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12866 = 8'ha6 == r_count_62_io_out ? io_r_166_b : _GEN_12865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12867 = 8'ha7 == r_count_62_io_out ? io_r_167_b : _GEN_12866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12868 = 8'ha8 == r_count_62_io_out ? io_r_168_b : _GEN_12867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12869 = 8'ha9 == r_count_62_io_out ? io_r_169_b : _GEN_12868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12870 = 8'haa == r_count_62_io_out ? io_r_170_b : _GEN_12869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12871 = 8'hab == r_count_62_io_out ? io_r_171_b : _GEN_12870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12872 = 8'hac == r_count_62_io_out ? io_r_172_b : _GEN_12871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12873 = 8'had == r_count_62_io_out ? io_r_173_b : _GEN_12872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12874 = 8'hae == r_count_62_io_out ? io_r_174_b : _GEN_12873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12875 = 8'haf == r_count_62_io_out ? io_r_175_b : _GEN_12874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12876 = 8'hb0 == r_count_62_io_out ? io_r_176_b : _GEN_12875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12877 = 8'hb1 == r_count_62_io_out ? io_r_177_b : _GEN_12876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12878 = 8'hb2 == r_count_62_io_out ? io_r_178_b : _GEN_12877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12879 = 8'hb3 == r_count_62_io_out ? io_r_179_b : _GEN_12878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12880 = 8'hb4 == r_count_62_io_out ? io_r_180_b : _GEN_12879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12881 = 8'hb5 == r_count_62_io_out ? io_r_181_b : _GEN_12880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12882 = 8'hb6 == r_count_62_io_out ? io_r_182_b : _GEN_12881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12883 = 8'hb7 == r_count_62_io_out ? io_r_183_b : _GEN_12882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12884 = 8'hb8 == r_count_62_io_out ? io_r_184_b : _GEN_12883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12885 = 8'hb9 == r_count_62_io_out ? io_r_185_b : _GEN_12884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12886 = 8'hba == r_count_62_io_out ? io_r_186_b : _GEN_12885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12887 = 8'hbb == r_count_62_io_out ? io_r_187_b : _GEN_12886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12888 = 8'hbc == r_count_62_io_out ? io_r_188_b : _GEN_12887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12889 = 8'hbd == r_count_62_io_out ? io_r_189_b : _GEN_12888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12890 = 8'hbe == r_count_62_io_out ? io_r_190_b : _GEN_12889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12891 = 8'hbf == r_count_62_io_out ? io_r_191_b : _GEN_12890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12892 = 8'hc0 == r_count_62_io_out ? io_r_192_b : _GEN_12891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12893 = 8'hc1 == r_count_62_io_out ? io_r_193_b : _GEN_12892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12894 = 8'hc2 == r_count_62_io_out ? io_r_194_b : _GEN_12893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12895 = 8'hc3 == r_count_62_io_out ? io_r_195_b : _GEN_12894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12896 = 8'hc4 == r_count_62_io_out ? io_r_196_b : _GEN_12895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12897 = 8'hc5 == r_count_62_io_out ? io_r_197_b : _GEN_12896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12898 = 8'hc6 == r_count_62_io_out ? io_r_198_b : _GEN_12897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12901 = 8'h1 == r_count_63_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12902 = 8'h2 == r_count_63_io_out ? io_r_2_b : _GEN_12901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12903 = 8'h3 == r_count_63_io_out ? io_r_3_b : _GEN_12902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12904 = 8'h4 == r_count_63_io_out ? io_r_4_b : _GEN_12903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12905 = 8'h5 == r_count_63_io_out ? io_r_5_b : _GEN_12904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12906 = 8'h6 == r_count_63_io_out ? io_r_6_b : _GEN_12905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12907 = 8'h7 == r_count_63_io_out ? io_r_7_b : _GEN_12906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12908 = 8'h8 == r_count_63_io_out ? io_r_8_b : _GEN_12907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12909 = 8'h9 == r_count_63_io_out ? io_r_9_b : _GEN_12908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12910 = 8'ha == r_count_63_io_out ? io_r_10_b : _GEN_12909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12911 = 8'hb == r_count_63_io_out ? io_r_11_b : _GEN_12910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12912 = 8'hc == r_count_63_io_out ? io_r_12_b : _GEN_12911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12913 = 8'hd == r_count_63_io_out ? io_r_13_b : _GEN_12912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12914 = 8'he == r_count_63_io_out ? io_r_14_b : _GEN_12913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12915 = 8'hf == r_count_63_io_out ? io_r_15_b : _GEN_12914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12916 = 8'h10 == r_count_63_io_out ? io_r_16_b : _GEN_12915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12917 = 8'h11 == r_count_63_io_out ? io_r_17_b : _GEN_12916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12918 = 8'h12 == r_count_63_io_out ? io_r_18_b : _GEN_12917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12919 = 8'h13 == r_count_63_io_out ? io_r_19_b : _GEN_12918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12920 = 8'h14 == r_count_63_io_out ? io_r_20_b : _GEN_12919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12921 = 8'h15 == r_count_63_io_out ? io_r_21_b : _GEN_12920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12922 = 8'h16 == r_count_63_io_out ? io_r_22_b : _GEN_12921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12923 = 8'h17 == r_count_63_io_out ? io_r_23_b : _GEN_12922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12924 = 8'h18 == r_count_63_io_out ? io_r_24_b : _GEN_12923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12925 = 8'h19 == r_count_63_io_out ? io_r_25_b : _GEN_12924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12926 = 8'h1a == r_count_63_io_out ? io_r_26_b : _GEN_12925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12927 = 8'h1b == r_count_63_io_out ? io_r_27_b : _GEN_12926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12928 = 8'h1c == r_count_63_io_out ? io_r_28_b : _GEN_12927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12929 = 8'h1d == r_count_63_io_out ? io_r_29_b : _GEN_12928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12930 = 8'h1e == r_count_63_io_out ? io_r_30_b : _GEN_12929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12931 = 8'h1f == r_count_63_io_out ? io_r_31_b : _GEN_12930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12932 = 8'h20 == r_count_63_io_out ? io_r_32_b : _GEN_12931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12933 = 8'h21 == r_count_63_io_out ? io_r_33_b : _GEN_12932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12934 = 8'h22 == r_count_63_io_out ? io_r_34_b : _GEN_12933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12935 = 8'h23 == r_count_63_io_out ? io_r_35_b : _GEN_12934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12936 = 8'h24 == r_count_63_io_out ? io_r_36_b : _GEN_12935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12937 = 8'h25 == r_count_63_io_out ? io_r_37_b : _GEN_12936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12938 = 8'h26 == r_count_63_io_out ? io_r_38_b : _GEN_12937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12939 = 8'h27 == r_count_63_io_out ? io_r_39_b : _GEN_12938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12940 = 8'h28 == r_count_63_io_out ? io_r_40_b : _GEN_12939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12941 = 8'h29 == r_count_63_io_out ? io_r_41_b : _GEN_12940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12942 = 8'h2a == r_count_63_io_out ? io_r_42_b : _GEN_12941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12943 = 8'h2b == r_count_63_io_out ? io_r_43_b : _GEN_12942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12944 = 8'h2c == r_count_63_io_out ? io_r_44_b : _GEN_12943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12945 = 8'h2d == r_count_63_io_out ? io_r_45_b : _GEN_12944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12946 = 8'h2e == r_count_63_io_out ? io_r_46_b : _GEN_12945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12947 = 8'h2f == r_count_63_io_out ? io_r_47_b : _GEN_12946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12948 = 8'h30 == r_count_63_io_out ? io_r_48_b : _GEN_12947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12949 = 8'h31 == r_count_63_io_out ? io_r_49_b : _GEN_12948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12950 = 8'h32 == r_count_63_io_out ? io_r_50_b : _GEN_12949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12951 = 8'h33 == r_count_63_io_out ? io_r_51_b : _GEN_12950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12952 = 8'h34 == r_count_63_io_out ? io_r_52_b : _GEN_12951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12953 = 8'h35 == r_count_63_io_out ? io_r_53_b : _GEN_12952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12954 = 8'h36 == r_count_63_io_out ? io_r_54_b : _GEN_12953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12955 = 8'h37 == r_count_63_io_out ? io_r_55_b : _GEN_12954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12956 = 8'h38 == r_count_63_io_out ? io_r_56_b : _GEN_12955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12957 = 8'h39 == r_count_63_io_out ? io_r_57_b : _GEN_12956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12958 = 8'h3a == r_count_63_io_out ? io_r_58_b : _GEN_12957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12959 = 8'h3b == r_count_63_io_out ? io_r_59_b : _GEN_12958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12960 = 8'h3c == r_count_63_io_out ? io_r_60_b : _GEN_12959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12961 = 8'h3d == r_count_63_io_out ? io_r_61_b : _GEN_12960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12962 = 8'h3e == r_count_63_io_out ? io_r_62_b : _GEN_12961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12963 = 8'h3f == r_count_63_io_out ? io_r_63_b : _GEN_12962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12964 = 8'h40 == r_count_63_io_out ? io_r_64_b : _GEN_12963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12965 = 8'h41 == r_count_63_io_out ? io_r_65_b : _GEN_12964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12966 = 8'h42 == r_count_63_io_out ? io_r_66_b : _GEN_12965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12967 = 8'h43 == r_count_63_io_out ? io_r_67_b : _GEN_12966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12968 = 8'h44 == r_count_63_io_out ? io_r_68_b : _GEN_12967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12969 = 8'h45 == r_count_63_io_out ? io_r_69_b : _GEN_12968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12970 = 8'h46 == r_count_63_io_out ? io_r_70_b : _GEN_12969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12971 = 8'h47 == r_count_63_io_out ? io_r_71_b : _GEN_12970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12972 = 8'h48 == r_count_63_io_out ? io_r_72_b : _GEN_12971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12973 = 8'h49 == r_count_63_io_out ? io_r_73_b : _GEN_12972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12974 = 8'h4a == r_count_63_io_out ? io_r_74_b : _GEN_12973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12975 = 8'h4b == r_count_63_io_out ? io_r_75_b : _GEN_12974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12976 = 8'h4c == r_count_63_io_out ? io_r_76_b : _GEN_12975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12977 = 8'h4d == r_count_63_io_out ? io_r_77_b : _GEN_12976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12978 = 8'h4e == r_count_63_io_out ? io_r_78_b : _GEN_12977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12979 = 8'h4f == r_count_63_io_out ? io_r_79_b : _GEN_12978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12980 = 8'h50 == r_count_63_io_out ? io_r_80_b : _GEN_12979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12981 = 8'h51 == r_count_63_io_out ? io_r_81_b : _GEN_12980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12982 = 8'h52 == r_count_63_io_out ? io_r_82_b : _GEN_12981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12983 = 8'h53 == r_count_63_io_out ? io_r_83_b : _GEN_12982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12984 = 8'h54 == r_count_63_io_out ? io_r_84_b : _GEN_12983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12985 = 8'h55 == r_count_63_io_out ? io_r_85_b : _GEN_12984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12986 = 8'h56 == r_count_63_io_out ? io_r_86_b : _GEN_12985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12987 = 8'h57 == r_count_63_io_out ? io_r_87_b : _GEN_12986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12988 = 8'h58 == r_count_63_io_out ? io_r_88_b : _GEN_12987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12989 = 8'h59 == r_count_63_io_out ? io_r_89_b : _GEN_12988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12990 = 8'h5a == r_count_63_io_out ? io_r_90_b : _GEN_12989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12991 = 8'h5b == r_count_63_io_out ? io_r_91_b : _GEN_12990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12992 = 8'h5c == r_count_63_io_out ? io_r_92_b : _GEN_12991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12993 = 8'h5d == r_count_63_io_out ? io_r_93_b : _GEN_12992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12994 = 8'h5e == r_count_63_io_out ? io_r_94_b : _GEN_12993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12995 = 8'h5f == r_count_63_io_out ? io_r_95_b : _GEN_12994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12996 = 8'h60 == r_count_63_io_out ? io_r_96_b : _GEN_12995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12997 = 8'h61 == r_count_63_io_out ? io_r_97_b : _GEN_12996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12998 = 8'h62 == r_count_63_io_out ? io_r_98_b : _GEN_12997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_12999 = 8'h63 == r_count_63_io_out ? io_r_99_b : _GEN_12998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13000 = 8'h64 == r_count_63_io_out ? io_r_100_b : _GEN_12999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13001 = 8'h65 == r_count_63_io_out ? io_r_101_b : _GEN_13000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13002 = 8'h66 == r_count_63_io_out ? io_r_102_b : _GEN_13001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13003 = 8'h67 == r_count_63_io_out ? io_r_103_b : _GEN_13002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13004 = 8'h68 == r_count_63_io_out ? io_r_104_b : _GEN_13003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13005 = 8'h69 == r_count_63_io_out ? io_r_105_b : _GEN_13004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13006 = 8'h6a == r_count_63_io_out ? io_r_106_b : _GEN_13005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13007 = 8'h6b == r_count_63_io_out ? io_r_107_b : _GEN_13006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13008 = 8'h6c == r_count_63_io_out ? io_r_108_b : _GEN_13007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13009 = 8'h6d == r_count_63_io_out ? io_r_109_b : _GEN_13008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13010 = 8'h6e == r_count_63_io_out ? io_r_110_b : _GEN_13009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13011 = 8'h6f == r_count_63_io_out ? io_r_111_b : _GEN_13010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13012 = 8'h70 == r_count_63_io_out ? io_r_112_b : _GEN_13011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13013 = 8'h71 == r_count_63_io_out ? io_r_113_b : _GEN_13012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13014 = 8'h72 == r_count_63_io_out ? io_r_114_b : _GEN_13013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13015 = 8'h73 == r_count_63_io_out ? io_r_115_b : _GEN_13014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13016 = 8'h74 == r_count_63_io_out ? io_r_116_b : _GEN_13015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13017 = 8'h75 == r_count_63_io_out ? io_r_117_b : _GEN_13016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13018 = 8'h76 == r_count_63_io_out ? io_r_118_b : _GEN_13017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13019 = 8'h77 == r_count_63_io_out ? io_r_119_b : _GEN_13018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13020 = 8'h78 == r_count_63_io_out ? io_r_120_b : _GEN_13019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13021 = 8'h79 == r_count_63_io_out ? io_r_121_b : _GEN_13020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13022 = 8'h7a == r_count_63_io_out ? io_r_122_b : _GEN_13021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13023 = 8'h7b == r_count_63_io_out ? io_r_123_b : _GEN_13022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13024 = 8'h7c == r_count_63_io_out ? io_r_124_b : _GEN_13023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13025 = 8'h7d == r_count_63_io_out ? io_r_125_b : _GEN_13024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13026 = 8'h7e == r_count_63_io_out ? io_r_126_b : _GEN_13025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13027 = 8'h7f == r_count_63_io_out ? io_r_127_b : _GEN_13026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13028 = 8'h80 == r_count_63_io_out ? io_r_128_b : _GEN_13027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13029 = 8'h81 == r_count_63_io_out ? io_r_129_b : _GEN_13028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13030 = 8'h82 == r_count_63_io_out ? io_r_130_b : _GEN_13029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13031 = 8'h83 == r_count_63_io_out ? io_r_131_b : _GEN_13030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13032 = 8'h84 == r_count_63_io_out ? io_r_132_b : _GEN_13031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13033 = 8'h85 == r_count_63_io_out ? io_r_133_b : _GEN_13032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13034 = 8'h86 == r_count_63_io_out ? io_r_134_b : _GEN_13033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13035 = 8'h87 == r_count_63_io_out ? io_r_135_b : _GEN_13034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13036 = 8'h88 == r_count_63_io_out ? io_r_136_b : _GEN_13035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13037 = 8'h89 == r_count_63_io_out ? io_r_137_b : _GEN_13036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13038 = 8'h8a == r_count_63_io_out ? io_r_138_b : _GEN_13037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13039 = 8'h8b == r_count_63_io_out ? io_r_139_b : _GEN_13038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13040 = 8'h8c == r_count_63_io_out ? io_r_140_b : _GEN_13039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13041 = 8'h8d == r_count_63_io_out ? io_r_141_b : _GEN_13040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13042 = 8'h8e == r_count_63_io_out ? io_r_142_b : _GEN_13041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13043 = 8'h8f == r_count_63_io_out ? io_r_143_b : _GEN_13042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13044 = 8'h90 == r_count_63_io_out ? io_r_144_b : _GEN_13043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13045 = 8'h91 == r_count_63_io_out ? io_r_145_b : _GEN_13044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13046 = 8'h92 == r_count_63_io_out ? io_r_146_b : _GEN_13045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13047 = 8'h93 == r_count_63_io_out ? io_r_147_b : _GEN_13046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13048 = 8'h94 == r_count_63_io_out ? io_r_148_b : _GEN_13047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13049 = 8'h95 == r_count_63_io_out ? io_r_149_b : _GEN_13048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13050 = 8'h96 == r_count_63_io_out ? io_r_150_b : _GEN_13049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13051 = 8'h97 == r_count_63_io_out ? io_r_151_b : _GEN_13050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13052 = 8'h98 == r_count_63_io_out ? io_r_152_b : _GEN_13051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13053 = 8'h99 == r_count_63_io_out ? io_r_153_b : _GEN_13052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13054 = 8'h9a == r_count_63_io_out ? io_r_154_b : _GEN_13053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13055 = 8'h9b == r_count_63_io_out ? io_r_155_b : _GEN_13054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13056 = 8'h9c == r_count_63_io_out ? io_r_156_b : _GEN_13055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13057 = 8'h9d == r_count_63_io_out ? io_r_157_b : _GEN_13056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13058 = 8'h9e == r_count_63_io_out ? io_r_158_b : _GEN_13057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13059 = 8'h9f == r_count_63_io_out ? io_r_159_b : _GEN_13058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13060 = 8'ha0 == r_count_63_io_out ? io_r_160_b : _GEN_13059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13061 = 8'ha1 == r_count_63_io_out ? io_r_161_b : _GEN_13060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13062 = 8'ha2 == r_count_63_io_out ? io_r_162_b : _GEN_13061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13063 = 8'ha3 == r_count_63_io_out ? io_r_163_b : _GEN_13062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13064 = 8'ha4 == r_count_63_io_out ? io_r_164_b : _GEN_13063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13065 = 8'ha5 == r_count_63_io_out ? io_r_165_b : _GEN_13064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13066 = 8'ha6 == r_count_63_io_out ? io_r_166_b : _GEN_13065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13067 = 8'ha7 == r_count_63_io_out ? io_r_167_b : _GEN_13066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13068 = 8'ha8 == r_count_63_io_out ? io_r_168_b : _GEN_13067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13069 = 8'ha9 == r_count_63_io_out ? io_r_169_b : _GEN_13068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13070 = 8'haa == r_count_63_io_out ? io_r_170_b : _GEN_13069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13071 = 8'hab == r_count_63_io_out ? io_r_171_b : _GEN_13070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13072 = 8'hac == r_count_63_io_out ? io_r_172_b : _GEN_13071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13073 = 8'had == r_count_63_io_out ? io_r_173_b : _GEN_13072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13074 = 8'hae == r_count_63_io_out ? io_r_174_b : _GEN_13073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13075 = 8'haf == r_count_63_io_out ? io_r_175_b : _GEN_13074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13076 = 8'hb0 == r_count_63_io_out ? io_r_176_b : _GEN_13075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13077 = 8'hb1 == r_count_63_io_out ? io_r_177_b : _GEN_13076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13078 = 8'hb2 == r_count_63_io_out ? io_r_178_b : _GEN_13077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13079 = 8'hb3 == r_count_63_io_out ? io_r_179_b : _GEN_13078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13080 = 8'hb4 == r_count_63_io_out ? io_r_180_b : _GEN_13079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13081 = 8'hb5 == r_count_63_io_out ? io_r_181_b : _GEN_13080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13082 = 8'hb6 == r_count_63_io_out ? io_r_182_b : _GEN_13081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13083 = 8'hb7 == r_count_63_io_out ? io_r_183_b : _GEN_13082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13084 = 8'hb8 == r_count_63_io_out ? io_r_184_b : _GEN_13083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13085 = 8'hb9 == r_count_63_io_out ? io_r_185_b : _GEN_13084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13086 = 8'hba == r_count_63_io_out ? io_r_186_b : _GEN_13085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13087 = 8'hbb == r_count_63_io_out ? io_r_187_b : _GEN_13086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13088 = 8'hbc == r_count_63_io_out ? io_r_188_b : _GEN_13087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13089 = 8'hbd == r_count_63_io_out ? io_r_189_b : _GEN_13088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13090 = 8'hbe == r_count_63_io_out ? io_r_190_b : _GEN_13089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13091 = 8'hbf == r_count_63_io_out ? io_r_191_b : _GEN_13090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13092 = 8'hc0 == r_count_63_io_out ? io_r_192_b : _GEN_13091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13093 = 8'hc1 == r_count_63_io_out ? io_r_193_b : _GEN_13092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13094 = 8'hc2 == r_count_63_io_out ? io_r_194_b : _GEN_13093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13095 = 8'hc3 == r_count_63_io_out ? io_r_195_b : _GEN_13094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13096 = 8'hc4 == r_count_63_io_out ? io_r_196_b : _GEN_13095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13097 = 8'hc5 == r_count_63_io_out ? io_r_197_b : _GEN_13096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13098 = 8'hc6 == r_count_63_io_out ? io_r_198_b : _GEN_13097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13101 = 8'h1 == r_count_64_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13102 = 8'h2 == r_count_64_io_out ? io_r_2_b : _GEN_13101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13103 = 8'h3 == r_count_64_io_out ? io_r_3_b : _GEN_13102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13104 = 8'h4 == r_count_64_io_out ? io_r_4_b : _GEN_13103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13105 = 8'h5 == r_count_64_io_out ? io_r_5_b : _GEN_13104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13106 = 8'h6 == r_count_64_io_out ? io_r_6_b : _GEN_13105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13107 = 8'h7 == r_count_64_io_out ? io_r_7_b : _GEN_13106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13108 = 8'h8 == r_count_64_io_out ? io_r_8_b : _GEN_13107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13109 = 8'h9 == r_count_64_io_out ? io_r_9_b : _GEN_13108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13110 = 8'ha == r_count_64_io_out ? io_r_10_b : _GEN_13109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13111 = 8'hb == r_count_64_io_out ? io_r_11_b : _GEN_13110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13112 = 8'hc == r_count_64_io_out ? io_r_12_b : _GEN_13111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13113 = 8'hd == r_count_64_io_out ? io_r_13_b : _GEN_13112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13114 = 8'he == r_count_64_io_out ? io_r_14_b : _GEN_13113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13115 = 8'hf == r_count_64_io_out ? io_r_15_b : _GEN_13114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13116 = 8'h10 == r_count_64_io_out ? io_r_16_b : _GEN_13115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13117 = 8'h11 == r_count_64_io_out ? io_r_17_b : _GEN_13116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13118 = 8'h12 == r_count_64_io_out ? io_r_18_b : _GEN_13117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13119 = 8'h13 == r_count_64_io_out ? io_r_19_b : _GEN_13118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13120 = 8'h14 == r_count_64_io_out ? io_r_20_b : _GEN_13119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13121 = 8'h15 == r_count_64_io_out ? io_r_21_b : _GEN_13120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13122 = 8'h16 == r_count_64_io_out ? io_r_22_b : _GEN_13121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13123 = 8'h17 == r_count_64_io_out ? io_r_23_b : _GEN_13122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13124 = 8'h18 == r_count_64_io_out ? io_r_24_b : _GEN_13123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13125 = 8'h19 == r_count_64_io_out ? io_r_25_b : _GEN_13124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13126 = 8'h1a == r_count_64_io_out ? io_r_26_b : _GEN_13125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13127 = 8'h1b == r_count_64_io_out ? io_r_27_b : _GEN_13126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13128 = 8'h1c == r_count_64_io_out ? io_r_28_b : _GEN_13127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13129 = 8'h1d == r_count_64_io_out ? io_r_29_b : _GEN_13128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13130 = 8'h1e == r_count_64_io_out ? io_r_30_b : _GEN_13129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13131 = 8'h1f == r_count_64_io_out ? io_r_31_b : _GEN_13130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13132 = 8'h20 == r_count_64_io_out ? io_r_32_b : _GEN_13131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13133 = 8'h21 == r_count_64_io_out ? io_r_33_b : _GEN_13132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13134 = 8'h22 == r_count_64_io_out ? io_r_34_b : _GEN_13133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13135 = 8'h23 == r_count_64_io_out ? io_r_35_b : _GEN_13134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13136 = 8'h24 == r_count_64_io_out ? io_r_36_b : _GEN_13135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13137 = 8'h25 == r_count_64_io_out ? io_r_37_b : _GEN_13136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13138 = 8'h26 == r_count_64_io_out ? io_r_38_b : _GEN_13137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13139 = 8'h27 == r_count_64_io_out ? io_r_39_b : _GEN_13138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13140 = 8'h28 == r_count_64_io_out ? io_r_40_b : _GEN_13139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13141 = 8'h29 == r_count_64_io_out ? io_r_41_b : _GEN_13140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13142 = 8'h2a == r_count_64_io_out ? io_r_42_b : _GEN_13141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13143 = 8'h2b == r_count_64_io_out ? io_r_43_b : _GEN_13142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13144 = 8'h2c == r_count_64_io_out ? io_r_44_b : _GEN_13143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13145 = 8'h2d == r_count_64_io_out ? io_r_45_b : _GEN_13144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13146 = 8'h2e == r_count_64_io_out ? io_r_46_b : _GEN_13145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13147 = 8'h2f == r_count_64_io_out ? io_r_47_b : _GEN_13146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13148 = 8'h30 == r_count_64_io_out ? io_r_48_b : _GEN_13147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13149 = 8'h31 == r_count_64_io_out ? io_r_49_b : _GEN_13148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13150 = 8'h32 == r_count_64_io_out ? io_r_50_b : _GEN_13149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13151 = 8'h33 == r_count_64_io_out ? io_r_51_b : _GEN_13150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13152 = 8'h34 == r_count_64_io_out ? io_r_52_b : _GEN_13151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13153 = 8'h35 == r_count_64_io_out ? io_r_53_b : _GEN_13152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13154 = 8'h36 == r_count_64_io_out ? io_r_54_b : _GEN_13153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13155 = 8'h37 == r_count_64_io_out ? io_r_55_b : _GEN_13154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13156 = 8'h38 == r_count_64_io_out ? io_r_56_b : _GEN_13155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13157 = 8'h39 == r_count_64_io_out ? io_r_57_b : _GEN_13156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13158 = 8'h3a == r_count_64_io_out ? io_r_58_b : _GEN_13157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13159 = 8'h3b == r_count_64_io_out ? io_r_59_b : _GEN_13158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13160 = 8'h3c == r_count_64_io_out ? io_r_60_b : _GEN_13159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13161 = 8'h3d == r_count_64_io_out ? io_r_61_b : _GEN_13160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13162 = 8'h3e == r_count_64_io_out ? io_r_62_b : _GEN_13161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13163 = 8'h3f == r_count_64_io_out ? io_r_63_b : _GEN_13162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13164 = 8'h40 == r_count_64_io_out ? io_r_64_b : _GEN_13163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13165 = 8'h41 == r_count_64_io_out ? io_r_65_b : _GEN_13164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13166 = 8'h42 == r_count_64_io_out ? io_r_66_b : _GEN_13165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13167 = 8'h43 == r_count_64_io_out ? io_r_67_b : _GEN_13166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13168 = 8'h44 == r_count_64_io_out ? io_r_68_b : _GEN_13167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13169 = 8'h45 == r_count_64_io_out ? io_r_69_b : _GEN_13168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13170 = 8'h46 == r_count_64_io_out ? io_r_70_b : _GEN_13169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13171 = 8'h47 == r_count_64_io_out ? io_r_71_b : _GEN_13170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13172 = 8'h48 == r_count_64_io_out ? io_r_72_b : _GEN_13171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13173 = 8'h49 == r_count_64_io_out ? io_r_73_b : _GEN_13172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13174 = 8'h4a == r_count_64_io_out ? io_r_74_b : _GEN_13173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13175 = 8'h4b == r_count_64_io_out ? io_r_75_b : _GEN_13174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13176 = 8'h4c == r_count_64_io_out ? io_r_76_b : _GEN_13175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13177 = 8'h4d == r_count_64_io_out ? io_r_77_b : _GEN_13176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13178 = 8'h4e == r_count_64_io_out ? io_r_78_b : _GEN_13177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13179 = 8'h4f == r_count_64_io_out ? io_r_79_b : _GEN_13178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13180 = 8'h50 == r_count_64_io_out ? io_r_80_b : _GEN_13179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13181 = 8'h51 == r_count_64_io_out ? io_r_81_b : _GEN_13180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13182 = 8'h52 == r_count_64_io_out ? io_r_82_b : _GEN_13181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13183 = 8'h53 == r_count_64_io_out ? io_r_83_b : _GEN_13182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13184 = 8'h54 == r_count_64_io_out ? io_r_84_b : _GEN_13183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13185 = 8'h55 == r_count_64_io_out ? io_r_85_b : _GEN_13184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13186 = 8'h56 == r_count_64_io_out ? io_r_86_b : _GEN_13185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13187 = 8'h57 == r_count_64_io_out ? io_r_87_b : _GEN_13186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13188 = 8'h58 == r_count_64_io_out ? io_r_88_b : _GEN_13187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13189 = 8'h59 == r_count_64_io_out ? io_r_89_b : _GEN_13188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13190 = 8'h5a == r_count_64_io_out ? io_r_90_b : _GEN_13189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13191 = 8'h5b == r_count_64_io_out ? io_r_91_b : _GEN_13190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13192 = 8'h5c == r_count_64_io_out ? io_r_92_b : _GEN_13191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13193 = 8'h5d == r_count_64_io_out ? io_r_93_b : _GEN_13192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13194 = 8'h5e == r_count_64_io_out ? io_r_94_b : _GEN_13193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13195 = 8'h5f == r_count_64_io_out ? io_r_95_b : _GEN_13194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13196 = 8'h60 == r_count_64_io_out ? io_r_96_b : _GEN_13195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13197 = 8'h61 == r_count_64_io_out ? io_r_97_b : _GEN_13196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13198 = 8'h62 == r_count_64_io_out ? io_r_98_b : _GEN_13197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13199 = 8'h63 == r_count_64_io_out ? io_r_99_b : _GEN_13198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13200 = 8'h64 == r_count_64_io_out ? io_r_100_b : _GEN_13199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13201 = 8'h65 == r_count_64_io_out ? io_r_101_b : _GEN_13200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13202 = 8'h66 == r_count_64_io_out ? io_r_102_b : _GEN_13201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13203 = 8'h67 == r_count_64_io_out ? io_r_103_b : _GEN_13202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13204 = 8'h68 == r_count_64_io_out ? io_r_104_b : _GEN_13203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13205 = 8'h69 == r_count_64_io_out ? io_r_105_b : _GEN_13204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13206 = 8'h6a == r_count_64_io_out ? io_r_106_b : _GEN_13205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13207 = 8'h6b == r_count_64_io_out ? io_r_107_b : _GEN_13206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13208 = 8'h6c == r_count_64_io_out ? io_r_108_b : _GEN_13207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13209 = 8'h6d == r_count_64_io_out ? io_r_109_b : _GEN_13208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13210 = 8'h6e == r_count_64_io_out ? io_r_110_b : _GEN_13209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13211 = 8'h6f == r_count_64_io_out ? io_r_111_b : _GEN_13210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13212 = 8'h70 == r_count_64_io_out ? io_r_112_b : _GEN_13211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13213 = 8'h71 == r_count_64_io_out ? io_r_113_b : _GEN_13212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13214 = 8'h72 == r_count_64_io_out ? io_r_114_b : _GEN_13213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13215 = 8'h73 == r_count_64_io_out ? io_r_115_b : _GEN_13214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13216 = 8'h74 == r_count_64_io_out ? io_r_116_b : _GEN_13215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13217 = 8'h75 == r_count_64_io_out ? io_r_117_b : _GEN_13216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13218 = 8'h76 == r_count_64_io_out ? io_r_118_b : _GEN_13217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13219 = 8'h77 == r_count_64_io_out ? io_r_119_b : _GEN_13218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13220 = 8'h78 == r_count_64_io_out ? io_r_120_b : _GEN_13219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13221 = 8'h79 == r_count_64_io_out ? io_r_121_b : _GEN_13220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13222 = 8'h7a == r_count_64_io_out ? io_r_122_b : _GEN_13221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13223 = 8'h7b == r_count_64_io_out ? io_r_123_b : _GEN_13222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13224 = 8'h7c == r_count_64_io_out ? io_r_124_b : _GEN_13223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13225 = 8'h7d == r_count_64_io_out ? io_r_125_b : _GEN_13224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13226 = 8'h7e == r_count_64_io_out ? io_r_126_b : _GEN_13225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13227 = 8'h7f == r_count_64_io_out ? io_r_127_b : _GEN_13226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13228 = 8'h80 == r_count_64_io_out ? io_r_128_b : _GEN_13227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13229 = 8'h81 == r_count_64_io_out ? io_r_129_b : _GEN_13228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13230 = 8'h82 == r_count_64_io_out ? io_r_130_b : _GEN_13229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13231 = 8'h83 == r_count_64_io_out ? io_r_131_b : _GEN_13230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13232 = 8'h84 == r_count_64_io_out ? io_r_132_b : _GEN_13231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13233 = 8'h85 == r_count_64_io_out ? io_r_133_b : _GEN_13232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13234 = 8'h86 == r_count_64_io_out ? io_r_134_b : _GEN_13233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13235 = 8'h87 == r_count_64_io_out ? io_r_135_b : _GEN_13234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13236 = 8'h88 == r_count_64_io_out ? io_r_136_b : _GEN_13235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13237 = 8'h89 == r_count_64_io_out ? io_r_137_b : _GEN_13236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13238 = 8'h8a == r_count_64_io_out ? io_r_138_b : _GEN_13237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13239 = 8'h8b == r_count_64_io_out ? io_r_139_b : _GEN_13238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13240 = 8'h8c == r_count_64_io_out ? io_r_140_b : _GEN_13239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13241 = 8'h8d == r_count_64_io_out ? io_r_141_b : _GEN_13240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13242 = 8'h8e == r_count_64_io_out ? io_r_142_b : _GEN_13241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13243 = 8'h8f == r_count_64_io_out ? io_r_143_b : _GEN_13242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13244 = 8'h90 == r_count_64_io_out ? io_r_144_b : _GEN_13243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13245 = 8'h91 == r_count_64_io_out ? io_r_145_b : _GEN_13244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13246 = 8'h92 == r_count_64_io_out ? io_r_146_b : _GEN_13245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13247 = 8'h93 == r_count_64_io_out ? io_r_147_b : _GEN_13246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13248 = 8'h94 == r_count_64_io_out ? io_r_148_b : _GEN_13247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13249 = 8'h95 == r_count_64_io_out ? io_r_149_b : _GEN_13248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13250 = 8'h96 == r_count_64_io_out ? io_r_150_b : _GEN_13249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13251 = 8'h97 == r_count_64_io_out ? io_r_151_b : _GEN_13250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13252 = 8'h98 == r_count_64_io_out ? io_r_152_b : _GEN_13251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13253 = 8'h99 == r_count_64_io_out ? io_r_153_b : _GEN_13252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13254 = 8'h9a == r_count_64_io_out ? io_r_154_b : _GEN_13253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13255 = 8'h9b == r_count_64_io_out ? io_r_155_b : _GEN_13254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13256 = 8'h9c == r_count_64_io_out ? io_r_156_b : _GEN_13255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13257 = 8'h9d == r_count_64_io_out ? io_r_157_b : _GEN_13256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13258 = 8'h9e == r_count_64_io_out ? io_r_158_b : _GEN_13257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13259 = 8'h9f == r_count_64_io_out ? io_r_159_b : _GEN_13258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13260 = 8'ha0 == r_count_64_io_out ? io_r_160_b : _GEN_13259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13261 = 8'ha1 == r_count_64_io_out ? io_r_161_b : _GEN_13260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13262 = 8'ha2 == r_count_64_io_out ? io_r_162_b : _GEN_13261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13263 = 8'ha3 == r_count_64_io_out ? io_r_163_b : _GEN_13262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13264 = 8'ha4 == r_count_64_io_out ? io_r_164_b : _GEN_13263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13265 = 8'ha5 == r_count_64_io_out ? io_r_165_b : _GEN_13264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13266 = 8'ha6 == r_count_64_io_out ? io_r_166_b : _GEN_13265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13267 = 8'ha7 == r_count_64_io_out ? io_r_167_b : _GEN_13266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13268 = 8'ha8 == r_count_64_io_out ? io_r_168_b : _GEN_13267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13269 = 8'ha9 == r_count_64_io_out ? io_r_169_b : _GEN_13268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13270 = 8'haa == r_count_64_io_out ? io_r_170_b : _GEN_13269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13271 = 8'hab == r_count_64_io_out ? io_r_171_b : _GEN_13270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13272 = 8'hac == r_count_64_io_out ? io_r_172_b : _GEN_13271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13273 = 8'had == r_count_64_io_out ? io_r_173_b : _GEN_13272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13274 = 8'hae == r_count_64_io_out ? io_r_174_b : _GEN_13273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13275 = 8'haf == r_count_64_io_out ? io_r_175_b : _GEN_13274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13276 = 8'hb0 == r_count_64_io_out ? io_r_176_b : _GEN_13275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13277 = 8'hb1 == r_count_64_io_out ? io_r_177_b : _GEN_13276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13278 = 8'hb2 == r_count_64_io_out ? io_r_178_b : _GEN_13277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13279 = 8'hb3 == r_count_64_io_out ? io_r_179_b : _GEN_13278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13280 = 8'hb4 == r_count_64_io_out ? io_r_180_b : _GEN_13279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13281 = 8'hb5 == r_count_64_io_out ? io_r_181_b : _GEN_13280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13282 = 8'hb6 == r_count_64_io_out ? io_r_182_b : _GEN_13281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13283 = 8'hb7 == r_count_64_io_out ? io_r_183_b : _GEN_13282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13284 = 8'hb8 == r_count_64_io_out ? io_r_184_b : _GEN_13283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13285 = 8'hb9 == r_count_64_io_out ? io_r_185_b : _GEN_13284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13286 = 8'hba == r_count_64_io_out ? io_r_186_b : _GEN_13285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13287 = 8'hbb == r_count_64_io_out ? io_r_187_b : _GEN_13286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13288 = 8'hbc == r_count_64_io_out ? io_r_188_b : _GEN_13287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13289 = 8'hbd == r_count_64_io_out ? io_r_189_b : _GEN_13288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13290 = 8'hbe == r_count_64_io_out ? io_r_190_b : _GEN_13289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13291 = 8'hbf == r_count_64_io_out ? io_r_191_b : _GEN_13290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13292 = 8'hc0 == r_count_64_io_out ? io_r_192_b : _GEN_13291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13293 = 8'hc1 == r_count_64_io_out ? io_r_193_b : _GEN_13292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13294 = 8'hc2 == r_count_64_io_out ? io_r_194_b : _GEN_13293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13295 = 8'hc3 == r_count_64_io_out ? io_r_195_b : _GEN_13294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13296 = 8'hc4 == r_count_64_io_out ? io_r_196_b : _GEN_13295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13297 = 8'hc5 == r_count_64_io_out ? io_r_197_b : _GEN_13296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13298 = 8'hc6 == r_count_64_io_out ? io_r_198_b : _GEN_13297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13301 = 8'h1 == r_count_65_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13302 = 8'h2 == r_count_65_io_out ? io_r_2_b : _GEN_13301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13303 = 8'h3 == r_count_65_io_out ? io_r_3_b : _GEN_13302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13304 = 8'h4 == r_count_65_io_out ? io_r_4_b : _GEN_13303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13305 = 8'h5 == r_count_65_io_out ? io_r_5_b : _GEN_13304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13306 = 8'h6 == r_count_65_io_out ? io_r_6_b : _GEN_13305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13307 = 8'h7 == r_count_65_io_out ? io_r_7_b : _GEN_13306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13308 = 8'h8 == r_count_65_io_out ? io_r_8_b : _GEN_13307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13309 = 8'h9 == r_count_65_io_out ? io_r_9_b : _GEN_13308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13310 = 8'ha == r_count_65_io_out ? io_r_10_b : _GEN_13309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13311 = 8'hb == r_count_65_io_out ? io_r_11_b : _GEN_13310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13312 = 8'hc == r_count_65_io_out ? io_r_12_b : _GEN_13311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13313 = 8'hd == r_count_65_io_out ? io_r_13_b : _GEN_13312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13314 = 8'he == r_count_65_io_out ? io_r_14_b : _GEN_13313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13315 = 8'hf == r_count_65_io_out ? io_r_15_b : _GEN_13314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13316 = 8'h10 == r_count_65_io_out ? io_r_16_b : _GEN_13315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13317 = 8'h11 == r_count_65_io_out ? io_r_17_b : _GEN_13316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13318 = 8'h12 == r_count_65_io_out ? io_r_18_b : _GEN_13317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13319 = 8'h13 == r_count_65_io_out ? io_r_19_b : _GEN_13318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13320 = 8'h14 == r_count_65_io_out ? io_r_20_b : _GEN_13319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13321 = 8'h15 == r_count_65_io_out ? io_r_21_b : _GEN_13320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13322 = 8'h16 == r_count_65_io_out ? io_r_22_b : _GEN_13321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13323 = 8'h17 == r_count_65_io_out ? io_r_23_b : _GEN_13322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13324 = 8'h18 == r_count_65_io_out ? io_r_24_b : _GEN_13323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13325 = 8'h19 == r_count_65_io_out ? io_r_25_b : _GEN_13324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13326 = 8'h1a == r_count_65_io_out ? io_r_26_b : _GEN_13325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13327 = 8'h1b == r_count_65_io_out ? io_r_27_b : _GEN_13326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13328 = 8'h1c == r_count_65_io_out ? io_r_28_b : _GEN_13327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13329 = 8'h1d == r_count_65_io_out ? io_r_29_b : _GEN_13328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13330 = 8'h1e == r_count_65_io_out ? io_r_30_b : _GEN_13329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13331 = 8'h1f == r_count_65_io_out ? io_r_31_b : _GEN_13330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13332 = 8'h20 == r_count_65_io_out ? io_r_32_b : _GEN_13331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13333 = 8'h21 == r_count_65_io_out ? io_r_33_b : _GEN_13332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13334 = 8'h22 == r_count_65_io_out ? io_r_34_b : _GEN_13333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13335 = 8'h23 == r_count_65_io_out ? io_r_35_b : _GEN_13334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13336 = 8'h24 == r_count_65_io_out ? io_r_36_b : _GEN_13335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13337 = 8'h25 == r_count_65_io_out ? io_r_37_b : _GEN_13336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13338 = 8'h26 == r_count_65_io_out ? io_r_38_b : _GEN_13337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13339 = 8'h27 == r_count_65_io_out ? io_r_39_b : _GEN_13338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13340 = 8'h28 == r_count_65_io_out ? io_r_40_b : _GEN_13339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13341 = 8'h29 == r_count_65_io_out ? io_r_41_b : _GEN_13340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13342 = 8'h2a == r_count_65_io_out ? io_r_42_b : _GEN_13341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13343 = 8'h2b == r_count_65_io_out ? io_r_43_b : _GEN_13342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13344 = 8'h2c == r_count_65_io_out ? io_r_44_b : _GEN_13343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13345 = 8'h2d == r_count_65_io_out ? io_r_45_b : _GEN_13344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13346 = 8'h2e == r_count_65_io_out ? io_r_46_b : _GEN_13345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13347 = 8'h2f == r_count_65_io_out ? io_r_47_b : _GEN_13346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13348 = 8'h30 == r_count_65_io_out ? io_r_48_b : _GEN_13347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13349 = 8'h31 == r_count_65_io_out ? io_r_49_b : _GEN_13348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13350 = 8'h32 == r_count_65_io_out ? io_r_50_b : _GEN_13349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13351 = 8'h33 == r_count_65_io_out ? io_r_51_b : _GEN_13350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13352 = 8'h34 == r_count_65_io_out ? io_r_52_b : _GEN_13351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13353 = 8'h35 == r_count_65_io_out ? io_r_53_b : _GEN_13352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13354 = 8'h36 == r_count_65_io_out ? io_r_54_b : _GEN_13353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13355 = 8'h37 == r_count_65_io_out ? io_r_55_b : _GEN_13354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13356 = 8'h38 == r_count_65_io_out ? io_r_56_b : _GEN_13355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13357 = 8'h39 == r_count_65_io_out ? io_r_57_b : _GEN_13356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13358 = 8'h3a == r_count_65_io_out ? io_r_58_b : _GEN_13357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13359 = 8'h3b == r_count_65_io_out ? io_r_59_b : _GEN_13358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13360 = 8'h3c == r_count_65_io_out ? io_r_60_b : _GEN_13359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13361 = 8'h3d == r_count_65_io_out ? io_r_61_b : _GEN_13360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13362 = 8'h3e == r_count_65_io_out ? io_r_62_b : _GEN_13361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13363 = 8'h3f == r_count_65_io_out ? io_r_63_b : _GEN_13362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13364 = 8'h40 == r_count_65_io_out ? io_r_64_b : _GEN_13363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13365 = 8'h41 == r_count_65_io_out ? io_r_65_b : _GEN_13364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13366 = 8'h42 == r_count_65_io_out ? io_r_66_b : _GEN_13365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13367 = 8'h43 == r_count_65_io_out ? io_r_67_b : _GEN_13366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13368 = 8'h44 == r_count_65_io_out ? io_r_68_b : _GEN_13367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13369 = 8'h45 == r_count_65_io_out ? io_r_69_b : _GEN_13368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13370 = 8'h46 == r_count_65_io_out ? io_r_70_b : _GEN_13369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13371 = 8'h47 == r_count_65_io_out ? io_r_71_b : _GEN_13370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13372 = 8'h48 == r_count_65_io_out ? io_r_72_b : _GEN_13371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13373 = 8'h49 == r_count_65_io_out ? io_r_73_b : _GEN_13372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13374 = 8'h4a == r_count_65_io_out ? io_r_74_b : _GEN_13373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13375 = 8'h4b == r_count_65_io_out ? io_r_75_b : _GEN_13374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13376 = 8'h4c == r_count_65_io_out ? io_r_76_b : _GEN_13375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13377 = 8'h4d == r_count_65_io_out ? io_r_77_b : _GEN_13376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13378 = 8'h4e == r_count_65_io_out ? io_r_78_b : _GEN_13377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13379 = 8'h4f == r_count_65_io_out ? io_r_79_b : _GEN_13378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13380 = 8'h50 == r_count_65_io_out ? io_r_80_b : _GEN_13379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13381 = 8'h51 == r_count_65_io_out ? io_r_81_b : _GEN_13380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13382 = 8'h52 == r_count_65_io_out ? io_r_82_b : _GEN_13381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13383 = 8'h53 == r_count_65_io_out ? io_r_83_b : _GEN_13382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13384 = 8'h54 == r_count_65_io_out ? io_r_84_b : _GEN_13383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13385 = 8'h55 == r_count_65_io_out ? io_r_85_b : _GEN_13384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13386 = 8'h56 == r_count_65_io_out ? io_r_86_b : _GEN_13385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13387 = 8'h57 == r_count_65_io_out ? io_r_87_b : _GEN_13386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13388 = 8'h58 == r_count_65_io_out ? io_r_88_b : _GEN_13387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13389 = 8'h59 == r_count_65_io_out ? io_r_89_b : _GEN_13388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13390 = 8'h5a == r_count_65_io_out ? io_r_90_b : _GEN_13389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13391 = 8'h5b == r_count_65_io_out ? io_r_91_b : _GEN_13390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13392 = 8'h5c == r_count_65_io_out ? io_r_92_b : _GEN_13391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13393 = 8'h5d == r_count_65_io_out ? io_r_93_b : _GEN_13392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13394 = 8'h5e == r_count_65_io_out ? io_r_94_b : _GEN_13393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13395 = 8'h5f == r_count_65_io_out ? io_r_95_b : _GEN_13394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13396 = 8'h60 == r_count_65_io_out ? io_r_96_b : _GEN_13395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13397 = 8'h61 == r_count_65_io_out ? io_r_97_b : _GEN_13396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13398 = 8'h62 == r_count_65_io_out ? io_r_98_b : _GEN_13397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13399 = 8'h63 == r_count_65_io_out ? io_r_99_b : _GEN_13398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13400 = 8'h64 == r_count_65_io_out ? io_r_100_b : _GEN_13399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13401 = 8'h65 == r_count_65_io_out ? io_r_101_b : _GEN_13400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13402 = 8'h66 == r_count_65_io_out ? io_r_102_b : _GEN_13401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13403 = 8'h67 == r_count_65_io_out ? io_r_103_b : _GEN_13402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13404 = 8'h68 == r_count_65_io_out ? io_r_104_b : _GEN_13403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13405 = 8'h69 == r_count_65_io_out ? io_r_105_b : _GEN_13404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13406 = 8'h6a == r_count_65_io_out ? io_r_106_b : _GEN_13405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13407 = 8'h6b == r_count_65_io_out ? io_r_107_b : _GEN_13406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13408 = 8'h6c == r_count_65_io_out ? io_r_108_b : _GEN_13407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13409 = 8'h6d == r_count_65_io_out ? io_r_109_b : _GEN_13408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13410 = 8'h6e == r_count_65_io_out ? io_r_110_b : _GEN_13409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13411 = 8'h6f == r_count_65_io_out ? io_r_111_b : _GEN_13410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13412 = 8'h70 == r_count_65_io_out ? io_r_112_b : _GEN_13411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13413 = 8'h71 == r_count_65_io_out ? io_r_113_b : _GEN_13412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13414 = 8'h72 == r_count_65_io_out ? io_r_114_b : _GEN_13413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13415 = 8'h73 == r_count_65_io_out ? io_r_115_b : _GEN_13414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13416 = 8'h74 == r_count_65_io_out ? io_r_116_b : _GEN_13415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13417 = 8'h75 == r_count_65_io_out ? io_r_117_b : _GEN_13416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13418 = 8'h76 == r_count_65_io_out ? io_r_118_b : _GEN_13417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13419 = 8'h77 == r_count_65_io_out ? io_r_119_b : _GEN_13418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13420 = 8'h78 == r_count_65_io_out ? io_r_120_b : _GEN_13419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13421 = 8'h79 == r_count_65_io_out ? io_r_121_b : _GEN_13420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13422 = 8'h7a == r_count_65_io_out ? io_r_122_b : _GEN_13421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13423 = 8'h7b == r_count_65_io_out ? io_r_123_b : _GEN_13422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13424 = 8'h7c == r_count_65_io_out ? io_r_124_b : _GEN_13423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13425 = 8'h7d == r_count_65_io_out ? io_r_125_b : _GEN_13424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13426 = 8'h7e == r_count_65_io_out ? io_r_126_b : _GEN_13425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13427 = 8'h7f == r_count_65_io_out ? io_r_127_b : _GEN_13426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13428 = 8'h80 == r_count_65_io_out ? io_r_128_b : _GEN_13427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13429 = 8'h81 == r_count_65_io_out ? io_r_129_b : _GEN_13428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13430 = 8'h82 == r_count_65_io_out ? io_r_130_b : _GEN_13429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13431 = 8'h83 == r_count_65_io_out ? io_r_131_b : _GEN_13430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13432 = 8'h84 == r_count_65_io_out ? io_r_132_b : _GEN_13431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13433 = 8'h85 == r_count_65_io_out ? io_r_133_b : _GEN_13432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13434 = 8'h86 == r_count_65_io_out ? io_r_134_b : _GEN_13433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13435 = 8'h87 == r_count_65_io_out ? io_r_135_b : _GEN_13434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13436 = 8'h88 == r_count_65_io_out ? io_r_136_b : _GEN_13435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13437 = 8'h89 == r_count_65_io_out ? io_r_137_b : _GEN_13436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13438 = 8'h8a == r_count_65_io_out ? io_r_138_b : _GEN_13437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13439 = 8'h8b == r_count_65_io_out ? io_r_139_b : _GEN_13438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13440 = 8'h8c == r_count_65_io_out ? io_r_140_b : _GEN_13439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13441 = 8'h8d == r_count_65_io_out ? io_r_141_b : _GEN_13440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13442 = 8'h8e == r_count_65_io_out ? io_r_142_b : _GEN_13441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13443 = 8'h8f == r_count_65_io_out ? io_r_143_b : _GEN_13442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13444 = 8'h90 == r_count_65_io_out ? io_r_144_b : _GEN_13443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13445 = 8'h91 == r_count_65_io_out ? io_r_145_b : _GEN_13444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13446 = 8'h92 == r_count_65_io_out ? io_r_146_b : _GEN_13445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13447 = 8'h93 == r_count_65_io_out ? io_r_147_b : _GEN_13446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13448 = 8'h94 == r_count_65_io_out ? io_r_148_b : _GEN_13447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13449 = 8'h95 == r_count_65_io_out ? io_r_149_b : _GEN_13448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13450 = 8'h96 == r_count_65_io_out ? io_r_150_b : _GEN_13449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13451 = 8'h97 == r_count_65_io_out ? io_r_151_b : _GEN_13450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13452 = 8'h98 == r_count_65_io_out ? io_r_152_b : _GEN_13451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13453 = 8'h99 == r_count_65_io_out ? io_r_153_b : _GEN_13452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13454 = 8'h9a == r_count_65_io_out ? io_r_154_b : _GEN_13453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13455 = 8'h9b == r_count_65_io_out ? io_r_155_b : _GEN_13454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13456 = 8'h9c == r_count_65_io_out ? io_r_156_b : _GEN_13455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13457 = 8'h9d == r_count_65_io_out ? io_r_157_b : _GEN_13456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13458 = 8'h9e == r_count_65_io_out ? io_r_158_b : _GEN_13457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13459 = 8'h9f == r_count_65_io_out ? io_r_159_b : _GEN_13458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13460 = 8'ha0 == r_count_65_io_out ? io_r_160_b : _GEN_13459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13461 = 8'ha1 == r_count_65_io_out ? io_r_161_b : _GEN_13460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13462 = 8'ha2 == r_count_65_io_out ? io_r_162_b : _GEN_13461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13463 = 8'ha3 == r_count_65_io_out ? io_r_163_b : _GEN_13462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13464 = 8'ha4 == r_count_65_io_out ? io_r_164_b : _GEN_13463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13465 = 8'ha5 == r_count_65_io_out ? io_r_165_b : _GEN_13464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13466 = 8'ha6 == r_count_65_io_out ? io_r_166_b : _GEN_13465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13467 = 8'ha7 == r_count_65_io_out ? io_r_167_b : _GEN_13466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13468 = 8'ha8 == r_count_65_io_out ? io_r_168_b : _GEN_13467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13469 = 8'ha9 == r_count_65_io_out ? io_r_169_b : _GEN_13468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13470 = 8'haa == r_count_65_io_out ? io_r_170_b : _GEN_13469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13471 = 8'hab == r_count_65_io_out ? io_r_171_b : _GEN_13470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13472 = 8'hac == r_count_65_io_out ? io_r_172_b : _GEN_13471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13473 = 8'had == r_count_65_io_out ? io_r_173_b : _GEN_13472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13474 = 8'hae == r_count_65_io_out ? io_r_174_b : _GEN_13473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13475 = 8'haf == r_count_65_io_out ? io_r_175_b : _GEN_13474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13476 = 8'hb0 == r_count_65_io_out ? io_r_176_b : _GEN_13475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13477 = 8'hb1 == r_count_65_io_out ? io_r_177_b : _GEN_13476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13478 = 8'hb2 == r_count_65_io_out ? io_r_178_b : _GEN_13477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13479 = 8'hb3 == r_count_65_io_out ? io_r_179_b : _GEN_13478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13480 = 8'hb4 == r_count_65_io_out ? io_r_180_b : _GEN_13479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13481 = 8'hb5 == r_count_65_io_out ? io_r_181_b : _GEN_13480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13482 = 8'hb6 == r_count_65_io_out ? io_r_182_b : _GEN_13481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13483 = 8'hb7 == r_count_65_io_out ? io_r_183_b : _GEN_13482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13484 = 8'hb8 == r_count_65_io_out ? io_r_184_b : _GEN_13483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13485 = 8'hb9 == r_count_65_io_out ? io_r_185_b : _GEN_13484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13486 = 8'hba == r_count_65_io_out ? io_r_186_b : _GEN_13485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13487 = 8'hbb == r_count_65_io_out ? io_r_187_b : _GEN_13486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13488 = 8'hbc == r_count_65_io_out ? io_r_188_b : _GEN_13487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13489 = 8'hbd == r_count_65_io_out ? io_r_189_b : _GEN_13488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13490 = 8'hbe == r_count_65_io_out ? io_r_190_b : _GEN_13489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13491 = 8'hbf == r_count_65_io_out ? io_r_191_b : _GEN_13490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13492 = 8'hc0 == r_count_65_io_out ? io_r_192_b : _GEN_13491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13493 = 8'hc1 == r_count_65_io_out ? io_r_193_b : _GEN_13492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13494 = 8'hc2 == r_count_65_io_out ? io_r_194_b : _GEN_13493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13495 = 8'hc3 == r_count_65_io_out ? io_r_195_b : _GEN_13494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13496 = 8'hc4 == r_count_65_io_out ? io_r_196_b : _GEN_13495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13497 = 8'hc5 == r_count_65_io_out ? io_r_197_b : _GEN_13496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13498 = 8'hc6 == r_count_65_io_out ? io_r_198_b : _GEN_13497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13501 = 8'h1 == r_count_66_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13502 = 8'h2 == r_count_66_io_out ? io_r_2_b : _GEN_13501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13503 = 8'h3 == r_count_66_io_out ? io_r_3_b : _GEN_13502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13504 = 8'h4 == r_count_66_io_out ? io_r_4_b : _GEN_13503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13505 = 8'h5 == r_count_66_io_out ? io_r_5_b : _GEN_13504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13506 = 8'h6 == r_count_66_io_out ? io_r_6_b : _GEN_13505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13507 = 8'h7 == r_count_66_io_out ? io_r_7_b : _GEN_13506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13508 = 8'h8 == r_count_66_io_out ? io_r_8_b : _GEN_13507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13509 = 8'h9 == r_count_66_io_out ? io_r_9_b : _GEN_13508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13510 = 8'ha == r_count_66_io_out ? io_r_10_b : _GEN_13509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13511 = 8'hb == r_count_66_io_out ? io_r_11_b : _GEN_13510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13512 = 8'hc == r_count_66_io_out ? io_r_12_b : _GEN_13511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13513 = 8'hd == r_count_66_io_out ? io_r_13_b : _GEN_13512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13514 = 8'he == r_count_66_io_out ? io_r_14_b : _GEN_13513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13515 = 8'hf == r_count_66_io_out ? io_r_15_b : _GEN_13514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13516 = 8'h10 == r_count_66_io_out ? io_r_16_b : _GEN_13515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13517 = 8'h11 == r_count_66_io_out ? io_r_17_b : _GEN_13516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13518 = 8'h12 == r_count_66_io_out ? io_r_18_b : _GEN_13517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13519 = 8'h13 == r_count_66_io_out ? io_r_19_b : _GEN_13518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13520 = 8'h14 == r_count_66_io_out ? io_r_20_b : _GEN_13519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13521 = 8'h15 == r_count_66_io_out ? io_r_21_b : _GEN_13520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13522 = 8'h16 == r_count_66_io_out ? io_r_22_b : _GEN_13521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13523 = 8'h17 == r_count_66_io_out ? io_r_23_b : _GEN_13522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13524 = 8'h18 == r_count_66_io_out ? io_r_24_b : _GEN_13523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13525 = 8'h19 == r_count_66_io_out ? io_r_25_b : _GEN_13524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13526 = 8'h1a == r_count_66_io_out ? io_r_26_b : _GEN_13525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13527 = 8'h1b == r_count_66_io_out ? io_r_27_b : _GEN_13526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13528 = 8'h1c == r_count_66_io_out ? io_r_28_b : _GEN_13527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13529 = 8'h1d == r_count_66_io_out ? io_r_29_b : _GEN_13528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13530 = 8'h1e == r_count_66_io_out ? io_r_30_b : _GEN_13529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13531 = 8'h1f == r_count_66_io_out ? io_r_31_b : _GEN_13530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13532 = 8'h20 == r_count_66_io_out ? io_r_32_b : _GEN_13531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13533 = 8'h21 == r_count_66_io_out ? io_r_33_b : _GEN_13532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13534 = 8'h22 == r_count_66_io_out ? io_r_34_b : _GEN_13533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13535 = 8'h23 == r_count_66_io_out ? io_r_35_b : _GEN_13534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13536 = 8'h24 == r_count_66_io_out ? io_r_36_b : _GEN_13535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13537 = 8'h25 == r_count_66_io_out ? io_r_37_b : _GEN_13536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13538 = 8'h26 == r_count_66_io_out ? io_r_38_b : _GEN_13537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13539 = 8'h27 == r_count_66_io_out ? io_r_39_b : _GEN_13538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13540 = 8'h28 == r_count_66_io_out ? io_r_40_b : _GEN_13539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13541 = 8'h29 == r_count_66_io_out ? io_r_41_b : _GEN_13540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13542 = 8'h2a == r_count_66_io_out ? io_r_42_b : _GEN_13541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13543 = 8'h2b == r_count_66_io_out ? io_r_43_b : _GEN_13542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13544 = 8'h2c == r_count_66_io_out ? io_r_44_b : _GEN_13543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13545 = 8'h2d == r_count_66_io_out ? io_r_45_b : _GEN_13544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13546 = 8'h2e == r_count_66_io_out ? io_r_46_b : _GEN_13545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13547 = 8'h2f == r_count_66_io_out ? io_r_47_b : _GEN_13546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13548 = 8'h30 == r_count_66_io_out ? io_r_48_b : _GEN_13547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13549 = 8'h31 == r_count_66_io_out ? io_r_49_b : _GEN_13548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13550 = 8'h32 == r_count_66_io_out ? io_r_50_b : _GEN_13549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13551 = 8'h33 == r_count_66_io_out ? io_r_51_b : _GEN_13550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13552 = 8'h34 == r_count_66_io_out ? io_r_52_b : _GEN_13551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13553 = 8'h35 == r_count_66_io_out ? io_r_53_b : _GEN_13552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13554 = 8'h36 == r_count_66_io_out ? io_r_54_b : _GEN_13553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13555 = 8'h37 == r_count_66_io_out ? io_r_55_b : _GEN_13554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13556 = 8'h38 == r_count_66_io_out ? io_r_56_b : _GEN_13555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13557 = 8'h39 == r_count_66_io_out ? io_r_57_b : _GEN_13556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13558 = 8'h3a == r_count_66_io_out ? io_r_58_b : _GEN_13557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13559 = 8'h3b == r_count_66_io_out ? io_r_59_b : _GEN_13558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13560 = 8'h3c == r_count_66_io_out ? io_r_60_b : _GEN_13559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13561 = 8'h3d == r_count_66_io_out ? io_r_61_b : _GEN_13560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13562 = 8'h3e == r_count_66_io_out ? io_r_62_b : _GEN_13561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13563 = 8'h3f == r_count_66_io_out ? io_r_63_b : _GEN_13562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13564 = 8'h40 == r_count_66_io_out ? io_r_64_b : _GEN_13563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13565 = 8'h41 == r_count_66_io_out ? io_r_65_b : _GEN_13564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13566 = 8'h42 == r_count_66_io_out ? io_r_66_b : _GEN_13565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13567 = 8'h43 == r_count_66_io_out ? io_r_67_b : _GEN_13566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13568 = 8'h44 == r_count_66_io_out ? io_r_68_b : _GEN_13567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13569 = 8'h45 == r_count_66_io_out ? io_r_69_b : _GEN_13568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13570 = 8'h46 == r_count_66_io_out ? io_r_70_b : _GEN_13569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13571 = 8'h47 == r_count_66_io_out ? io_r_71_b : _GEN_13570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13572 = 8'h48 == r_count_66_io_out ? io_r_72_b : _GEN_13571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13573 = 8'h49 == r_count_66_io_out ? io_r_73_b : _GEN_13572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13574 = 8'h4a == r_count_66_io_out ? io_r_74_b : _GEN_13573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13575 = 8'h4b == r_count_66_io_out ? io_r_75_b : _GEN_13574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13576 = 8'h4c == r_count_66_io_out ? io_r_76_b : _GEN_13575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13577 = 8'h4d == r_count_66_io_out ? io_r_77_b : _GEN_13576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13578 = 8'h4e == r_count_66_io_out ? io_r_78_b : _GEN_13577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13579 = 8'h4f == r_count_66_io_out ? io_r_79_b : _GEN_13578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13580 = 8'h50 == r_count_66_io_out ? io_r_80_b : _GEN_13579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13581 = 8'h51 == r_count_66_io_out ? io_r_81_b : _GEN_13580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13582 = 8'h52 == r_count_66_io_out ? io_r_82_b : _GEN_13581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13583 = 8'h53 == r_count_66_io_out ? io_r_83_b : _GEN_13582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13584 = 8'h54 == r_count_66_io_out ? io_r_84_b : _GEN_13583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13585 = 8'h55 == r_count_66_io_out ? io_r_85_b : _GEN_13584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13586 = 8'h56 == r_count_66_io_out ? io_r_86_b : _GEN_13585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13587 = 8'h57 == r_count_66_io_out ? io_r_87_b : _GEN_13586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13588 = 8'h58 == r_count_66_io_out ? io_r_88_b : _GEN_13587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13589 = 8'h59 == r_count_66_io_out ? io_r_89_b : _GEN_13588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13590 = 8'h5a == r_count_66_io_out ? io_r_90_b : _GEN_13589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13591 = 8'h5b == r_count_66_io_out ? io_r_91_b : _GEN_13590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13592 = 8'h5c == r_count_66_io_out ? io_r_92_b : _GEN_13591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13593 = 8'h5d == r_count_66_io_out ? io_r_93_b : _GEN_13592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13594 = 8'h5e == r_count_66_io_out ? io_r_94_b : _GEN_13593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13595 = 8'h5f == r_count_66_io_out ? io_r_95_b : _GEN_13594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13596 = 8'h60 == r_count_66_io_out ? io_r_96_b : _GEN_13595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13597 = 8'h61 == r_count_66_io_out ? io_r_97_b : _GEN_13596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13598 = 8'h62 == r_count_66_io_out ? io_r_98_b : _GEN_13597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13599 = 8'h63 == r_count_66_io_out ? io_r_99_b : _GEN_13598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13600 = 8'h64 == r_count_66_io_out ? io_r_100_b : _GEN_13599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13601 = 8'h65 == r_count_66_io_out ? io_r_101_b : _GEN_13600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13602 = 8'h66 == r_count_66_io_out ? io_r_102_b : _GEN_13601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13603 = 8'h67 == r_count_66_io_out ? io_r_103_b : _GEN_13602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13604 = 8'h68 == r_count_66_io_out ? io_r_104_b : _GEN_13603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13605 = 8'h69 == r_count_66_io_out ? io_r_105_b : _GEN_13604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13606 = 8'h6a == r_count_66_io_out ? io_r_106_b : _GEN_13605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13607 = 8'h6b == r_count_66_io_out ? io_r_107_b : _GEN_13606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13608 = 8'h6c == r_count_66_io_out ? io_r_108_b : _GEN_13607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13609 = 8'h6d == r_count_66_io_out ? io_r_109_b : _GEN_13608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13610 = 8'h6e == r_count_66_io_out ? io_r_110_b : _GEN_13609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13611 = 8'h6f == r_count_66_io_out ? io_r_111_b : _GEN_13610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13612 = 8'h70 == r_count_66_io_out ? io_r_112_b : _GEN_13611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13613 = 8'h71 == r_count_66_io_out ? io_r_113_b : _GEN_13612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13614 = 8'h72 == r_count_66_io_out ? io_r_114_b : _GEN_13613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13615 = 8'h73 == r_count_66_io_out ? io_r_115_b : _GEN_13614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13616 = 8'h74 == r_count_66_io_out ? io_r_116_b : _GEN_13615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13617 = 8'h75 == r_count_66_io_out ? io_r_117_b : _GEN_13616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13618 = 8'h76 == r_count_66_io_out ? io_r_118_b : _GEN_13617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13619 = 8'h77 == r_count_66_io_out ? io_r_119_b : _GEN_13618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13620 = 8'h78 == r_count_66_io_out ? io_r_120_b : _GEN_13619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13621 = 8'h79 == r_count_66_io_out ? io_r_121_b : _GEN_13620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13622 = 8'h7a == r_count_66_io_out ? io_r_122_b : _GEN_13621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13623 = 8'h7b == r_count_66_io_out ? io_r_123_b : _GEN_13622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13624 = 8'h7c == r_count_66_io_out ? io_r_124_b : _GEN_13623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13625 = 8'h7d == r_count_66_io_out ? io_r_125_b : _GEN_13624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13626 = 8'h7e == r_count_66_io_out ? io_r_126_b : _GEN_13625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13627 = 8'h7f == r_count_66_io_out ? io_r_127_b : _GEN_13626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13628 = 8'h80 == r_count_66_io_out ? io_r_128_b : _GEN_13627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13629 = 8'h81 == r_count_66_io_out ? io_r_129_b : _GEN_13628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13630 = 8'h82 == r_count_66_io_out ? io_r_130_b : _GEN_13629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13631 = 8'h83 == r_count_66_io_out ? io_r_131_b : _GEN_13630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13632 = 8'h84 == r_count_66_io_out ? io_r_132_b : _GEN_13631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13633 = 8'h85 == r_count_66_io_out ? io_r_133_b : _GEN_13632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13634 = 8'h86 == r_count_66_io_out ? io_r_134_b : _GEN_13633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13635 = 8'h87 == r_count_66_io_out ? io_r_135_b : _GEN_13634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13636 = 8'h88 == r_count_66_io_out ? io_r_136_b : _GEN_13635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13637 = 8'h89 == r_count_66_io_out ? io_r_137_b : _GEN_13636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13638 = 8'h8a == r_count_66_io_out ? io_r_138_b : _GEN_13637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13639 = 8'h8b == r_count_66_io_out ? io_r_139_b : _GEN_13638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13640 = 8'h8c == r_count_66_io_out ? io_r_140_b : _GEN_13639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13641 = 8'h8d == r_count_66_io_out ? io_r_141_b : _GEN_13640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13642 = 8'h8e == r_count_66_io_out ? io_r_142_b : _GEN_13641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13643 = 8'h8f == r_count_66_io_out ? io_r_143_b : _GEN_13642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13644 = 8'h90 == r_count_66_io_out ? io_r_144_b : _GEN_13643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13645 = 8'h91 == r_count_66_io_out ? io_r_145_b : _GEN_13644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13646 = 8'h92 == r_count_66_io_out ? io_r_146_b : _GEN_13645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13647 = 8'h93 == r_count_66_io_out ? io_r_147_b : _GEN_13646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13648 = 8'h94 == r_count_66_io_out ? io_r_148_b : _GEN_13647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13649 = 8'h95 == r_count_66_io_out ? io_r_149_b : _GEN_13648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13650 = 8'h96 == r_count_66_io_out ? io_r_150_b : _GEN_13649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13651 = 8'h97 == r_count_66_io_out ? io_r_151_b : _GEN_13650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13652 = 8'h98 == r_count_66_io_out ? io_r_152_b : _GEN_13651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13653 = 8'h99 == r_count_66_io_out ? io_r_153_b : _GEN_13652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13654 = 8'h9a == r_count_66_io_out ? io_r_154_b : _GEN_13653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13655 = 8'h9b == r_count_66_io_out ? io_r_155_b : _GEN_13654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13656 = 8'h9c == r_count_66_io_out ? io_r_156_b : _GEN_13655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13657 = 8'h9d == r_count_66_io_out ? io_r_157_b : _GEN_13656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13658 = 8'h9e == r_count_66_io_out ? io_r_158_b : _GEN_13657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13659 = 8'h9f == r_count_66_io_out ? io_r_159_b : _GEN_13658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13660 = 8'ha0 == r_count_66_io_out ? io_r_160_b : _GEN_13659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13661 = 8'ha1 == r_count_66_io_out ? io_r_161_b : _GEN_13660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13662 = 8'ha2 == r_count_66_io_out ? io_r_162_b : _GEN_13661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13663 = 8'ha3 == r_count_66_io_out ? io_r_163_b : _GEN_13662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13664 = 8'ha4 == r_count_66_io_out ? io_r_164_b : _GEN_13663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13665 = 8'ha5 == r_count_66_io_out ? io_r_165_b : _GEN_13664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13666 = 8'ha6 == r_count_66_io_out ? io_r_166_b : _GEN_13665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13667 = 8'ha7 == r_count_66_io_out ? io_r_167_b : _GEN_13666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13668 = 8'ha8 == r_count_66_io_out ? io_r_168_b : _GEN_13667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13669 = 8'ha9 == r_count_66_io_out ? io_r_169_b : _GEN_13668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13670 = 8'haa == r_count_66_io_out ? io_r_170_b : _GEN_13669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13671 = 8'hab == r_count_66_io_out ? io_r_171_b : _GEN_13670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13672 = 8'hac == r_count_66_io_out ? io_r_172_b : _GEN_13671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13673 = 8'had == r_count_66_io_out ? io_r_173_b : _GEN_13672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13674 = 8'hae == r_count_66_io_out ? io_r_174_b : _GEN_13673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13675 = 8'haf == r_count_66_io_out ? io_r_175_b : _GEN_13674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13676 = 8'hb0 == r_count_66_io_out ? io_r_176_b : _GEN_13675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13677 = 8'hb1 == r_count_66_io_out ? io_r_177_b : _GEN_13676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13678 = 8'hb2 == r_count_66_io_out ? io_r_178_b : _GEN_13677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13679 = 8'hb3 == r_count_66_io_out ? io_r_179_b : _GEN_13678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13680 = 8'hb4 == r_count_66_io_out ? io_r_180_b : _GEN_13679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13681 = 8'hb5 == r_count_66_io_out ? io_r_181_b : _GEN_13680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13682 = 8'hb6 == r_count_66_io_out ? io_r_182_b : _GEN_13681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13683 = 8'hb7 == r_count_66_io_out ? io_r_183_b : _GEN_13682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13684 = 8'hb8 == r_count_66_io_out ? io_r_184_b : _GEN_13683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13685 = 8'hb9 == r_count_66_io_out ? io_r_185_b : _GEN_13684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13686 = 8'hba == r_count_66_io_out ? io_r_186_b : _GEN_13685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13687 = 8'hbb == r_count_66_io_out ? io_r_187_b : _GEN_13686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13688 = 8'hbc == r_count_66_io_out ? io_r_188_b : _GEN_13687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13689 = 8'hbd == r_count_66_io_out ? io_r_189_b : _GEN_13688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13690 = 8'hbe == r_count_66_io_out ? io_r_190_b : _GEN_13689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13691 = 8'hbf == r_count_66_io_out ? io_r_191_b : _GEN_13690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13692 = 8'hc0 == r_count_66_io_out ? io_r_192_b : _GEN_13691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13693 = 8'hc1 == r_count_66_io_out ? io_r_193_b : _GEN_13692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13694 = 8'hc2 == r_count_66_io_out ? io_r_194_b : _GEN_13693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13695 = 8'hc3 == r_count_66_io_out ? io_r_195_b : _GEN_13694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13696 = 8'hc4 == r_count_66_io_out ? io_r_196_b : _GEN_13695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13697 = 8'hc5 == r_count_66_io_out ? io_r_197_b : _GEN_13696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13698 = 8'hc6 == r_count_66_io_out ? io_r_198_b : _GEN_13697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13701 = 8'h1 == r_count_67_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13702 = 8'h2 == r_count_67_io_out ? io_r_2_b : _GEN_13701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13703 = 8'h3 == r_count_67_io_out ? io_r_3_b : _GEN_13702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13704 = 8'h4 == r_count_67_io_out ? io_r_4_b : _GEN_13703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13705 = 8'h5 == r_count_67_io_out ? io_r_5_b : _GEN_13704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13706 = 8'h6 == r_count_67_io_out ? io_r_6_b : _GEN_13705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13707 = 8'h7 == r_count_67_io_out ? io_r_7_b : _GEN_13706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13708 = 8'h8 == r_count_67_io_out ? io_r_8_b : _GEN_13707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13709 = 8'h9 == r_count_67_io_out ? io_r_9_b : _GEN_13708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13710 = 8'ha == r_count_67_io_out ? io_r_10_b : _GEN_13709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13711 = 8'hb == r_count_67_io_out ? io_r_11_b : _GEN_13710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13712 = 8'hc == r_count_67_io_out ? io_r_12_b : _GEN_13711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13713 = 8'hd == r_count_67_io_out ? io_r_13_b : _GEN_13712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13714 = 8'he == r_count_67_io_out ? io_r_14_b : _GEN_13713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13715 = 8'hf == r_count_67_io_out ? io_r_15_b : _GEN_13714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13716 = 8'h10 == r_count_67_io_out ? io_r_16_b : _GEN_13715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13717 = 8'h11 == r_count_67_io_out ? io_r_17_b : _GEN_13716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13718 = 8'h12 == r_count_67_io_out ? io_r_18_b : _GEN_13717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13719 = 8'h13 == r_count_67_io_out ? io_r_19_b : _GEN_13718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13720 = 8'h14 == r_count_67_io_out ? io_r_20_b : _GEN_13719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13721 = 8'h15 == r_count_67_io_out ? io_r_21_b : _GEN_13720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13722 = 8'h16 == r_count_67_io_out ? io_r_22_b : _GEN_13721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13723 = 8'h17 == r_count_67_io_out ? io_r_23_b : _GEN_13722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13724 = 8'h18 == r_count_67_io_out ? io_r_24_b : _GEN_13723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13725 = 8'h19 == r_count_67_io_out ? io_r_25_b : _GEN_13724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13726 = 8'h1a == r_count_67_io_out ? io_r_26_b : _GEN_13725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13727 = 8'h1b == r_count_67_io_out ? io_r_27_b : _GEN_13726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13728 = 8'h1c == r_count_67_io_out ? io_r_28_b : _GEN_13727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13729 = 8'h1d == r_count_67_io_out ? io_r_29_b : _GEN_13728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13730 = 8'h1e == r_count_67_io_out ? io_r_30_b : _GEN_13729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13731 = 8'h1f == r_count_67_io_out ? io_r_31_b : _GEN_13730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13732 = 8'h20 == r_count_67_io_out ? io_r_32_b : _GEN_13731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13733 = 8'h21 == r_count_67_io_out ? io_r_33_b : _GEN_13732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13734 = 8'h22 == r_count_67_io_out ? io_r_34_b : _GEN_13733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13735 = 8'h23 == r_count_67_io_out ? io_r_35_b : _GEN_13734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13736 = 8'h24 == r_count_67_io_out ? io_r_36_b : _GEN_13735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13737 = 8'h25 == r_count_67_io_out ? io_r_37_b : _GEN_13736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13738 = 8'h26 == r_count_67_io_out ? io_r_38_b : _GEN_13737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13739 = 8'h27 == r_count_67_io_out ? io_r_39_b : _GEN_13738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13740 = 8'h28 == r_count_67_io_out ? io_r_40_b : _GEN_13739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13741 = 8'h29 == r_count_67_io_out ? io_r_41_b : _GEN_13740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13742 = 8'h2a == r_count_67_io_out ? io_r_42_b : _GEN_13741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13743 = 8'h2b == r_count_67_io_out ? io_r_43_b : _GEN_13742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13744 = 8'h2c == r_count_67_io_out ? io_r_44_b : _GEN_13743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13745 = 8'h2d == r_count_67_io_out ? io_r_45_b : _GEN_13744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13746 = 8'h2e == r_count_67_io_out ? io_r_46_b : _GEN_13745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13747 = 8'h2f == r_count_67_io_out ? io_r_47_b : _GEN_13746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13748 = 8'h30 == r_count_67_io_out ? io_r_48_b : _GEN_13747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13749 = 8'h31 == r_count_67_io_out ? io_r_49_b : _GEN_13748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13750 = 8'h32 == r_count_67_io_out ? io_r_50_b : _GEN_13749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13751 = 8'h33 == r_count_67_io_out ? io_r_51_b : _GEN_13750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13752 = 8'h34 == r_count_67_io_out ? io_r_52_b : _GEN_13751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13753 = 8'h35 == r_count_67_io_out ? io_r_53_b : _GEN_13752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13754 = 8'h36 == r_count_67_io_out ? io_r_54_b : _GEN_13753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13755 = 8'h37 == r_count_67_io_out ? io_r_55_b : _GEN_13754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13756 = 8'h38 == r_count_67_io_out ? io_r_56_b : _GEN_13755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13757 = 8'h39 == r_count_67_io_out ? io_r_57_b : _GEN_13756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13758 = 8'h3a == r_count_67_io_out ? io_r_58_b : _GEN_13757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13759 = 8'h3b == r_count_67_io_out ? io_r_59_b : _GEN_13758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13760 = 8'h3c == r_count_67_io_out ? io_r_60_b : _GEN_13759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13761 = 8'h3d == r_count_67_io_out ? io_r_61_b : _GEN_13760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13762 = 8'h3e == r_count_67_io_out ? io_r_62_b : _GEN_13761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13763 = 8'h3f == r_count_67_io_out ? io_r_63_b : _GEN_13762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13764 = 8'h40 == r_count_67_io_out ? io_r_64_b : _GEN_13763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13765 = 8'h41 == r_count_67_io_out ? io_r_65_b : _GEN_13764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13766 = 8'h42 == r_count_67_io_out ? io_r_66_b : _GEN_13765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13767 = 8'h43 == r_count_67_io_out ? io_r_67_b : _GEN_13766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13768 = 8'h44 == r_count_67_io_out ? io_r_68_b : _GEN_13767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13769 = 8'h45 == r_count_67_io_out ? io_r_69_b : _GEN_13768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13770 = 8'h46 == r_count_67_io_out ? io_r_70_b : _GEN_13769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13771 = 8'h47 == r_count_67_io_out ? io_r_71_b : _GEN_13770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13772 = 8'h48 == r_count_67_io_out ? io_r_72_b : _GEN_13771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13773 = 8'h49 == r_count_67_io_out ? io_r_73_b : _GEN_13772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13774 = 8'h4a == r_count_67_io_out ? io_r_74_b : _GEN_13773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13775 = 8'h4b == r_count_67_io_out ? io_r_75_b : _GEN_13774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13776 = 8'h4c == r_count_67_io_out ? io_r_76_b : _GEN_13775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13777 = 8'h4d == r_count_67_io_out ? io_r_77_b : _GEN_13776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13778 = 8'h4e == r_count_67_io_out ? io_r_78_b : _GEN_13777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13779 = 8'h4f == r_count_67_io_out ? io_r_79_b : _GEN_13778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13780 = 8'h50 == r_count_67_io_out ? io_r_80_b : _GEN_13779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13781 = 8'h51 == r_count_67_io_out ? io_r_81_b : _GEN_13780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13782 = 8'h52 == r_count_67_io_out ? io_r_82_b : _GEN_13781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13783 = 8'h53 == r_count_67_io_out ? io_r_83_b : _GEN_13782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13784 = 8'h54 == r_count_67_io_out ? io_r_84_b : _GEN_13783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13785 = 8'h55 == r_count_67_io_out ? io_r_85_b : _GEN_13784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13786 = 8'h56 == r_count_67_io_out ? io_r_86_b : _GEN_13785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13787 = 8'h57 == r_count_67_io_out ? io_r_87_b : _GEN_13786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13788 = 8'h58 == r_count_67_io_out ? io_r_88_b : _GEN_13787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13789 = 8'h59 == r_count_67_io_out ? io_r_89_b : _GEN_13788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13790 = 8'h5a == r_count_67_io_out ? io_r_90_b : _GEN_13789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13791 = 8'h5b == r_count_67_io_out ? io_r_91_b : _GEN_13790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13792 = 8'h5c == r_count_67_io_out ? io_r_92_b : _GEN_13791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13793 = 8'h5d == r_count_67_io_out ? io_r_93_b : _GEN_13792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13794 = 8'h5e == r_count_67_io_out ? io_r_94_b : _GEN_13793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13795 = 8'h5f == r_count_67_io_out ? io_r_95_b : _GEN_13794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13796 = 8'h60 == r_count_67_io_out ? io_r_96_b : _GEN_13795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13797 = 8'h61 == r_count_67_io_out ? io_r_97_b : _GEN_13796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13798 = 8'h62 == r_count_67_io_out ? io_r_98_b : _GEN_13797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13799 = 8'h63 == r_count_67_io_out ? io_r_99_b : _GEN_13798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13800 = 8'h64 == r_count_67_io_out ? io_r_100_b : _GEN_13799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13801 = 8'h65 == r_count_67_io_out ? io_r_101_b : _GEN_13800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13802 = 8'h66 == r_count_67_io_out ? io_r_102_b : _GEN_13801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13803 = 8'h67 == r_count_67_io_out ? io_r_103_b : _GEN_13802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13804 = 8'h68 == r_count_67_io_out ? io_r_104_b : _GEN_13803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13805 = 8'h69 == r_count_67_io_out ? io_r_105_b : _GEN_13804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13806 = 8'h6a == r_count_67_io_out ? io_r_106_b : _GEN_13805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13807 = 8'h6b == r_count_67_io_out ? io_r_107_b : _GEN_13806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13808 = 8'h6c == r_count_67_io_out ? io_r_108_b : _GEN_13807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13809 = 8'h6d == r_count_67_io_out ? io_r_109_b : _GEN_13808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13810 = 8'h6e == r_count_67_io_out ? io_r_110_b : _GEN_13809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13811 = 8'h6f == r_count_67_io_out ? io_r_111_b : _GEN_13810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13812 = 8'h70 == r_count_67_io_out ? io_r_112_b : _GEN_13811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13813 = 8'h71 == r_count_67_io_out ? io_r_113_b : _GEN_13812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13814 = 8'h72 == r_count_67_io_out ? io_r_114_b : _GEN_13813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13815 = 8'h73 == r_count_67_io_out ? io_r_115_b : _GEN_13814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13816 = 8'h74 == r_count_67_io_out ? io_r_116_b : _GEN_13815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13817 = 8'h75 == r_count_67_io_out ? io_r_117_b : _GEN_13816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13818 = 8'h76 == r_count_67_io_out ? io_r_118_b : _GEN_13817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13819 = 8'h77 == r_count_67_io_out ? io_r_119_b : _GEN_13818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13820 = 8'h78 == r_count_67_io_out ? io_r_120_b : _GEN_13819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13821 = 8'h79 == r_count_67_io_out ? io_r_121_b : _GEN_13820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13822 = 8'h7a == r_count_67_io_out ? io_r_122_b : _GEN_13821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13823 = 8'h7b == r_count_67_io_out ? io_r_123_b : _GEN_13822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13824 = 8'h7c == r_count_67_io_out ? io_r_124_b : _GEN_13823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13825 = 8'h7d == r_count_67_io_out ? io_r_125_b : _GEN_13824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13826 = 8'h7e == r_count_67_io_out ? io_r_126_b : _GEN_13825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13827 = 8'h7f == r_count_67_io_out ? io_r_127_b : _GEN_13826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13828 = 8'h80 == r_count_67_io_out ? io_r_128_b : _GEN_13827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13829 = 8'h81 == r_count_67_io_out ? io_r_129_b : _GEN_13828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13830 = 8'h82 == r_count_67_io_out ? io_r_130_b : _GEN_13829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13831 = 8'h83 == r_count_67_io_out ? io_r_131_b : _GEN_13830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13832 = 8'h84 == r_count_67_io_out ? io_r_132_b : _GEN_13831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13833 = 8'h85 == r_count_67_io_out ? io_r_133_b : _GEN_13832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13834 = 8'h86 == r_count_67_io_out ? io_r_134_b : _GEN_13833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13835 = 8'h87 == r_count_67_io_out ? io_r_135_b : _GEN_13834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13836 = 8'h88 == r_count_67_io_out ? io_r_136_b : _GEN_13835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13837 = 8'h89 == r_count_67_io_out ? io_r_137_b : _GEN_13836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13838 = 8'h8a == r_count_67_io_out ? io_r_138_b : _GEN_13837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13839 = 8'h8b == r_count_67_io_out ? io_r_139_b : _GEN_13838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13840 = 8'h8c == r_count_67_io_out ? io_r_140_b : _GEN_13839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13841 = 8'h8d == r_count_67_io_out ? io_r_141_b : _GEN_13840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13842 = 8'h8e == r_count_67_io_out ? io_r_142_b : _GEN_13841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13843 = 8'h8f == r_count_67_io_out ? io_r_143_b : _GEN_13842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13844 = 8'h90 == r_count_67_io_out ? io_r_144_b : _GEN_13843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13845 = 8'h91 == r_count_67_io_out ? io_r_145_b : _GEN_13844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13846 = 8'h92 == r_count_67_io_out ? io_r_146_b : _GEN_13845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13847 = 8'h93 == r_count_67_io_out ? io_r_147_b : _GEN_13846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13848 = 8'h94 == r_count_67_io_out ? io_r_148_b : _GEN_13847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13849 = 8'h95 == r_count_67_io_out ? io_r_149_b : _GEN_13848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13850 = 8'h96 == r_count_67_io_out ? io_r_150_b : _GEN_13849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13851 = 8'h97 == r_count_67_io_out ? io_r_151_b : _GEN_13850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13852 = 8'h98 == r_count_67_io_out ? io_r_152_b : _GEN_13851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13853 = 8'h99 == r_count_67_io_out ? io_r_153_b : _GEN_13852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13854 = 8'h9a == r_count_67_io_out ? io_r_154_b : _GEN_13853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13855 = 8'h9b == r_count_67_io_out ? io_r_155_b : _GEN_13854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13856 = 8'h9c == r_count_67_io_out ? io_r_156_b : _GEN_13855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13857 = 8'h9d == r_count_67_io_out ? io_r_157_b : _GEN_13856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13858 = 8'h9e == r_count_67_io_out ? io_r_158_b : _GEN_13857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13859 = 8'h9f == r_count_67_io_out ? io_r_159_b : _GEN_13858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13860 = 8'ha0 == r_count_67_io_out ? io_r_160_b : _GEN_13859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13861 = 8'ha1 == r_count_67_io_out ? io_r_161_b : _GEN_13860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13862 = 8'ha2 == r_count_67_io_out ? io_r_162_b : _GEN_13861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13863 = 8'ha3 == r_count_67_io_out ? io_r_163_b : _GEN_13862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13864 = 8'ha4 == r_count_67_io_out ? io_r_164_b : _GEN_13863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13865 = 8'ha5 == r_count_67_io_out ? io_r_165_b : _GEN_13864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13866 = 8'ha6 == r_count_67_io_out ? io_r_166_b : _GEN_13865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13867 = 8'ha7 == r_count_67_io_out ? io_r_167_b : _GEN_13866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13868 = 8'ha8 == r_count_67_io_out ? io_r_168_b : _GEN_13867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13869 = 8'ha9 == r_count_67_io_out ? io_r_169_b : _GEN_13868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13870 = 8'haa == r_count_67_io_out ? io_r_170_b : _GEN_13869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13871 = 8'hab == r_count_67_io_out ? io_r_171_b : _GEN_13870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13872 = 8'hac == r_count_67_io_out ? io_r_172_b : _GEN_13871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13873 = 8'had == r_count_67_io_out ? io_r_173_b : _GEN_13872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13874 = 8'hae == r_count_67_io_out ? io_r_174_b : _GEN_13873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13875 = 8'haf == r_count_67_io_out ? io_r_175_b : _GEN_13874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13876 = 8'hb0 == r_count_67_io_out ? io_r_176_b : _GEN_13875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13877 = 8'hb1 == r_count_67_io_out ? io_r_177_b : _GEN_13876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13878 = 8'hb2 == r_count_67_io_out ? io_r_178_b : _GEN_13877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13879 = 8'hb3 == r_count_67_io_out ? io_r_179_b : _GEN_13878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13880 = 8'hb4 == r_count_67_io_out ? io_r_180_b : _GEN_13879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13881 = 8'hb5 == r_count_67_io_out ? io_r_181_b : _GEN_13880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13882 = 8'hb6 == r_count_67_io_out ? io_r_182_b : _GEN_13881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13883 = 8'hb7 == r_count_67_io_out ? io_r_183_b : _GEN_13882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13884 = 8'hb8 == r_count_67_io_out ? io_r_184_b : _GEN_13883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13885 = 8'hb9 == r_count_67_io_out ? io_r_185_b : _GEN_13884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13886 = 8'hba == r_count_67_io_out ? io_r_186_b : _GEN_13885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13887 = 8'hbb == r_count_67_io_out ? io_r_187_b : _GEN_13886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13888 = 8'hbc == r_count_67_io_out ? io_r_188_b : _GEN_13887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13889 = 8'hbd == r_count_67_io_out ? io_r_189_b : _GEN_13888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13890 = 8'hbe == r_count_67_io_out ? io_r_190_b : _GEN_13889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13891 = 8'hbf == r_count_67_io_out ? io_r_191_b : _GEN_13890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13892 = 8'hc0 == r_count_67_io_out ? io_r_192_b : _GEN_13891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13893 = 8'hc1 == r_count_67_io_out ? io_r_193_b : _GEN_13892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13894 = 8'hc2 == r_count_67_io_out ? io_r_194_b : _GEN_13893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13895 = 8'hc3 == r_count_67_io_out ? io_r_195_b : _GEN_13894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13896 = 8'hc4 == r_count_67_io_out ? io_r_196_b : _GEN_13895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13897 = 8'hc5 == r_count_67_io_out ? io_r_197_b : _GEN_13896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13898 = 8'hc6 == r_count_67_io_out ? io_r_198_b : _GEN_13897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13901 = 8'h1 == r_count_68_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13902 = 8'h2 == r_count_68_io_out ? io_r_2_b : _GEN_13901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13903 = 8'h3 == r_count_68_io_out ? io_r_3_b : _GEN_13902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13904 = 8'h4 == r_count_68_io_out ? io_r_4_b : _GEN_13903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13905 = 8'h5 == r_count_68_io_out ? io_r_5_b : _GEN_13904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13906 = 8'h6 == r_count_68_io_out ? io_r_6_b : _GEN_13905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13907 = 8'h7 == r_count_68_io_out ? io_r_7_b : _GEN_13906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13908 = 8'h8 == r_count_68_io_out ? io_r_8_b : _GEN_13907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13909 = 8'h9 == r_count_68_io_out ? io_r_9_b : _GEN_13908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13910 = 8'ha == r_count_68_io_out ? io_r_10_b : _GEN_13909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13911 = 8'hb == r_count_68_io_out ? io_r_11_b : _GEN_13910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13912 = 8'hc == r_count_68_io_out ? io_r_12_b : _GEN_13911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13913 = 8'hd == r_count_68_io_out ? io_r_13_b : _GEN_13912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13914 = 8'he == r_count_68_io_out ? io_r_14_b : _GEN_13913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13915 = 8'hf == r_count_68_io_out ? io_r_15_b : _GEN_13914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13916 = 8'h10 == r_count_68_io_out ? io_r_16_b : _GEN_13915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13917 = 8'h11 == r_count_68_io_out ? io_r_17_b : _GEN_13916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13918 = 8'h12 == r_count_68_io_out ? io_r_18_b : _GEN_13917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13919 = 8'h13 == r_count_68_io_out ? io_r_19_b : _GEN_13918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13920 = 8'h14 == r_count_68_io_out ? io_r_20_b : _GEN_13919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13921 = 8'h15 == r_count_68_io_out ? io_r_21_b : _GEN_13920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13922 = 8'h16 == r_count_68_io_out ? io_r_22_b : _GEN_13921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13923 = 8'h17 == r_count_68_io_out ? io_r_23_b : _GEN_13922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13924 = 8'h18 == r_count_68_io_out ? io_r_24_b : _GEN_13923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13925 = 8'h19 == r_count_68_io_out ? io_r_25_b : _GEN_13924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13926 = 8'h1a == r_count_68_io_out ? io_r_26_b : _GEN_13925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13927 = 8'h1b == r_count_68_io_out ? io_r_27_b : _GEN_13926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13928 = 8'h1c == r_count_68_io_out ? io_r_28_b : _GEN_13927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13929 = 8'h1d == r_count_68_io_out ? io_r_29_b : _GEN_13928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13930 = 8'h1e == r_count_68_io_out ? io_r_30_b : _GEN_13929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13931 = 8'h1f == r_count_68_io_out ? io_r_31_b : _GEN_13930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13932 = 8'h20 == r_count_68_io_out ? io_r_32_b : _GEN_13931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13933 = 8'h21 == r_count_68_io_out ? io_r_33_b : _GEN_13932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13934 = 8'h22 == r_count_68_io_out ? io_r_34_b : _GEN_13933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13935 = 8'h23 == r_count_68_io_out ? io_r_35_b : _GEN_13934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13936 = 8'h24 == r_count_68_io_out ? io_r_36_b : _GEN_13935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13937 = 8'h25 == r_count_68_io_out ? io_r_37_b : _GEN_13936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13938 = 8'h26 == r_count_68_io_out ? io_r_38_b : _GEN_13937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13939 = 8'h27 == r_count_68_io_out ? io_r_39_b : _GEN_13938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13940 = 8'h28 == r_count_68_io_out ? io_r_40_b : _GEN_13939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13941 = 8'h29 == r_count_68_io_out ? io_r_41_b : _GEN_13940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13942 = 8'h2a == r_count_68_io_out ? io_r_42_b : _GEN_13941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13943 = 8'h2b == r_count_68_io_out ? io_r_43_b : _GEN_13942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13944 = 8'h2c == r_count_68_io_out ? io_r_44_b : _GEN_13943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13945 = 8'h2d == r_count_68_io_out ? io_r_45_b : _GEN_13944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13946 = 8'h2e == r_count_68_io_out ? io_r_46_b : _GEN_13945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13947 = 8'h2f == r_count_68_io_out ? io_r_47_b : _GEN_13946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13948 = 8'h30 == r_count_68_io_out ? io_r_48_b : _GEN_13947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13949 = 8'h31 == r_count_68_io_out ? io_r_49_b : _GEN_13948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13950 = 8'h32 == r_count_68_io_out ? io_r_50_b : _GEN_13949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13951 = 8'h33 == r_count_68_io_out ? io_r_51_b : _GEN_13950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13952 = 8'h34 == r_count_68_io_out ? io_r_52_b : _GEN_13951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13953 = 8'h35 == r_count_68_io_out ? io_r_53_b : _GEN_13952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13954 = 8'h36 == r_count_68_io_out ? io_r_54_b : _GEN_13953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13955 = 8'h37 == r_count_68_io_out ? io_r_55_b : _GEN_13954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13956 = 8'h38 == r_count_68_io_out ? io_r_56_b : _GEN_13955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13957 = 8'h39 == r_count_68_io_out ? io_r_57_b : _GEN_13956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13958 = 8'h3a == r_count_68_io_out ? io_r_58_b : _GEN_13957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13959 = 8'h3b == r_count_68_io_out ? io_r_59_b : _GEN_13958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13960 = 8'h3c == r_count_68_io_out ? io_r_60_b : _GEN_13959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13961 = 8'h3d == r_count_68_io_out ? io_r_61_b : _GEN_13960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13962 = 8'h3e == r_count_68_io_out ? io_r_62_b : _GEN_13961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13963 = 8'h3f == r_count_68_io_out ? io_r_63_b : _GEN_13962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13964 = 8'h40 == r_count_68_io_out ? io_r_64_b : _GEN_13963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13965 = 8'h41 == r_count_68_io_out ? io_r_65_b : _GEN_13964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13966 = 8'h42 == r_count_68_io_out ? io_r_66_b : _GEN_13965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13967 = 8'h43 == r_count_68_io_out ? io_r_67_b : _GEN_13966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13968 = 8'h44 == r_count_68_io_out ? io_r_68_b : _GEN_13967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13969 = 8'h45 == r_count_68_io_out ? io_r_69_b : _GEN_13968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13970 = 8'h46 == r_count_68_io_out ? io_r_70_b : _GEN_13969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13971 = 8'h47 == r_count_68_io_out ? io_r_71_b : _GEN_13970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13972 = 8'h48 == r_count_68_io_out ? io_r_72_b : _GEN_13971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13973 = 8'h49 == r_count_68_io_out ? io_r_73_b : _GEN_13972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13974 = 8'h4a == r_count_68_io_out ? io_r_74_b : _GEN_13973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13975 = 8'h4b == r_count_68_io_out ? io_r_75_b : _GEN_13974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13976 = 8'h4c == r_count_68_io_out ? io_r_76_b : _GEN_13975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13977 = 8'h4d == r_count_68_io_out ? io_r_77_b : _GEN_13976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13978 = 8'h4e == r_count_68_io_out ? io_r_78_b : _GEN_13977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13979 = 8'h4f == r_count_68_io_out ? io_r_79_b : _GEN_13978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13980 = 8'h50 == r_count_68_io_out ? io_r_80_b : _GEN_13979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13981 = 8'h51 == r_count_68_io_out ? io_r_81_b : _GEN_13980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13982 = 8'h52 == r_count_68_io_out ? io_r_82_b : _GEN_13981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13983 = 8'h53 == r_count_68_io_out ? io_r_83_b : _GEN_13982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13984 = 8'h54 == r_count_68_io_out ? io_r_84_b : _GEN_13983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13985 = 8'h55 == r_count_68_io_out ? io_r_85_b : _GEN_13984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13986 = 8'h56 == r_count_68_io_out ? io_r_86_b : _GEN_13985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13987 = 8'h57 == r_count_68_io_out ? io_r_87_b : _GEN_13986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13988 = 8'h58 == r_count_68_io_out ? io_r_88_b : _GEN_13987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13989 = 8'h59 == r_count_68_io_out ? io_r_89_b : _GEN_13988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13990 = 8'h5a == r_count_68_io_out ? io_r_90_b : _GEN_13989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13991 = 8'h5b == r_count_68_io_out ? io_r_91_b : _GEN_13990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13992 = 8'h5c == r_count_68_io_out ? io_r_92_b : _GEN_13991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13993 = 8'h5d == r_count_68_io_out ? io_r_93_b : _GEN_13992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13994 = 8'h5e == r_count_68_io_out ? io_r_94_b : _GEN_13993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13995 = 8'h5f == r_count_68_io_out ? io_r_95_b : _GEN_13994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13996 = 8'h60 == r_count_68_io_out ? io_r_96_b : _GEN_13995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13997 = 8'h61 == r_count_68_io_out ? io_r_97_b : _GEN_13996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13998 = 8'h62 == r_count_68_io_out ? io_r_98_b : _GEN_13997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_13999 = 8'h63 == r_count_68_io_out ? io_r_99_b : _GEN_13998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14000 = 8'h64 == r_count_68_io_out ? io_r_100_b : _GEN_13999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14001 = 8'h65 == r_count_68_io_out ? io_r_101_b : _GEN_14000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14002 = 8'h66 == r_count_68_io_out ? io_r_102_b : _GEN_14001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14003 = 8'h67 == r_count_68_io_out ? io_r_103_b : _GEN_14002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14004 = 8'h68 == r_count_68_io_out ? io_r_104_b : _GEN_14003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14005 = 8'h69 == r_count_68_io_out ? io_r_105_b : _GEN_14004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14006 = 8'h6a == r_count_68_io_out ? io_r_106_b : _GEN_14005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14007 = 8'h6b == r_count_68_io_out ? io_r_107_b : _GEN_14006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14008 = 8'h6c == r_count_68_io_out ? io_r_108_b : _GEN_14007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14009 = 8'h6d == r_count_68_io_out ? io_r_109_b : _GEN_14008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14010 = 8'h6e == r_count_68_io_out ? io_r_110_b : _GEN_14009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14011 = 8'h6f == r_count_68_io_out ? io_r_111_b : _GEN_14010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14012 = 8'h70 == r_count_68_io_out ? io_r_112_b : _GEN_14011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14013 = 8'h71 == r_count_68_io_out ? io_r_113_b : _GEN_14012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14014 = 8'h72 == r_count_68_io_out ? io_r_114_b : _GEN_14013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14015 = 8'h73 == r_count_68_io_out ? io_r_115_b : _GEN_14014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14016 = 8'h74 == r_count_68_io_out ? io_r_116_b : _GEN_14015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14017 = 8'h75 == r_count_68_io_out ? io_r_117_b : _GEN_14016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14018 = 8'h76 == r_count_68_io_out ? io_r_118_b : _GEN_14017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14019 = 8'h77 == r_count_68_io_out ? io_r_119_b : _GEN_14018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14020 = 8'h78 == r_count_68_io_out ? io_r_120_b : _GEN_14019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14021 = 8'h79 == r_count_68_io_out ? io_r_121_b : _GEN_14020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14022 = 8'h7a == r_count_68_io_out ? io_r_122_b : _GEN_14021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14023 = 8'h7b == r_count_68_io_out ? io_r_123_b : _GEN_14022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14024 = 8'h7c == r_count_68_io_out ? io_r_124_b : _GEN_14023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14025 = 8'h7d == r_count_68_io_out ? io_r_125_b : _GEN_14024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14026 = 8'h7e == r_count_68_io_out ? io_r_126_b : _GEN_14025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14027 = 8'h7f == r_count_68_io_out ? io_r_127_b : _GEN_14026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14028 = 8'h80 == r_count_68_io_out ? io_r_128_b : _GEN_14027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14029 = 8'h81 == r_count_68_io_out ? io_r_129_b : _GEN_14028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14030 = 8'h82 == r_count_68_io_out ? io_r_130_b : _GEN_14029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14031 = 8'h83 == r_count_68_io_out ? io_r_131_b : _GEN_14030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14032 = 8'h84 == r_count_68_io_out ? io_r_132_b : _GEN_14031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14033 = 8'h85 == r_count_68_io_out ? io_r_133_b : _GEN_14032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14034 = 8'h86 == r_count_68_io_out ? io_r_134_b : _GEN_14033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14035 = 8'h87 == r_count_68_io_out ? io_r_135_b : _GEN_14034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14036 = 8'h88 == r_count_68_io_out ? io_r_136_b : _GEN_14035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14037 = 8'h89 == r_count_68_io_out ? io_r_137_b : _GEN_14036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14038 = 8'h8a == r_count_68_io_out ? io_r_138_b : _GEN_14037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14039 = 8'h8b == r_count_68_io_out ? io_r_139_b : _GEN_14038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14040 = 8'h8c == r_count_68_io_out ? io_r_140_b : _GEN_14039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14041 = 8'h8d == r_count_68_io_out ? io_r_141_b : _GEN_14040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14042 = 8'h8e == r_count_68_io_out ? io_r_142_b : _GEN_14041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14043 = 8'h8f == r_count_68_io_out ? io_r_143_b : _GEN_14042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14044 = 8'h90 == r_count_68_io_out ? io_r_144_b : _GEN_14043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14045 = 8'h91 == r_count_68_io_out ? io_r_145_b : _GEN_14044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14046 = 8'h92 == r_count_68_io_out ? io_r_146_b : _GEN_14045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14047 = 8'h93 == r_count_68_io_out ? io_r_147_b : _GEN_14046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14048 = 8'h94 == r_count_68_io_out ? io_r_148_b : _GEN_14047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14049 = 8'h95 == r_count_68_io_out ? io_r_149_b : _GEN_14048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14050 = 8'h96 == r_count_68_io_out ? io_r_150_b : _GEN_14049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14051 = 8'h97 == r_count_68_io_out ? io_r_151_b : _GEN_14050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14052 = 8'h98 == r_count_68_io_out ? io_r_152_b : _GEN_14051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14053 = 8'h99 == r_count_68_io_out ? io_r_153_b : _GEN_14052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14054 = 8'h9a == r_count_68_io_out ? io_r_154_b : _GEN_14053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14055 = 8'h9b == r_count_68_io_out ? io_r_155_b : _GEN_14054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14056 = 8'h9c == r_count_68_io_out ? io_r_156_b : _GEN_14055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14057 = 8'h9d == r_count_68_io_out ? io_r_157_b : _GEN_14056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14058 = 8'h9e == r_count_68_io_out ? io_r_158_b : _GEN_14057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14059 = 8'h9f == r_count_68_io_out ? io_r_159_b : _GEN_14058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14060 = 8'ha0 == r_count_68_io_out ? io_r_160_b : _GEN_14059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14061 = 8'ha1 == r_count_68_io_out ? io_r_161_b : _GEN_14060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14062 = 8'ha2 == r_count_68_io_out ? io_r_162_b : _GEN_14061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14063 = 8'ha3 == r_count_68_io_out ? io_r_163_b : _GEN_14062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14064 = 8'ha4 == r_count_68_io_out ? io_r_164_b : _GEN_14063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14065 = 8'ha5 == r_count_68_io_out ? io_r_165_b : _GEN_14064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14066 = 8'ha6 == r_count_68_io_out ? io_r_166_b : _GEN_14065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14067 = 8'ha7 == r_count_68_io_out ? io_r_167_b : _GEN_14066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14068 = 8'ha8 == r_count_68_io_out ? io_r_168_b : _GEN_14067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14069 = 8'ha9 == r_count_68_io_out ? io_r_169_b : _GEN_14068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14070 = 8'haa == r_count_68_io_out ? io_r_170_b : _GEN_14069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14071 = 8'hab == r_count_68_io_out ? io_r_171_b : _GEN_14070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14072 = 8'hac == r_count_68_io_out ? io_r_172_b : _GEN_14071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14073 = 8'had == r_count_68_io_out ? io_r_173_b : _GEN_14072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14074 = 8'hae == r_count_68_io_out ? io_r_174_b : _GEN_14073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14075 = 8'haf == r_count_68_io_out ? io_r_175_b : _GEN_14074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14076 = 8'hb0 == r_count_68_io_out ? io_r_176_b : _GEN_14075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14077 = 8'hb1 == r_count_68_io_out ? io_r_177_b : _GEN_14076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14078 = 8'hb2 == r_count_68_io_out ? io_r_178_b : _GEN_14077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14079 = 8'hb3 == r_count_68_io_out ? io_r_179_b : _GEN_14078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14080 = 8'hb4 == r_count_68_io_out ? io_r_180_b : _GEN_14079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14081 = 8'hb5 == r_count_68_io_out ? io_r_181_b : _GEN_14080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14082 = 8'hb6 == r_count_68_io_out ? io_r_182_b : _GEN_14081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14083 = 8'hb7 == r_count_68_io_out ? io_r_183_b : _GEN_14082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14084 = 8'hb8 == r_count_68_io_out ? io_r_184_b : _GEN_14083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14085 = 8'hb9 == r_count_68_io_out ? io_r_185_b : _GEN_14084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14086 = 8'hba == r_count_68_io_out ? io_r_186_b : _GEN_14085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14087 = 8'hbb == r_count_68_io_out ? io_r_187_b : _GEN_14086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14088 = 8'hbc == r_count_68_io_out ? io_r_188_b : _GEN_14087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14089 = 8'hbd == r_count_68_io_out ? io_r_189_b : _GEN_14088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14090 = 8'hbe == r_count_68_io_out ? io_r_190_b : _GEN_14089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14091 = 8'hbf == r_count_68_io_out ? io_r_191_b : _GEN_14090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14092 = 8'hc0 == r_count_68_io_out ? io_r_192_b : _GEN_14091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14093 = 8'hc1 == r_count_68_io_out ? io_r_193_b : _GEN_14092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14094 = 8'hc2 == r_count_68_io_out ? io_r_194_b : _GEN_14093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14095 = 8'hc3 == r_count_68_io_out ? io_r_195_b : _GEN_14094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14096 = 8'hc4 == r_count_68_io_out ? io_r_196_b : _GEN_14095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14097 = 8'hc5 == r_count_68_io_out ? io_r_197_b : _GEN_14096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14098 = 8'hc6 == r_count_68_io_out ? io_r_198_b : _GEN_14097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14101 = 8'h1 == r_count_69_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14102 = 8'h2 == r_count_69_io_out ? io_r_2_b : _GEN_14101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14103 = 8'h3 == r_count_69_io_out ? io_r_3_b : _GEN_14102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14104 = 8'h4 == r_count_69_io_out ? io_r_4_b : _GEN_14103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14105 = 8'h5 == r_count_69_io_out ? io_r_5_b : _GEN_14104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14106 = 8'h6 == r_count_69_io_out ? io_r_6_b : _GEN_14105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14107 = 8'h7 == r_count_69_io_out ? io_r_7_b : _GEN_14106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14108 = 8'h8 == r_count_69_io_out ? io_r_8_b : _GEN_14107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14109 = 8'h9 == r_count_69_io_out ? io_r_9_b : _GEN_14108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14110 = 8'ha == r_count_69_io_out ? io_r_10_b : _GEN_14109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14111 = 8'hb == r_count_69_io_out ? io_r_11_b : _GEN_14110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14112 = 8'hc == r_count_69_io_out ? io_r_12_b : _GEN_14111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14113 = 8'hd == r_count_69_io_out ? io_r_13_b : _GEN_14112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14114 = 8'he == r_count_69_io_out ? io_r_14_b : _GEN_14113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14115 = 8'hf == r_count_69_io_out ? io_r_15_b : _GEN_14114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14116 = 8'h10 == r_count_69_io_out ? io_r_16_b : _GEN_14115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14117 = 8'h11 == r_count_69_io_out ? io_r_17_b : _GEN_14116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14118 = 8'h12 == r_count_69_io_out ? io_r_18_b : _GEN_14117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14119 = 8'h13 == r_count_69_io_out ? io_r_19_b : _GEN_14118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14120 = 8'h14 == r_count_69_io_out ? io_r_20_b : _GEN_14119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14121 = 8'h15 == r_count_69_io_out ? io_r_21_b : _GEN_14120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14122 = 8'h16 == r_count_69_io_out ? io_r_22_b : _GEN_14121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14123 = 8'h17 == r_count_69_io_out ? io_r_23_b : _GEN_14122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14124 = 8'h18 == r_count_69_io_out ? io_r_24_b : _GEN_14123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14125 = 8'h19 == r_count_69_io_out ? io_r_25_b : _GEN_14124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14126 = 8'h1a == r_count_69_io_out ? io_r_26_b : _GEN_14125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14127 = 8'h1b == r_count_69_io_out ? io_r_27_b : _GEN_14126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14128 = 8'h1c == r_count_69_io_out ? io_r_28_b : _GEN_14127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14129 = 8'h1d == r_count_69_io_out ? io_r_29_b : _GEN_14128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14130 = 8'h1e == r_count_69_io_out ? io_r_30_b : _GEN_14129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14131 = 8'h1f == r_count_69_io_out ? io_r_31_b : _GEN_14130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14132 = 8'h20 == r_count_69_io_out ? io_r_32_b : _GEN_14131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14133 = 8'h21 == r_count_69_io_out ? io_r_33_b : _GEN_14132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14134 = 8'h22 == r_count_69_io_out ? io_r_34_b : _GEN_14133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14135 = 8'h23 == r_count_69_io_out ? io_r_35_b : _GEN_14134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14136 = 8'h24 == r_count_69_io_out ? io_r_36_b : _GEN_14135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14137 = 8'h25 == r_count_69_io_out ? io_r_37_b : _GEN_14136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14138 = 8'h26 == r_count_69_io_out ? io_r_38_b : _GEN_14137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14139 = 8'h27 == r_count_69_io_out ? io_r_39_b : _GEN_14138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14140 = 8'h28 == r_count_69_io_out ? io_r_40_b : _GEN_14139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14141 = 8'h29 == r_count_69_io_out ? io_r_41_b : _GEN_14140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14142 = 8'h2a == r_count_69_io_out ? io_r_42_b : _GEN_14141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14143 = 8'h2b == r_count_69_io_out ? io_r_43_b : _GEN_14142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14144 = 8'h2c == r_count_69_io_out ? io_r_44_b : _GEN_14143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14145 = 8'h2d == r_count_69_io_out ? io_r_45_b : _GEN_14144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14146 = 8'h2e == r_count_69_io_out ? io_r_46_b : _GEN_14145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14147 = 8'h2f == r_count_69_io_out ? io_r_47_b : _GEN_14146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14148 = 8'h30 == r_count_69_io_out ? io_r_48_b : _GEN_14147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14149 = 8'h31 == r_count_69_io_out ? io_r_49_b : _GEN_14148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14150 = 8'h32 == r_count_69_io_out ? io_r_50_b : _GEN_14149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14151 = 8'h33 == r_count_69_io_out ? io_r_51_b : _GEN_14150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14152 = 8'h34 == r_count_69_io_out ? io_r_52_b : _GEN_14151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14153 = 8'h35 == r_count_69_io_out ? io_r_53_b : _GEN_14152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14154 = 8'h36 == r_count_69_io_out ? io_r_54_b : _GEN_14153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14155 = 8'h37 == r_count_69_io_out ? io_r_55_b : _GEN_14154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14156 = 8'h38 == r_count_69_io_out ? io_r_56_b : _GEN_14155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14157 = 8'h39 == r_count_69_io_out ? io_r_57_b : _GEN_14156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14158 = 8'h3a == r_count_69_io_out ? io_r_58_b : _GEN_14157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14159 = 8'h3b == r_count_69_io_out ? io_r_59_b : _GEN_14158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14160 = 8'h3c == r_count_69_io_out ? io_r_60_b : _GEN_14159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14161 = 8'h3d == r_count_69_io_out ? io_r_61_b : _GEN_14160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14162 = 8'h3e == r_count_69_io_out ? io_r_62_b : _GEN_14161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14163 = 8'h3f == r_count_69_io_out ? io_r_63_b : _GEN_14162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14164 = 8'h40 == r_count_69_io_out ? io_r_64_b : _GEN_14163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14165 = 8'h41 == r_count_69_io_out ? io_r_65_b : _GEN_14164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14166 = 8'h42 == r_count_69_io_out ? io_r_66_b : _GEN_14165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14167 = 8'h43 == r_count_69_io_out ? io_r_67_b : _GEN_14166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14168 = 8'h44 == r_count_69_io_out ? io_r_68_b : _GEN_14167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14169 = 8'h45 == r_count_69_io_out ? io_r_69_b : _GEN_14168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14170 = 8'h46 == r_count_69_io_out ? io_r_70_b : _GEN_14169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14171 = 8'h47 == r_count_69_io_out ? io_r_71_b : _GEN_14170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14172 = 8'h48 == r_count_69_io_out ? io_r_72_b : _GEN_14171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14173 = 8'h49 == r_count_69_io_out ? io_r_73_b : _GEN_14172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14174 = 8'h4a == r_count_69_io_out ? io_r_74_b : _GEN_14173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14175 = 8'h4b == r_count_69_io_out ? io_r_75_b : _GEN_14174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14176 = 8'h4c == r_count_69_io_out ? io_r_76_b : _GEN_14175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14177 = 8'h4d == r_count_69_io_out ? io_r_77_b : _GEN_14176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14178 = 8'h4e == r_count_69_io_out ? io_r_78_b : _GEN_14177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14179 = 8'h4f == r_count_69_io_out ? io_r_79_b : _GEN_14178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14180 = 8'h50 == r_count_69_io_out ? io_r_80_b : _GEN_14179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14181 = 8'h51 == r_count_69_io_out ? io_r_81_b : _GEN_14180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14182 = 8'h52 == r_count_69_io_out ? io_r_82_b : _GEN_14181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14183 = 8'h53 == r_count_69_io_out ? io_r_83_b : _GEN_14182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14184 = 8'h54 == r_count_69_io_out ? io_r_84_b : _GEN_14183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14185 = 8'h55 == r_count_69_io_out ? io_r_85_b : _GEN_14184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14186 = 8'h56 == r_count_69_io_out ? io_r_86_b : _GEN_14185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14187 = 8'h57 == r_count_69_io_out ? io_r_87_b : _GEN_14186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14188 = 8'h58 == r_count_69_io_out ? io_r_88_b : _GEN_14187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14189 = 8'h59 == r_count_69_io_out ? io_r_89_b : _GEN_14188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14190 = 8'h5a == r_count_69_io_out ? io_r_90_b : _GEN_14189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14191 = 8'h5b == r_count_69_io_out ? io_r_91_b : _GEN_14190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14192 = 8'h5c == r_count_69_io_out ? io_r_92_b : _GEN_14191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14193 = 8'h5d == r_count_69_io_out ? io_r_93_b : _GEN_14192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14194 = 8'h5e == r_count_69_io_out ? io_r_94_b : _GEN_14193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14195 = 8'h5f == r_count_69_io_out ? io_r_95_b : _GEN_14194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14196 = 8'h60 == r_count_69_io_out ? io_r_96_b : _GEN_14195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14197 = 8'h61 == r_count_69_io_out ? io_r_97_b : _GEN_14196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14198 = 8'h62 == r_count_69_io_out ? io_r_98_b : _GEN_14197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14199 = 8'h63 == r_count_69_io_out ? io_r_99_b : _GEN_14198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14200 = 8'h64 == r_count_69_io_out ? io_r_100_b : _GEN_14199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14201 = 8'h65 == r_count_69_io_out ? io_r_101_b : _GEN_14200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14202 = 8'h66 == r_count_69_io_out ? io_r_102_b : _GEN_14201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14203 = 8'h67 == r_count_69_io_out ? io_r_103_b : _GEN_14202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14204 = 8'h68 == r_count_69_io_out ? io_r_104_b : _GEN_14203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14205 = 8'h69 == r_count_69_io_out ? io_r_105_b : _GEN_14204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14206 = 8'h6a == r_count_69_io_out ? io_r_106_b : _GEN_14205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14207 = 8'h6b == r_count_69_io_out ? io_r_107_b : _GEN_14206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14208 = 8'h6c == r_count_69_io_out ? io_r_108_b : _GEN_14207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14209 = 8'h6d == r_count_69_io_out ? io_r_109_b : _GEN_14208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14210 = 8'h6e == r_count_69_io_out ? io_r_110_b : _GEN_14209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14211 = 8'h6f == r_count_69_io_out ? io_r_111_b : _GEN_14210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14212 = 8'h70 == r_count_69_io_out ? io_r_112_b : _GEN_14211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14213 = 8'h71 == r_count_69_io_out ? io_r_113_b : _GEN_14212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14214 = 8'h72 == r_count_69_io_out ? io_r_114_b : _GEN_14213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14215 = 8'h73 == r_count_69_io_out ? io_r_115_b : _GEN_14214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14216 = 8'h74 == r_count_69_io_out ? io_r_116_b : _GEN_14215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14217 = 8'h75 == r_count_69_io_out ? io_r_117_b : _GEN_14216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14218 = 8'h76 == r_count_69_io_out ? io_r_118_b : _GEN_14217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14219 = 8'h77 == r_count_69_io_out ? io_r_119_b : _GEN_14218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14220 = 8'h78 == r_count_69_io_out ? io_r_120_b : _GEN_14219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14221 = 8'h79 == r_count_69_io_out ? io_r_121_b : _GEN_14220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14222 = 8'h7a == r_count_69_io_out ? io_r_122_b : _GEN_14221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14223 = 8'h7b == r_count_69_io_out ? io_r_123_b : _GEN_14222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14224 = 8'h7c == r_count_69_io_out ? io_r_124_b : _GEN_14223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14225 = 8'h7d == r_count_69_io_out ? io_r_125_b : _GEN_14224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14226 = 8'h7e == r_count_69_io_out ? io_r_126_b : _GEN_14225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14227 = 8'h7f == r_count_69_io_out ? io_r_127_b : _GEN_14226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14228 = 8'h80 == r_count_69_io_out ? io_r_128_b : _GEN_14227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14229 = 8'h81 == r_count_69_io_out ? io_r_129_b : _GEN_14228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14230 = 8'h82 == r_count_69_io_out ? io_r_130_b : _GEN_14229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14231 = 8'h83 == r_count_69_io_out ? io_r_131_b : _GEN_14230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14232 = 8'h84 == r_count_69_io_out ? io_r_132_b : _GEN_14231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14233 = 8'h85 == r_count_69_io_out ? io_r_133_b : _GEN_14232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14234 = 8'h86 == r_count_69_io_out ? io_r_134_b : _GEN_14233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14235 = 8'h87 == r_count_69_io_out ? io_r_135_b : _GEN_14234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14236 = 8'h88 == r_count_69_io_out ? io_r_136_b : _GEN_14235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14237 = 8'h89 == r_count_69_io_out ? io_r_137_b : _GEN_14236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14238 = 8'h8a == r_count_69_io_out ? io_r_138_b : _GEN_14237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14239 = 8'h8b == r_count_69_io_out ? io_r_139_b : _GEN_14238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14240 = 8'h8c == r_count_69_io_out ? io_r_140_b : _GEN_14239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14241 = 8'h8d == r_count_69_io_out ? io_r_141_b : _GEN_14240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14242 = 8'h8e == r_count_69_io_out ? io_r_142_b : _GEN_14241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14243 = 8'h8f == r_count_69_io_out ? io_r_143_b : _GEN_14242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14244 = 8'h90 == r_count_69_io_out ? io_r_144_b : _GEN_14243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14245 = 8'h91 == r_count_69_io_out ? io_r_145_b : _GEN_14244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14246 = 8'h92 == r_count_69_io_out ? io_r_146_b : _GEN_14245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14247 = 8'h93 == r_count_69_io_out ? io_r_147_b : _GEN_14246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14248 = 8'h94 == r_count_69_io_out ? io_r_148_b : _GEN_14247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14249 = 8'h95 == r_count_69_io_out ? io_r_149_b : _GEN_14248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14250 = 8'h96 == r_count_69_io_out ? io_r_150_b : _GEN_14249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14251 = 8'h97 == r_count_69_io_out ? io_r_151_b : _GEN_14250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14252 = 8'h98 == r_count_69_io_out ? io_r_152_b : _GEN_14251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14253 = 8'h99 == r_count_69_io_out ? io_r_153_b : _GEN_14252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14254 = 8'h9a == r_count_69_io_out ? io_r_154_b : _GEN_14253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14255 = 8'h9b == r_count_69_io_out ? io_r_155_b : _GEN_14254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14256 = 8'h9c == r_count_69_io_out ? io_r_156_b : _GEN_14255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14257 = 8'h9d == r_count_69_io_out ? io_r_157_b : _GEN_14256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14258 = 8'h9e == r_count_69_io_out ? io_r_158_b : _GEN_14257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14259 = 8'h9f == r_count_69_io_out ? io_r_159_b : _GEN_14258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14260 = 8'ha0 == r_count_69_io_out ? io_r_160_b : _GEN_14259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14261 = 8'ha1 == r_count_69_io_out ? io_r_161_b : _GEN_14260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14262 = 8'ha2 == r_count_69_io_out ? io_r_162_b : _GEN_14261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14263 = 8'ha3 == r_count_69_io_out ? io_r_163_b : _GEN_14262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14264 = 8'ha4 == r_count_69_io_out ? io_r_164_b : _GEN_14263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14265 = 8'ha5 == r_count_69_io_out ? io_r_165_b : _GEN_14264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14266 = 8'ha6 == r_count_69_io_out ? io_r_166_b : _GEN_14265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14267 = 8'ha7 == r_count_69_io_out ? io_r_167_b : _GEN_14266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14268 = 8'ha8 == r_count_69_io_out ? io_r_168_b : _GEN_14267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14269 = 8'ha9 == r_count_69_io_out ? io_r_169_b : _GEN_14268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14270 = 8'haa == r_count_69_io_out ? io_r_170_b : _GEN_14269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14271 = 8'hab == r_count_69_io_out ? io_r_171_b : _GEN_14270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14272 = 8'hac == r_count_69_io_out ? io_r_172_b : _GEN_14271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14273 = 8'had == r_count_69_io_out ? io_r_173_b : _GEN_14272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14274 = 8'hae == r_count_69_io_out ? io_r_174_b : _GEN_14273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14275 = 8'haf == r_count_69_io_out ? io_r_175_b : _GEN_14274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14276 = 8'hb0 == r_count_69_io_out ? io_r_176_b : _GEN_14275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14277 = 8'hb1 == r_count_69_io_out ? io_r_177_b : _GEN_14276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14278 = 8'hb2 == r_count_69_io_out ? io_r_178_b : _GEN_14277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14279 = 8'hb3 == r_count_69_io_out ? io_r_179_b : _GEN_14278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14280 = 8'hb4 == r_count_69_io_out ? io_r_180_b : _GEN_14279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14281 = 8'hb5 == r_count_69_io_out ? io_r_181_b : _GEN_14280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14282 = 8'hb6 == r_count_69_io_out ? io_r_182_b : _GEN_14281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14283 = 8'hb7 == r_count_69_io_out ? io_r_183_b : _GEN_14282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14284 = 8'hb8 == r_count_69_io_out ? io_r_184_b : _GEN_14283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14285 = 8'hb9 == r_count_69_io_out ? io_r_185_b : _GEN_14284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14286 = 8'hba == r_count_69_io_out ? io_r_186_b : _GEN_14285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14287 = 8'hbb == r_count_69_io_out ? io_r_187_b : _GEN_14286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14288 = 8'hbc == r_count_69_io_out ? io_r_188_b : _GEN_14287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14289 = 8'hbd == r_count_69_io_out ? io_r_189_b : _GEN_14288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14290 = 8'hbe == r_count_69_io_out ? io_r_190_b : _GEN_14289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14291 = 8'hbf == r_count_69_io_out ? io_r_191_b : _GEN_14290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14292 = 8'hc0 == r_count_69_io_out ? io_r_192_b : _GEN_14291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14293 = 8'hc1 == r_count_69_io_out ? io_r_193_b : _GEN_14292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14294 = 8'hc2 == r_count_69_io_out ? io_r_194_b : _GEN_14293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14295 = 8'hc3 == r_count_69_io_out ? io_r_195_b : _GEN_14294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14296 = 8'hc4 == r_count_69_io_out ? io_r_196_b : _GEN_14295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14297 = 8'hc5 == r_count_69_io_out ? io_r_197_b : _GEN_14296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14298 = 8'hc6 == r_count_69_io_out ? io_r_198_b : _GEN_14297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14301 = 8'h1 == r_count_70_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14302 = 8'h2 == r_count_70_io_out ? io_r_2_b : _GEN_14301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14303 = 8'h3 == r_count_70_io_out ? io_r_3_b : _GEN_14302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14304 = 8'h4 == r_count_70_io_out ? io_r_4_b : _GEN_14303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14305 = 8'h5 == r_count_70_io_out ? io_r_5_b : _GEN_14304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14306 = 8'h6 == r_count_70_io_out ? io_r_6_b : _GEN_14305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14307 = 8'h7 == r_count_70_io_out ? io_r_7_b : _GEN_14306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14308 = 8'h8 == r_count_70_io_out ? io_r_8_b : _GEN_14307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14309 = 8'h9 == r_count_70_io_out ? io_r_9_b : _GEN_14308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14310 = 8'ha == r_count_70_io_out ? io_r_10_b : _GEN_14309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14311 = 8'hb == r_count_70_io_out ? io_r_11_b : _GEN_14310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14312 = 8'hc == r_count_70_io_out ? io_r_12_b : _GEN_14311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14313 = 8'hd == r_count_70_io_out ? io_r_13_b : _GEN_14312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14314 = 8'he == r_count_70_io_out ? io_r_14_b : _GEN_14313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14315 = 8'hf == r_count_70_io_out ? io_r_15_b : _GEN_14314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14316 = 8'h10 == r_count_70_io_out ? io_r_16_b : _GEN_14315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14317 = 8'h11 == r_count_70_io_out ? io_r_17_b : _GEN_14316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14318 = 8'h12 == r_count_70_io_out ? io_r_18_b : _GEN_14317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14319 = 8'h13 == r_count_70_io_out ? io_r_19_b : _GEN_14318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14320 = 8'h14 == r_count_70_io_out ? io_r_20_b : _GEN_14319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14321 = 8'h15 == r_count_70_io_out ? io_r_21_b : _GEN_14320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14322 = 8'h16 == r_count_70_io_out ? io_r_22_b : _GEN_14321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14323 = 8'h17 == r_count_70_io_out ? io_r_23_b : _GEN_14322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14324 = 8'h18 == r_count_70_io_out ? io_r_24_b : _GEN_14323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14325 = 8'h19 == r_count_70_io_out ? io_r_25_b : _GEN_14324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14326 = 8'h1a == r_count_70_io_out ? io_r_26_b : _GEN_14325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14327 = 8'h1b == r_count_70_io_out ? io_r_27_b : _GEN_14326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14328 = 8'h1c == r_count_70_io_out ? io_r_28_b : _GEN_14327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14329 = 8'h1d == r_count_70_io_out ? io_r_29_b : _GEN_14328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14330 = 8'h1e == r_count_70_io_out ? io_r_30_b : _GEN_14329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14331 = 8'h1f == r_count_70_io_out ? io_r_31_b : _GEN_14330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14332 = 8'h20 == r_count_70_io_out ? io_r_32_b : _GEN_14331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14333 = 8'h21 == r_count_70_io_out ? io_r_33_b : _GEN_14332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14334 = 8'h22 == r_count_70_io_out ? io_r_34_b : _GEN_14333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14335 = 8'h23 == r_count_70_io_out ? io_r_35_b : _GEN_14334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14336 = 8'h24 == r_count_70_io_out ? io_r_36_b : _GEN_14335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14337 = 8'h25 == r_count_70_io_out ? io_r_37_b : _GEN_14336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14338 = 8'h26 == r_count_70_io_out ? io_r_38_b : _GEN_14337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14339 = 8'h27 == r_count_70_io_out ? io_r_39_b : _GEN_14338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14340 = 8'h28 == r_count_70_io_out ? io_r_40_b : _GEN_14339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14341 = 8'h29 == r_count_70_io_out ? io_r_41_b : _GEN_14340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14342 = 8'h2a == r_count_70_io_out ? io_r_42_b : _GEN_14341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14343 = 8'h2b == r_count_70_io_out ? io_r_43_b : _GEN_14342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14344 = 8'h2c == r_count_70_io_out ? io_r_44_b : _GEN_14343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14345 = 8'h2d == r_count_70_io_out ? io_r_45_b : _GEN_14344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14346 = 8'h2e == r_count_70_io_out ? io_r_46_b : _GEN_14345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14347 = 8'h2f == r_count_70_io_out ? io_r_47_b : _GEN_14346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14348 = 8'h30 == r_count_70_io_out ? io_r_48_b : _GEN_14347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14349 = 8'h31 == r_count_70_io_out ? io_r_49_b : _GEN_14348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14350 = 8'h32 == r_count_70_io_out ? io_r_50_b : _GEN_14349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14351 = 8'h33 == r_count_70_io_out ? io_r_51_b : _GEN_14350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14352 = 8'h34 == r_count_70_io_out ? io_r_52_b : _GEN_14351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14353 = 8'h35 == r_count_70_io_out ? io_r_53_b : _GEN_14352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14354 = 8'h36 == r_count_70_io_out ? io_r_54_b : _GEN_14353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14355 = 8'h37 == r_count_70_io_out ? io_r_55_b : _GEN_14354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14356 = 8'h38 == r_count_70_io_out ? io_r_56_b : _GEN_14355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14357 = 8'h39 == r_count_70_io_out ? io_r_57_b : _GEN_14356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14358 = 8'h3a == r_count_70_io_out ? io_r_58_b : _GEN_14357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14359 = 8'h3b == r_count_70_io_out ? io_r_59_b : _GEN_14358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14360 = 8'h3c == r_count_70_io_out ? io_r_60_b : _GEN_14359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14361 = 8'h3d == r_count_70_io_out ? io_r_61_b : _GEN_14360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14362 = 8'h3e == r_count_70_io_out ? io_r_62_b : _GEN_14361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14363 = 8'h3f == r_count_70_io_out ? io_r_63_b : _GEN_14362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14364 = 8'h40 == r_count_70_io_out ? io_r_64_b : _GEN_14363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14365 = 8'h41 == r_count_70_io_out ? io_r_65_b : _GEN_14364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14366 = 8'h42 == r_count_70_io_out ? io_r_66_b : _GEN_14365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14367 = 8'h43 == r_count_70_io_out ? io_r_67_b : _GEN_14366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14368 = 8'h44 == r_count_70_io_out ? io_r_68_b : _GEN_14367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14369 = 8'h45 == r_count_70_io_out ? io_r_69_b : _GEN_14368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14370 = 8'h46 == r_count_70_io_out ? io_r_70_b : _GEN_14369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14371 = 8'h47 == r_count_70_io_out ? io_r_71_b : _GEN_14370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14372 = 8'h48 == r_count_70_io_out ? io_r_72_b : _GEN_14371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14373 = 8'h49 == r_count_70_io_out ? io_r_73_b : _GEN_14372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14374 = 8'h4a == r_count_70_io_out ? io_r_74_b : _GEN_14373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14375 = 8'h4b == r_count_70_io_out ? io_r_75_b : _GEN_14374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14376 = 8'h4c == r_count_70_io_out ? io_r_76_b : _GEN_14375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14377 = 8'h4d == r_count_70_io_out ? io_r_77_b : _GEN_14376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14378 = 8'h4e == r_count_70_io_out ? io_r_78_b : _GEN_14377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14379 = 8'h4f == r_count_70_io_out ? io_r_79_b : _GEN_14378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14380 = 8'h50 == r_count_70_io_out ? io_r_80_b : _GEN_14379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14381 = 8'h51 == r_count_70_io_out ? io_r_81_b : _GEN_14380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14382 = 8'h52 == r_count_70_io_out ? io_r_82_b : _GEN_14381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14383 = 8'h53 == r_count_70_io_out ? io_r_83_b : _GEN_14382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14384 = 8'h54 == r_count_70_io_out ? io_r_84_b : _GEN_14383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14385 = 8'h55 == r_count_70_io_out ? io_r_85_b : _GEN_14384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14386 = 8'h56 == r_count_70_io_out ? io_r_86_b : _GEN_14385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14387 = 8'h57 == r_count_70_io_out ? io_r_87_b : _GEN_14386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14388 = 8'h58 == r_count_70_io_out ? io_r_88_b : _GEN_14387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14389 = 8'h59 == r_count_70_io_out ? io_r_89_b : _GEN_14388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14390 = 8'h5a == r_count_70_io_out ? io_r_90_b : _GEN_14389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14391 = 8'h5b == r_count_70_io_out ? io_r_91_b : _GEN_14390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14392 = 8'h5c == r_count_70_io_out ? io_r_92_b : _GEN_14391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14393 = 8'h5d == r_count_70_io_out ? io_r_93_b : _GEN_14392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14394 = 8'h5e == r_count_70_io_out ? io_r_94_b : _GEN_14393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14395 = 8'h5f == r_count_70_io_out ? io_r_95_b : _GEN_14394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14396 = 8'h60 == r_count_70_io_out ? io_r_96_b : _GEN_14395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14397 = 8'h61 == r_count_70_io_out ? io_r_97_b : _GEN_14396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14398 = 8'h62 == r_count_70_io_out ? io_r_98_b : _GEN_14397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14399 = 8'h63 == r_count_70_io_out ? io_r_99_b : _GEN_14398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14400 = 8'h64 == r_count_70_io_out ? io_r_100_b : _GEN_14399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14401 = 8'h65 == r_count_70_io_out ? io_r_101_b : _GEN_14400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14402 = 8'h66 == r_count_70_io_out ? io_r_102_b : _GEN_14401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14403 = 8'h67 == r_count_70_io_out ? io_r_103_b : _GEN_14402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14404 = 8'h68 == r_count_70_io_out ? io_r_104_b : _GEN_14403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14405 = 8'h69 == r_count_70_io_out ? io_r_105_b : _GEN_14404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14406 = 8'h6a == r_count_70_io_out ? io_r_106_b : _GEN_14405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14407 = 8'h6b == r_count_70_io_out ? io_r_107_b : _GEN_14406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14408 = 8'h6c == r_count_70_io_out ? io_r_108_b : _GEN_14407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14409 = 8'h6d == r_count_70_io_out ? io_r_109_b : _GEN_14408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14410 = 8'h6e == r_count_70_io_out ? io_r_110_b : _GEN_14409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14411 = 8'h6f == r_count_70_io_out ? io_r_111_b : _GEN_14410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14412 = 8'h70 == r_count_70_io_out ? io_r_112_b : _GEN_14411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14413 = 8'h71 == r_count_70_io_out ? io_r_113_b : _GEN_14412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14414 = 8'h72 == r_count_70_io_out ? io_r_114_b : _GEN_14413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14415 = 8'h73 == r_count_70_io_out ? io_r_115_b : _GEN_14414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14416 = 8'h74 == r_count_70_io_out ? io_r_116_b : _GEN_14415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14417 = 8'h75 == r_count_70_io_out ? io_r_117_b : _GEN_14416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14418 = 8'h76 == r_count_70_io_out ? io_r_118_b : _GEN_14417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14419 = 8'h77 == r_count_70_io_out ? io_r_119_b : _GEN_14418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14420 = 8'h78 == r_count_70_io_out ? io_r_120_b : _GEN_14419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14421 = 8'h79 == r_count_70_io_out ? io_r_121_b : _GEN_14420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14422 = 8'h7a == r_count_70_io_out ? io_r_122_b : _GEN_14421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14423 = 8'h7b == r_count_70_io_out ? io_r_123_b : _GEN_14422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14424 = 8'h7c == r_count_70_io_out ? io_r_124_b : _GEN_14423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14425 = 8'h7d == r_count_70_io_out ? io_r_125_b : _GEN_14424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14426 = 8'h7e == r_count_70_io_out ? io_r_126_b : _GEN_14425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14427 = 8'h7f == r_count_70_io_out ? io_r_127_b : _GEN_14426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14428 = 8'h80 == r_count_70_io_out ? io_r_128_b : _GEN_14427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14429 = 8'h81 == r_count_70_io_out ? io_r_129_b : _GEN_14428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14430 = 8'h82 == r_count_70_io_out ? io_r_130_b : _GEN_14429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14431 = 8'h83 == r_count_70_io_out ? io_r_131_b : _GEN_14430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14432 = 8'h84 == r_count_70_io_out ? io_r_132_b : _GEN_14431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14433 = 8'h85 == r_count_70_io_out ? io_r_133_b : _GEN_14432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14434 = 8'h86 == r_count_70_io_out ? io_r_134_b : _GEN_14433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14435 = 8'h87 == r_count_70_io_out ? io_r_135_b : _GEN_14434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14436 = 8'h88 == r_count_70_io_out ? io_r_136_b : _GEN_14435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14437 = 8'h89 == r_count_70_io_out ? io_r_137_b : _GEN_14436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14438 = 8'h8a == r_count_70_io_out ? io_r_138_b : _GEN_14437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14439 = 8'h8b == r_count_70_io_out ? io_r_139_b : _GEN_14438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14440 = 8'h8c == r_count_70_io_out ? io_r_140_b : _GEN_14439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14441 = 8'h8d == r_count_70_io_out ? io_r_141_b : _GEN_14440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14442 = 8'h8e == r_count_70_io_out ? io_r_142_b : _GEN_14441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14443 = 8'h8f == r_count_70_io_out ? io_r_143_b : _GEN_14442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14444 = 8'h90 == r_count_70_io_out ? io_r_144_b : _GEN_14443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14445 = 8'h91 == r_count_70_io_out ? io_r_145_b : _GEN_14444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14446 = 8'h92 == r_count_70_io_out ? io_r_146_b : _GEN_14445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14447 = 8'h93 == r_count_70_io_out ? io_r_147_b : _GEN_14446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14448 = 8'h94 == r_count_70_io_out ? io_r_148_b : _GEN_14447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14449 = 8'h95 == r_count_70_io_out ? io_r_149_b : _GEN_14448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14450 = 8'h96 == r_count_70_io_out ? io_r_150_b : _GEN_14449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14451 = 8'h97 == r_count_70_io_out ? io_r_151_b : _GEN_14450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14452 = 8'h98 == r_count_70_io_out ? io_r_152_b : _GEN_14451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14453 = 8'h99 == r_count_70_io_out ? io_r_153_b : _GEN_14452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14454 = 8'h9a == r_count_70_io_out ? io_r_154_b : _GEN_14453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14455 = 8'h9b == r_count_70_io_out ? io_r_155_b : _GEN_14454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14456 = 8'h9c == r_count_70_io_out ? io_r_156_b : _GEN_14455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14457 = 8'h9d == r_count_70_io_out ? io_r_157_b : _GEN_14456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14458 = 8'h9e == r_count_70_io_out ? io_r_158_b : _GEN_14457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14459 = 8'h9f == r_count_70_io_out ? io_r_159_b : _GEN_14458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14460 = 8'ha0 == r_count_70_io_out ? io_r_160_b : _GEN_14459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14461 = 8'ha1 == r_count_70_io_out ? io_r_161_b : _GEN_14460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14462 = 8'ha2 == r_count_70_io_out ? io_r_162_b : _GEN_14461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14463 = 8'ha3 == r_count_70_io_out ? io_r_163_b : _GEN_14462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14464 = 8'ha4 == r_count_70_io_out ? io_r_164_b : _GEN_14463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14465 = 8'ha5 == r_count_70_io_out ? io_r_165_b : _GEN_14464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14466 = 8'ha6 == r_count_70_io_out ? io_r_166_b : _GEN_14465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14467 = 8'ha7 == r_count_70_io_out ? io_r_167_b : _GEN_14466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14468 = 8'ha8 == r_count_70_io_out ? io_r_168_b : _GEN_14467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14469 = 8'ha9 == r_count_70_io_out ? io_r_169_b : _GEN_14468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14470 = 8'haa == r_count_70_io_out ? io_r_170_b : _GEN_14469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14471 = 8'hab == r_count_70_io_out ? io_r_171_b : _GEN_14470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14472 = 8'hac == r_count_70_io_out ? io_r_172_b : _GEN_14471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14473 = 8'had == r_count_70_io_out ? io_r_173_b : _GEN_14472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14474 = 8'hae == r_count_70_io_out ? io_r_174_b : _GEN_14473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14475 = 8'haf == r_count_70_io_out ? io_r_175_b : _GEN_14474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14476 = 8'hb0 == r_count_70_io_out ? io_r_176_b : _GEN_14475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14477 = 8'hb1 == r_count_70_io_out ? io_r_177_b : _GEN_14476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14478 = 8'hb2 == r_count_70_io_out ? io_r_178_b : _GEN_14477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14479 = 8'hb3 == r_count_70_io_out ? io_r_179_b : _GEN_14478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14480 = 8'hb4 == r_count_70_io_out ? io_r_180_b : _GEN_14479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14481 = 8'hb5 == r_count_70_io_out ? io_r_181_b : _GEN_14480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14482 = 8'hb6 == r_count_70_io_out ? io_r_182_b : _GEN_14481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14483 = 8'hb7 == r_count_70_io_out ? io_r_183_b : _GEN_14482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14484 = 8'hb8 == r_count_70_io_out ? io_r_184_b : _GEN_14483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14485 = 8'hb9 == r_count_70_io_out ? io_r_185_b : _GEN_14484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14486 = 8'hba == r_count_70_io_out ? io_r_186_b : _GEN_14485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14487 = 8'hbb == r_count_70_io_out ? io_r_187_b : _GEN_14486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14488 = 8'hbc == r_count_70_io_out ? io_r_188_b : _GEN_14487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14489 = 8'hbd == r_count_70_io_out ? io_r_189_b : _GEN_14488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14490 = 8'hbe == r_count_70_io_out ? io_r_190_b : _GEN_14489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14491 = 8'hbf == r_count_70_io_out ? io_r_191_b : _GEN_14490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14492 = 8'hc0 == r_count_70_io_out ? io_r_192_b : _GEN_14491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14493 = 8'hc1 == r_count_70_io_out ? io_r_193_b : _GEN_14492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14494 = 8'hc2 == r_count_70_io_out ? io_r_194_b : _GEN_14493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14495 = 8'hc3 == r_count_70_io_out ? io_r_195_b : _GEN_14494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14496 = 8'hc4 == r_count_70_io_out ? io_r_196_b : _GEN_14495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14497 = 8'hc5 == r_count_70_io_out ? io_r_197_b : _GEN_14496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14498 = 8'hc6 == r_count_70_io_out ? io_r_198_b : _GEN_14497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14501 = 8'h1 == r_count_71_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14502 = 8'h2 == r_count_71_io_out ? io_r_2_b : _GEN_14501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14503 = 8'h3 == r_count_71_io_out ? io_r_3_b : _GEN_14502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14504 = 8'h4 == r_count_71_io_out ? io_r_4_b : _GEN_14503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14505 = 8'h5 == r_count_71_io_out ? io_r_5_b : _GEN_14504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14506 = 8'h6 == r_count_71_io_out ? io_r_6_b : _GEN_14505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14507 = 8'h7 == r_count_71_io_out ? io_r_7_b : _GEN_14506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14508 = 8'h8 == r_count_71_io_out ? io_r_8_b : _GEN_14507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14509 = 8'h9 == r_count_71_io_out ? io_r_9_b : _GEN_14508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14510 = 8'ha == r_count_71_io_out ? io_r_10_b : _GEN_14509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14511 = 8'hb == r_count_71_io_out ? io_r_11_b : _GEN_14510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14512 = 8'hc == r_count_71_io_out ? io_r_12_b : _GEN_14511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14513 = 8'hd == r_count_71_io_out ? io_r_13_b : _GEN_14512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14514 = 8'he == r_count_71_io_out ? io_r_14_b : _GEN_14513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14515 = 8'hf == r_count_71_io_out ? io_r_15_b : _GEN_14514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14516 = 8'h10 == r_count_71_io_out ? io_r_16_b : _GEN_14515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14517 = 8'h11 == r_count_71_io_out ? io_r_17_b : _GEN_14516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14518 = 8'h12 == r_count_71_io_out ? io_r_18_b : _GEN_14517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14519 = 8'h13 == r_count_71_io_out ? io_r_19_b : _GEN_14518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14520 = 8'h14 == r_count_71_io_out ? io_r_20_b : _GEN_14519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14521 = 8'h15 == r_count_71_io_out ? io_r_21_b : _GEN_14520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14522 = 8'h16 == r_count_71_io_out ? io_r_22_b : _GEN_14521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14523 = 8'h17 == r_count_71_io_out ? io_r_23_b : _GEN_14522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14524 = 8'h18 == r_count_71_io_out ? io_r_24_b : _GEN_14523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14525 = 8'h19 == r_count_71_io_out ? io_r_25_b : _GEN_14524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14526 = 8'h1a == r_count_71_io_out ? io_r_26_b : _GEN_14525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14527 = 8'h1b == r_count_71_io_out ? io_r_27_b : _GEN_14526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14528 = 8'h1c == r_count_71_io_out ? io_r_28_b : _GEN_14527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14529 = 8'h1d == r_count_71_io_out ? io_r_29_b : _GEN_14528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14530 = 8'h1e == r_count_71_io_out ? io_r_30_b : _GEN_14529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14531 = 8'h1f == r_count_71_io_out ? io_r_31_b : _GEN_14530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14532 = 8'h20 == r_count_71_io_out ? io_r_32_b : _GEN_14531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14533 = 8'h21 == r_count_71_io_out ? io_r_33_b : _GEN_14532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14534 = 8'h22 == r_count_71_io_out ? io_r_34_b : _GEN_14533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14535 = 8'h23 == r_count_71_io_out ? io_r_35_b : _GEN_14534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14536 = 8'h24 == r_count_71_io_out ? io_r_36_b : _GEN_14535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14537 = 8'h25 == r_count_71_io_out ? io_r_37_b : _GEN_14536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14538 = 8'h26 == r_count_71_io_out ? io_r_38_b : _GEN_14537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14539 = 8'h27 == r_count_71_io_out ? io_r_39_b : _GEN_14538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14540 = 8'h28 == r_count_71_io_out ? io_r_40_b : _GEN_14539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14541 = 8'h29 == r_count_71_io_out ? io_r_41_b : _GEN_14540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14542 = 8'h2a == r_count_71_io_out ? io_r_42_b : _GEN_14541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14543 = 8'h2b == r_count_71_io_out ? io_r_43_b : _GEN_14542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14544 = 8'h2c == r_count_71_io_out ? io_r_44_b : _GEN_14543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14545 = 8'h2d == r_count_71_io_out ? io_r_45_b : _GEN_14544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14546 = 8'h2e == r_count_71_io_out ? io_r_46_b : _GEN_14545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14547 = 8'h2f == r_count_71_io_out ? io_r_47_b : _GEN_14546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14548 = 8'h30 == r_count_71_io_out ? io_r_48_b : _GEN_14547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14549 = 8'h31 == r_count_71_io_out ? io_r_49_b : _GEN_14548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14550 = 8'h32 == r_count_71_io_out ? io_r_50_b : _GEN_14549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14551 = 8'h33 == r_count_71_io_out ? io_r_51_b : _GEN_14550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14552 = 8'h34 == r_count_71_io_out ? io_r_52_b : _GEN_14551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14553 = 8'h35 == r_count_71_io_out ? io_r_53_b : _GEN_14552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14554 = 8'h36 == r_count_71_io_out ? io_r_54_b : _GEN_14553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14555 = 8'h37 == r_count_71_io_out ? io_r_55_b : _GEN_14554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14556 = 8'h38 == r_count_71_io_out ? io_r_56_b : _GEN_14555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14557 = 8'h39 == r_count_71_io_out ? io_r_57_b : _GEN_14556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14558 = 8'h3a == r_count_71_io_out ? io_r_58_b : _GEN_14557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14559 = 8'h3b == r_count_71_io_out ? io_r_59_b : _GEN_14558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14560 = 8'h3c == r_count_71_io_out ? io_r_60_b : _GEN_14559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14561 = 8'h3d == r_count_71_io_out ? io_r_61_b : _GEN_14560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14562 = 8'h3e == r_count_71_io_out ? io_r_62_b : _GEN_14561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14563 = 8'h3f == r_count_71_io_out ? io_r_63_b : _GEN_14562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14564 = 8'h40 == r_count_71_io_out ? io_r_64_b : _GEN_14563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14565 = 8'h41 == r_count_71_io_out ? io_r_65_b : _GEN_14564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14566 = 8'h42 == r_count_71_io_out ? io_r_66_b : _GEN_14565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14567 = 8'h43 == r_count_71_io_out ? io_r_67_b : _GEN_14566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14568 = 8'h44 == r_count_71_io_out ? io_r_68_b : _GEN_14567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14569 = 8'h45 == r_count_71_io_out ? io_r_69_b : _GEN_14568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14570 = 8'h46 == r_count_71_io_out ? io_r_70_b : _GEN_14569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14571 = 8'h47 == r_count_71_io_out ? io_r_71_b : _GEN_14570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14572 = 8'h48 == r_count_71_io_out ? io_r_72_b : _GEN_14571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14573 = 8'h49 == r_count_71_io_out ? io_r_73_b : _GEN_14572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14574 = 8'h4a == r_count_71_io_out ? io_r_74_b : _GEN_14573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14575 = 8'h4b == r_count_71_io_out ? io_r_75_b : _GEN_14574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14576 = 8'h4c == r_count_71_io_out ? io_r_76_b : _GEN_14575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14577 = 8'h4d == r_count_71_io_out ? io_r_77_b : _GEN_14576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14578 = 8'h4e == r_count_71_io_out ? io_r_78_b : _GEN_14577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14579 = 8'h4f == r_count_71_io_out ? io_r_79_b : _GEN_14578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14580 = 8'h50 == r_count_71_io_out ? io_r_80_b : _GEN_14579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14581 = 8'h51 == r_count_71_io_out ? io_r_81_b : _GEN_14580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14582 = 8'h52 == r_count_71_io_out ? io_r_82_b : _GEN_14581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14583 = 8'h53 == r_count_71_io_out ? io_r_83_b : _GEN_14582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14584 = 8'h54 == r_count_71_io_out ? io_r_84_b : _GEN_14583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14585 = 8'h55 == r_count_71_io_out ? io_r_85_b : _GEN_14584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14586 = 8'h56 == r_count_71_io_out ? io_r_86_b : _GEN_14585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14587 = 8'h57 == r_count_71_io_out ? io_r_87_b : _GEN_14586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14588 = 8'h58 == r_count_71_io_out ? io_r_88_b : _GEN_14587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14589 = 8'h59 == r_count_71_io_out ? io_r_89_b : _GEN_14588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14590 = 8'h5a == r_count_71_io_out ? io_r_90_b : _GEN_14589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14591 = 8'h5b == r_count_71_io_out ? io_r_91_b : _GEN_14590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14592 = 8'h5c == r_count_71_io_out ? io_r_92_b : _GEN_14591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14593 = 8'h5d == r_count_71_io_out ? io_r_93_b : _GEN_14592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14594 = 8'h5e == r_count_71_io_out ? io_r_94_b : _GEN_14593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14595 = 8'h5f == r_count_71_io_out ? io_r_95_b : _GEN_14594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14596 = 8'h60 == r_count_71_io_out ? io_r_96_b : _GEN_14595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14597 = 8'h61 == r_count_71_io_out ? io_r_97_b : _GEN_14596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14598 = 8'h62 == r_count_71_io_out ? io_r_98_b : _GEN_14597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14599 = 8'h63 == r_count_71_io_out ? io_r_99_b : _GEN_14598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14600 = 8'h64 == r_count_71_io_out ? io_r_100_b : _GEN_14599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14601 = 8'h65 == r_count_71_io_out ? io_r_101_b : _GEN_14600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14602 = 8'h66 == r_count_71_io_out ? io_r_102_b : _GEN_14601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14603 = 8'h67 == r_count_71_io_out ? io_r_103_b : _GEN_14602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14604 = 8'h68 == r_count_71_io_out ? io_r_104_b : _GEN_14603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14605 = 8'h69 == r_count_71_io_out ? io_r_105_b : _GEN_14604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14606 = 8'h6a == r_count_71_io_out ? io_r_106_b : _GEN_14605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14607 = 8'h6b == r_count_71_io_out ? io_r_107_b : _GEN_14606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14608 = 8'h6c == r_count_71_io_out ? io_r_108_b : _GEN_14607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14609 = 8'h6d == r_count_71_io_out ? io_r_109_b : _GEN_14608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14610 = 8'h6e == r_count_71_io_out ? io_r_110_b : _GEN_14609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14611 = 8'h6f == r_count_71_io_out ? io_r_111_b : _GEN_14610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14612 = 8'h70 == r_count_71_io_out ? io_r_112_b : _GEN_14611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14613 = 8'h71 == r_count_71_io_out ? io_r_113_b : _GEN_14612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14614 = 8'h72 == r_count_71_io_out ? io_r_114_b : _GEN_14613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14615 = 8'h73 == r_count_71_io_out ? io_r_115_b : _GEN_14614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14616 = 8'h74 == r_count_71_io_out ? io_r_116_b : _GEN_14615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14617 = 8'h75 == r_count_71_io_out ? io_r_117_b : _GEN_14616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14618 = 8'h76 == r_count_71_io_out ? io_r_118_b : _GEN_14617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14619 = 8'h77 == r_count_71_io_out ? io_r_119_b : _GEN_14618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14620 = 8'h78 == r_count_71_io_out ? io_r_120_b : _GEN_14619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14621 = 8'h79 == r_count_71_io_out ? io_r_121_b : _GEN_14620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14622 = 8'h7a == r_count_71_io_out ? io_r_122_b : _GEN_14621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14623 = 8'h7b == r_count_71_io_out ? io_r_123_b : _GEN_14622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14624 = 8'h7c == r_count_71_io_out ? io_r_124_b : _GEN_14623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14625 = 8'h7d == r_count_71_io_out ? io_r_125_b : _GEN_14624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14626 = 8'h7e == r_count_71_io_out ? io_r_126_b : _GEN_14625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14627 = 8'h7f == r_count_71_io_out ? io_r_127_b : _GEN_14626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14628 = 8'h80 == r_count_71_io_out ? io_r_128_b : _GEN_14627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14629 = 8'h81 == r_count_71_io_out ? io_r_129_b : _GEN_14628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14630 = 8'h82 == r_count_71_io_out ? io_r_130_b : _GEN_14629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14631 = 8'h83 == r_count_71_io_out ? io_r_131_b : _GEN_14630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14632 = 8'h84 == r_count_71_io_out ? io_r_132_b : _GEN_14631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14633 = 8'h85 == r_count_71_io_out ? io_r_133_b : _GEN_14632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14634 = 8'h86 == r_count_71_io_out ? io_r_134_b : _GEN_14633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14635 = 8'h87 == r_count_71_io_out ? io_r_135_b : _GEN_14634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14636 = 8'h88 == r_count_71_io_out ? io_r_136_b : _GEN_14635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14637 = 8'h89 == r_count_71_io_out ? io_r_137_b : _GEN_14636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14638 = 8'h8a == r_count_71_io_out ? io_r_138_b : _GEN_14637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14639 = 8'h8b == r_count_71_io_out ? io_r_139_b : _GEN_14638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14640 = 8'h8c == r_count_71_io_out ? io_r_140_b : _GEN_14639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14641 = 8'h8d == r_count_71_io_out ? io_r_141_b : _GEN_14640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14642 = 8'h8e == r_count_71_io_out ? io_r_142_b : _GEN_14641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14643 = 8'h8f == r_count_71_io_out ? io_r_143_b : _GEN_14642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14644 = 8'h90 == r_count_71_io_out ? io_r_144_b : _GEN_14643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14645 = 8'h91 == r_count_71_io_out ? io_r_145_b : _GEN_14644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14646 = 8'h92 == r_count_71_io_out ? io_r_146_b : _GEN_14645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14647 = 8'h93 == r_count_71_io_out ? io_r_147_b : _GEN_14646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14648 = 8'h94 == r_count_71_io_out ? io_r_148_b : _GEN_14647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14649 = 8'h95 == r_count_71_io_out ? io_r_149_b : _GEN_14648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14650 = 8'h96 == r_count_71_io_out ? io_r_150_b : _GEN_14649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14651 = 8'h97 == r_count_71_io_out ? io_r_151_b : _GEN_14650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14652 = 8'h98 == r_count_71_io_out ? io_r_152_b : _GEN_14651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14653 = 8'h99 == r_count_71_io_out ? io_r_153_b : _GEN_14652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14654 = 8'h9a == r_count_71_io_out ? io_r_154_b : _GEN_14653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14655 = 8'h9b == r_count_71_io_out ? io_r_155_b : _GEN_14654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14656 = 8'h9c == r_count_71_io_out ? io_r_156_b : _GEN_14655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14657 = 8'h9d == r_count_71_io_out ? io_r_157_b : _GEN_14656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14658 = 8'h9e == r_count_71_io_out ? io_r_158_b : _GEN_14657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14659 = 8'h9f == r_count_71_io_out ? io_r_159_b : _GEN_14658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14660 = 8'ha0 == r_count_71_io_out ? io_r_160_b : _GEN_14659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14661 = 8'ha1 == r_count_71_io_out ? io_r_161_b : _GEN_14660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14662 = 8'ha2 == r_count_71_io_out ? io_r_162_b : _GEN_14661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14663 = 8'ha3 == r_count_71_io_out ? io_r_163_b : _GEN_14662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14664 = 8'ha4 == r_count_71_io_out ? io_r_164_b : _GEN_14663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14665 = 8'ha5 == r_count_71_io_out ? io_r_165_b : _GEN_14664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14666 = 8'ha6 == r_count_71_io_out ? io_r_166_b : _GEN_14665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14667 = 8'ha7 == r_count_71_io_out ? io_r_167_b : _GEN_14666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14668 = 8'ha8 == r_count_71_io_out ? io_r_168_b : _GEN_14667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14669 = 8'ha9 == r_count_71_io_out ? io_r_169_b : _GEN_14668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14670 = 8'haa == r_count_71_io_out ? io_r_170_b : _GEN_14669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14671 = 8'hab == r_count_71_io_out ? io_r_171_b : _GEN_14670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14672 = 8'hac == r_count_71_io_out ? io_r_172_b : _GEN_14671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14673 = 8'had == r_count_71_io_out ? io_r_173_b : _GEN_14672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14674 = 8'hae == r_count_71_io_out ? io_r_174_b : _GEN_14673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14675 = 8'haf == r_count_71_io_out ? io_r_175_b : _GEN_14674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14676 = 8'hb0 == r_count_71_io_out ? io_r_176_b : _GEN_14675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14677 = 8'hb1 == r_count_71_io_out ? io_r_177_b : _GEN_14676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14678 = 8'hb2 == r_count_71_io_out ? io_r_178_b : _GEN_14677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14679 = 8'hb3 == r_count_71_io_out ? io_r_179_b : _GEN_14678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14680 = 8'hb4 == r_count_71_io_out ? io_r_180_b : _GEN_14679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14681 = 8'hb5 == r_count_71_io_out ? io_r_181_b : _GEN_14680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14682 = 8'hb6 == r_count_71_io_out ? io_r_182_b : _GEN_14681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14683 = 8'hb7 == r_count_71_io_out ? io_r_183_b : _GEN_14682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14684 = 8'hb8 == r_count_71_io_out ? io_r_184_b : _GEN_14683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14685 = 8'hb9 == r_count_71_io_out ? io_r_185_b : _GEN_14684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14686 = 8'hba == r_count_71_io_out ? io_r_186_b : _GEN_14685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14687 = 8'hbb == r_count_71_io_out ? io_r_187_b : _GEN_14686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14688 = 8'hbc == r_count_71_io_out ? io_r_188_b : _GEN_14687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14689 = 8'hbd == r_count_71_io_out ? io_r_189_b : _GEN_14688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14690 = 8'hbe == r_count_71_io_out ? io_r_190_b : _GEN_14689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14691 = 8'hbf == r_count_71_io_out ? io_r_191_b : _GEN_14690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14692 = 8'hc0 == r_count_71_io_out ? io_r_192_b : _GEN_14691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14693 = 8'hc1 == r_count_71_io_out ? io_r_193_b : _GEN_14692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14694 = 8'hc2 == r_count_71_io_out ? io_r_194_b : _GEN_14693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14695 = 8'hc3 == r_count_71_io_out ? io_r_195_b : _GEN_14694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14696 = 8'hc4 == r_count_71_io_out ? io_r_196_b : _GEN_14695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14697 = 8'hc5 == r_count_71_io_out ? io_r_197_b : _GEN_14696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14698 = 8'hc6 == r_count_71_io_out ? io_r_198_b : _GEN_14697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14701 = 8'h1 == r_count_72_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14702 = 8'h2 == r_count_72_io_out ? io_r_2_b : _GEN_14701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14703 = 8'h3 == r_count_72_io_out ? io_r_3_b : _GEN_14702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14704 = 8'h4 == r_count_72_io_out ? io_r_4_b : _GEN_14703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14705 = 8'h5 == r_count_72_io_out ? io_r_5_b : _GEN_14704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14706 = 8'h6 == r_count_72_io_out ? io_r_6_b : _GEN_14705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14707 = 8'h7 == r_count_72_io_out ? io_r_7_b : _GEN_14706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14708 = 8'h8 == r_count_72_io_out ? io_r_8_b : _GEN_14707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14709 = 8'h9 == r_count_72_io_out ? io_r_9_b : _GEN_14708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14710 = 8'ha == r_count_72_io_out ? io_r_10_b : _GEN_14709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14711 = 8'hb == r_count_72_io_out ? io_r_11_b : _GEN_14710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14712 = 8'hc == r_count_72_io_out ? io_r_12_b : _GEN_14711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14713 = 8'hd == r_count_72_io_out ? io_r_13_b : _GEN_14712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14714 = 8'he == r_count_72_io_out ? io_r_14_b : _GEN_14713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14715 = 8'hf == r_count_72_io_out ? io_r_15_b : _GEN_14714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14716 = 8'h10 == r_count_72_io_out ? io_r_16_b : _GEN_14715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14717 = 8'h11 == r_count_72_io_out ? io_r_17_b : _GEN_14716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14718 = 8'h12 == r_count_72_io_out ? io_r_18_b : _GEN_14717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14719 = 8'h13 == r_count_72_io_out ? io_r_19_b : _GEN_14718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14720 = 8'h14 == r_count_72_io_out ? io_r_20_b : _GEN_14719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14721 = 8'h15 == r_count_72_io_out ? io_r_21_b : _GEN_14720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14722 = 8'h16 == r_count_72_io_out ? io_r_22_b : _GEN_14721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14723 = 8'h17 == r_count_72_io_out ? io_r_23_b : _GEN_14722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14724 = 8'h18 == r_count_72_io_out ? io_r_24_b : _GEN_14723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14725 = 8'h19 == r_count_72_io_out ? io_r_25_b : _GEN_14724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14726 = 8'h1a == r_count_72_io_out ? io_r_26_b : _GEN_14725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14727 = 8'h1b == r_count_72_io_out ? io_r_27_b : _GEN_14726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14728 = 8'h1c == r_count_72_io_out ? io_r_28_b : _GEN_14727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14729 = 8'h1d == r_count_72_io_out ? io_r_29_b : _GEN_14728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14730 = 8'h1e == r_count_72_io_out ? io_r_30_b : _GEN_14729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14731 = 8'h1f == r_count_72_io_out ? io_r_31_b : _GEN_14730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14732 = 8'h20 == r_count_72_io_out ? io_r_32_b : _GEN_14731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14733 = 8'h21 == r_count_72_io_out ? io_r_33_b : _GEN_14732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14734 = 8'h22 == r_count_72_io_out ? io_r_34_b : _GEN_14733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14735 = 8'h23 == r_count_72_io_out ? io_r_35_b : _GEN_14734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14736 = 8'h24 == r_count_72_io_out ? io_r_36_b : _GEN_14735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14737 = 8'h25 == r_count_72_io_out ? io_r_37_b : _GEN_14736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14738 = 8'h26 == r_count_72_io_out ? io_r_38_b : _GEN_14737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14739 = 8'h27 == r_count_72_io_out ? io_r_39_b : _GEN_14738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14740 = 8'h28 == r_count_72_io_out ? io_r_40_b : _GEN_14739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14741 = 8'h29 == r_count_72_io_out ? io_r_41_b : _GEN_14740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14742 = 8'h2a == r_count_72_io_out ? io_r_42_b : _GEN_14741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14743 = 8'h2b == r_count_72_io_out ? io_r_43_b : _GEN_14742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14744 = 8'h2c == r_count_72_io_out ? io_r_44_b : _GEN_14743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14745 = 8'h2d == r_count_72_io_out ? io_r_45_b : _GEN_14744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14746 = 8'h2e == r_count_72_io_out ? io_r_46_b : _GEN_14745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14747 = 8'h2f == r_count_72_io_out ? io_r_47_b : _GEN_14746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14748 = 8'h30 == r_count_72_io_out ? io_r_48_b : _GEN_14747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14749 = 8'h31 == r_count_72_io_out ? io_r_49_b : _GEN_14748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14750 = 8'h32 == r_count_72_io_out ? io_r_50_b : _GEN_14749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14751 = 8'h33 == r_count_72_io_out ? io_r_51_b : _GEN_14750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14752 = 8'h34 == r_count_72_io_out ? io_r_52_b : _GEN_14751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14753 = 8'h35 == r_count_72_io_out ? io_r_53_b : _GEN_14752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14754 = 8'h36 == r_count_72_io_out ? io_r_54_b : _GEN_14753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14755 = 8'h37 == r_count_72_io_out ? io_r_55_b : _GEN_14754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14756 = 8'h38 == r_count_72_io_out ? io_r_56_b : _GEN_14755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14757 = 8'h39 == r_count_72_io_out ? io_r_57_b : _GEN_14756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14758 = 8'h3a == r_count_72_io_out ? io_r_58_b : _GEN_14757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14759 = 8'h3b == r_count_72_io_out ? io_r_59_b : _GEN_14758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14760 = 8'h3c == r_count_72_io_out ? io_r_60_b : _GEN_14759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14761 = 8'h3d == r_count_72_io_out ? io_r_61_b : _GEN_14760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14762 = 8'h3e == r_count_72_io_out ? io_r_62_b : _GEN_14761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14763 = 8'h3f == r_count_72_io_out ? io_r_63_b : _GEN_14762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14764 = 8'h40 == r_count_72_io_out ? io_r_64_b : _GEN_14763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14765 = 8'h41 == r_count_72_io_out ? io_r_65_b : _GEN_14764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14766 = 8'h42 == r_count_72_io_out ? io_r_66_b : _GEN_14765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14767 = 8'h43 == r_count_72_io_out ? io_r_67_b : _GEN_14766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14768 = 8'h44 == r_count_72_io_out ? io_r_68_b : _GEN_14767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14769 = 8'h45 == r_count_72_io_out ? io_r_69_b : _GEN_14768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14770 = 8'h46 == r_count_72_io_out ? io_r_70_b : _GEN_14769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14771 = 8'h47 == r_count_72_io_out ? io_r_71_b : _GEN_14770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14772 = 8'h48 == r_count_72_io_out ? io_r_72_b : _GEN_14771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14773 = 8'h49 == r_count_72_io_out ? io_r_73_b : _GEN_14772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14774 = 8'h4a == r_count_72_io_out ? io_r_74_b : _GEN_14773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14775 = 8'h4b == r_count_72_io_out ? io_r_75_b : _GEN_14774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14776 = 8'h4c == r_count_72_io_out ? io_r_76_b : _GEN_14775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14777 = 8'h4d == r_count_72_io_out ? io_r_77_b : _GEN_14776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14778 = 8'h4e == r_count_72_io_out ? io_r_78_b : _GEN_14777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14779 = 8'h4f == r_count_72_io_out ? io_r_79_b : _GEN_14778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14780 = 8'h50 == r_count_72_io_out ? io_r_80_b : _GEN_14779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14781 = 8'h51 == r_count_72_io_out ? io_r_81_b : _GEN_14780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14782 = 8'h52 == r_count_72_io_out ? io_r_82_b : _GEN_14781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14783 = 8'h53 == r_count_72_io_out ? io_r_83_b : _GEN_14782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14784 = 8'h54 == r_count_72_io_out ? io_r_84_b : _GEN_14783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14785 = 8'h55 == r_count_72_io_out ? io_r_85_b : _GEN_14784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14786 = 8'h56 == r_count_72_io_out ? io_r_86_b : _GEN_14785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14787 = 8'h57 == r_count_72_io_out ? io_r_87_b : _GEN_14786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14788 = 8'h58 == r_count_72_io_out ? io_r_88_b : _GEN_14787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14789 = 8'h59 == r_count_72_io_out ? io_r_89_b : _GEN_14788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14790 = 8'h5a == r_count_72_io_out ? io_r_90_b : _GEN_14789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14791 = 8'h5b == r_count_72_io_out ? io_r_91_b : _GEN_14790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14792 = 8'h5c == r_count_72_io_out ? io_r_92_b : _GEN_14791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14793 = 8'h5d == r_count_72_io_out ? io_r_93_b : _GEN_14792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14794 = 8'h5e == r_count_72_io_out ? io_r_94_b : _GEN_14793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14795 = 8'h5f == r_count_72_io_out ? io_r_95_b : _GEN_14794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14796 = 8'h60 == r_count_72_io_out ? io_r_96_b : _GEN_14795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14797 = 8'h61 == r_count_72_io_out ? io_r_97_b : _GEN_14796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14798 = 8'h62 == r_count_72_io_out ? io_r_98_b : _GEN_14797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14799 = 8'h63 == r_count_72_io_out ? io_r_99_b : _GEN_14798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14800 = 8'h64 == r_count_72_io_out ? io_r_100_b : _GEN_14799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14801 = 8'h65 == r_count_72_io_out ? io_r_101_b : _GEN_14800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14802 = 8'h66 == r_count_72_io_out ? io_r_102_b : _GEN_14801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14803 = 8'h67 == r_count_72_io_out ? io_r_103_b : _GEN_14802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14804 = 8'h68 == r_count_72_io_out ? io_r_104_b : _GEN_14803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14805 = 8'h69 == r_count_72_io_out ? io_r_105_b : _GEN_14804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14806 = 8'h6a == r_count_72_io_out ? io_r_106_b : _GEN_14805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14807 = 8'h6b == r_count_72_io_out ? io_r_107_b : _GEN_14806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14808 = 8'h6c == r_count_72_io_out ? io_r_108_b : _GEN_14807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14809 = 8'h6d == r_count_72_io_out ? io_r_109_b : _GEN_14808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14810 = 8'h6e == r_count_72_io_out ? io_r_110_b : _GEN_14809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14811 = 8'h6f == r_count_72_io_out ? io_r_111_b : _GEN_14810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14812 = 8'h70 == r_count_72_io_out ? io_r_112_b : _GEN_14811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14813 = 8'h71 == r_count_72_io_out ? io_r_113_b : _GEN_14812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14814 = 8'h72 == r_count_72_io_out ? io_r_114_b : _GEN_14813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14815 = 8'h73 == r_count_72_io_out ? io_r_115_b : _GEN_14814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14816 = 8'h74 == r_count_72_io_out ? io_r_116_b : _GEN_14815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14817 = 8'h75 == r_count_72_io_out ? io_r_117_b : _GEN_14816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14818 = 8'h76 == r_count_72_io_out ? io_r_118_b : _GEN_14817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14819 = 8'h77 == r_count_72_io_out ? io_r_119_b : _GEN_14818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14820 = 8'h78 == r_count_72_io_out ? io_r_120_b : _GEN_14819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14821 = 8'h79 == r_count_72_io_out ? io_r_121_b : _GEN_14820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14822 = 8'h7a == r_count_72_io_out ? io_r_122_b : _GEN_14821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14823 = 8'h7b == r_count_72_io_out ? io_r_123_b : _GEN_14822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14824 = 8'h7c == r_count_72_io_out ? io_r_124_b : _GEN_14823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14825 = 8'h7d == r_count_72_io_out ? io_r_125_b : _GEN_14824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14826 = 8'h7e == r_count_72_io_out ? io_r_126_b : _GEN_14825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14827 = 8'h7f == r_count_72_io_out ? io_r_127_b : _GEN_14826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14828 = 8'h80 == r_count_72_io_out ? io_r_128_b : _GEN_14827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14829 = 8'h81 == r_count_72_io_out ? io_r_129_b : _GEN_14828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14830 = 8'h82 == r_count_72_io_out ? io_r_130_b : _GEN_14829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14831 = 8'h83 == r_count_72_io_out ? io_r_131_b : _GEN_14830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14832 = 8'h84 == r_count_72_io_out ? io_r_132_b : _GEN_14831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14833 = 8'h85 == r_count_72_io_out ? io_r_133_b : _GEN_14832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14834 = 8'h86 == r_count_72_io_out ? io_r_134_b : _GEN_14833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14835 = 8'h87 == r_count_72_io_out ? io_r_135_b : _GEN_14834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14836 = 8'h88 == r_count_72_io_out ? io_r_136_b : _GEN_14835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14837 = 8'h89 == r_count_72_io_out ? io_r_137_b : _GEN_14836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14838 = 8'h8a == r_count_72_io_out ? io_r_138_b : _GEN_14837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14839 = 8'h8b == r_count_72_io_out ? io_r_139_b : _GEN_14838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14840 = 8'h8c == r_count_72_io_out ? io_r_140_b : _GEN_14839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14841 = 8'h8d == r_count_72_io_out ? io_r_141_b : _GEN_14840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14842 = 8'h8e == r_count_72_io_out ? io_r_142_b : _GEN_14841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14843 = 8'h8f == r_count_72_io_out ? io_r_143_b : _GEN_14842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14844 = 8'h90 == r_count_72_io_out ? io_r_144_b : _GEN_14843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14845 = 8'h91 == r_count_72_io_out ? io_r_145_b : _GEN_14844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14846 = 8'h92 == r_count_72_io_out ? io_r_146_b : _GEN_14845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14847 = 8'h93 == r_count_72_io_out ? io_r_147_b : _GEN_14846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14848 = 8'h94 == r_count_72_io_out ? io_r_148_b : _GEN_14847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14849 = 8'h95 == r_count_72_io_out ? io_r_149_b : _GEN_14848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14850 = 8'h96 == r_count_72_io_out ? io_r_150_b : _GEN_14849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14851 = 8'h97 == r_count_72_io_out ? io_r_151_b : _GEN_14850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14852 = 8'h98 == r_count_72_io_out ? io_r_152_b : _GEN_14851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14853 = 8'h99 == r_count_72_io_out ? io_r_153_b : _GEN_14852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14854 = 8'h9a == r_count_72_io_out ? io_r_154_b : _GEN_14853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14855 = 8'h9b == r_count_72_io_out ? io_r_155_b : _GEN_14854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14856 = 8'h9c == r_count_72_io_out ? io_r_156_b : _GEN_14855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14857 = 8'h9d == r_count_72_io_out ? io_r_157_b : _GEN_14856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14858 = 8'h9e == r_count_72_io_out ? io_r_158_b : _GEN_14857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14859 = 8'h9f == r_count_72_io_out ? io_r_159_b : _GEN_14858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14860 = 8'ha0 == r_count_72_io_out ? io_r_160_b : _GEN_14859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14861 = 8'ha1 == r_count_72_io_out ? io_r_161_b : _GEN_14860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14862 = 8'ha2 == r_count_72_io_out ? io_r_162_b : _GEN_14861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14863 = 8'ha3 == r_count_72_io_out ? io_r_163_b : _GEN_14862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14864 = 8'ha4 == r_count_72_io_out ? io_r_164_b : _GEN_14863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14865 = 8'ha5 == r_count_72_io_out ? io_r_165_b : _GEN_14864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14866 = 8'ha6 == r_count_72_io_out ? io_r_166_b : _GEN_14865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14867 = 8'ha7 == r_count_72_io_out ? io_r_167_b : _GEN_14866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14868 = 8'ha8 == r_count_72_io_out ? io_r_168_b : _GEN_14867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14869 = 8'ha9 == r_count_72_io_out ? io_r_169_b : _GEN_14868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14870 = 8'haa == r_count_72_io_out ? io_r_170_b : _GEN_14869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14871 = 8'hab == r_count_72_io_out ? io_r_171_b : _GEN_14870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14872 = 8'hac == r_count_72_io_out ? io_r_172_b : _GEN_14871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14873 = 8'had == r_count_72_io_out ? io_r_173_b : _GEN_14872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14874 = 8'hae == r_count_72_io_out ? io_r_174_b : _GEN_14873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14875 = 8'haf == r_count_72_io_out ? io_r_175_b : _GEN_14874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14876 = 8'hb0 == r_count_72_io_out ? io_r_176_b : _GEN_14875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14877 = 8'hb1 == r_count_72_io_out ? io_r_177_b : _GEN_14876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14878 = 8'hb2 == r_count_72_io_out ? io_r_178_b : _GEN_14877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14879 = 8'hb3 == r_count_72_io_out ? io_r_179_b : _GEN_14878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14880 = 8'hb4 == r_count_72_io_out ? io_r_180_b : _GEN_14879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14881 = 8'hb5 == r_count_72_io_out ? io_r_181_b : _GEN_14880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14882 = 8'hb6 == r_count_72_io_out ? io_r_182_b : _GEN_14881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14883 = 8'hb7 == r_count_72_io_out ? io_r_183_b : _GEN_14882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14884 = 8'hb8 == r_count_72_io_out ? io_r_184_b : _GEN_14883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14885 = 8'hb9 == r_count_72_io_out ? io_r_185_b : _GEN_14884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14886 = 8'hba == r_count_72_io_out ? io_r_186_b : _GEN_14885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14887 = 8'hbb == r_count_72_io_out ? io_r_187_b : _GEN_14886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14888 = 8'hbc == r_count_72_io_out ? io_r_188_b : _GEN_14887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14889 = 8'hbd == r_count_72_io_out ? io_r_189_b : _GEN_14888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14890 = 8'hbe == r_count_72_io_out ? io_r_190_b : _GEN_14889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14891 = 8'hbf == r_count_72_io_out ? io_r_191_b : _GEN_14890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14892 = 8'hc0 == r_count_72_io_out ? io_r_192_b : _GEN_14891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14893 = 8'hc1 == r_count_72_io_out ? io_r_193_b : _GEN_14892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14894 = 8'hc2 == r_count_72_io_out ? io_r_194_b : _GEN_14893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14895 = 8'hc3 == r_count_72_io_out ? io_r_195_b : _GEN_14894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14896 = 8'hc4 == r_count_72_io_out ? io_r_196_b : _GEN_14895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14897 = 8'hc5 == r_count_72_io_out ? io_r_197_b : _GEN_14896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14898 = 8'hc6 == r_count_72_io_out ? io_r_198_b : _GEN_14897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14901 = 8'h1 == r_count_73_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14902 = 8'h2 == r_count_73_io_out ? io_r_2_b : _GEN_14901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14903 = 8'h3 == r_count_73_io_out ? io_r_3_b : _GEN_14902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14904 = 8'h4 == r_count_73_io_out ? io_r_4_b : _GEN_14903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14905 = 8'h5 == r_count_73_io_out ? io_r_5_b : _GEN_14904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14906 = 8'h6 == r_count_73_io_out ? io_r_6_b : _GEN_14905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14907 = 8'h7 == r_count_73_io_out ? io_r_7_b : _GEN_14906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14908 = 8'h8 == r_count_73_io_out ? io_r_8_b : _GEN_14907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14909 = 8'h9 == r_count_73_io_out ? io_r_9_b : _GEN_14908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14910 = 8'ha == r_count_73_io_out ? io_r_10_b : _GEN_14909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14911 = 8'hb == r_count_73_io_out ? io_r_11_b : _GEN_14910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14912 = 8'hc == r_count_73_io_out ? io_r_12_b : _GEN_14911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14913 = 8'hd == r_count_73_io_out ? io_r_13_b : _GEN_14912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14914 = 8'he == r_count_73_io_out ? io_r_14_b : _GEN_14913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14915 = 8'hf == r_count_73_io_out ? io_r_15_b : _GEN_14914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14916 = 8'h10 == r_count_73_io_out ? io_r_16_b : _GEN_14915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14917 = 8'h11 == r_count_73_io_out ? io_r_17_b : _GEN_14916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14918 = 8'h12 == r_count_73_io_out ? io_r_18_b : _GEN_14917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14919 = 8'h13 == r_count_73_io_out ? io_r_19_b : _GEN_14918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14920 = 8'h14 == r_count_73_io_out ? io_r_20_b : _GEN_14919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14921 = 8'h15 == r_count_73_io_out ? io_r_21_b : _GEN_14920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14922 = 8'h16 == r_count_73_io_out ? io_r_22_b : _GEN_14921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14923 = 8'h17 == r_count_73_io_out ? io_r_23_b : _GEN_14922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14924 = 8'h18 == r_count_73_io_out ? io_r_24_b : _GEN_14923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14925 = 8'h19 == r_count_73_io_out ? io_r_25_b : _GEN_14924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14926 = 8'h1a == r_count_73_io_out ? io_r_26_b : _GEN_14925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14927 = 8'h1b == r_count_73_io_out ? io_r_27_b : _GEN_14926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14928 = 8'h1c == r_count_73_io_out ? io_r_28_b : _GEN_14927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14929 = 8'h1d == r_count_73_io_out ? io_r_29_b : _GEN_14928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14930 = 8'h1e == r_count_73_io_out ? io_r_30_b : _GEN_14929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14931 = 8'h1f == r_count_73_io_out ? io_r_31_b : _GEN_14930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14932 = 8'h20 == r_count_73_io_out ? io_r_32_b : _GEN_14931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14933 = 8'h21 == r_count_73_io_out ? io_r_33_b : _GEN_14932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14934 = 8'h22 == r_count_73_io_out ? io_r_34_b : _GEN_14933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14935 = 8'h23 == r_count_73_io_out ? io_r_35_b : _GEN_14934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14936 = 8'h24 == r_count_73_io_out ? io_r_36_b : _GEN_14935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14937 = 8'h25 == r_count_73_io_out ? io_r_37_b : _GEN_14936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14938 = 8'h26 == r_count_73_io_out ? io_r_38_b : _GEN_14937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14939 = 8'h27 == r_count_73_io_out ? io_r_39_b : _GEN_14938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14940 = 8'h28 == r_count_73_io_out ? io_r_40_b : _GEN_14939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14941 = 8'h29 == r_count_73_io_out ? io_r_41_b : _GEN_14940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14942 = 8'h2a == r_count_73_io_out ? io_r_42_b : _GEN_14941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14943 = 8'h2b == r_count_73_io_out ? io_r_43_b : _GEN_14942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14944 = 8'h2c == r_count_73_io_out ? io_r_44_b : _GEN_14943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14945 = 8'h2d == r_count_73_io_out ? io_r_45_b : _GEN_14944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14946 = 8'h2e == r_count_73_io_out ? io_r_46_b : _GEN_14945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14947 = 8'h2f == r_count_73_io_out ? io_r_47_b : _GEN_14946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14948 = 8'h30 == r_count_73_io_out ? io_r_48_b : _GEN_14947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14949 = 8'h31 == r_count_73_io_out ? io_r_49_b : _GEN_14948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14950 = 8'h32 == r_count_73_io_out ? io_r_50_b : _GEN_14949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14951 = 8'h33 == r_count_73_io_out ? io_r_51_b : _GEN_14950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14952 = 8'h34 == r_count_73_io_out ? io_r_52_b : _GEN_14951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14953 = 8'h35 == r_count_73_io_out ? io_r_53_b : _GEN_14952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14954 = 8'h36 == r_count_73_io_out ? io_r_54_b : _GEN_14953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14955 = 8'h37 == r_count_73_io_out ? io_r_55_b : _GEN_14954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14956 = 8'h38 == r_count_73_io_out ? io_r_56_b : _GEN_14955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14957 = 8'h39 == r_count_73_io_out ? io_r_57_b : _GEN_14956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14958 = 8'h3a == r_count_73_io_out ? io_r_58_b : _GEN_14957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14959 = 8'h3b == r_count_73_io_out ? io_r_59_b : _GEN_14958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14960 = 8'h3c == r_count_73_io_out ? io_r_60_b : _GEN_14959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14961 = 8'h3d == r_count_73_io_out ? io_r_61_b : _GEN_14960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14962 = 8'h3e == r_count_73_io_out ? io_r_62_b : _GEN_14961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14963 = 8'h3f == r_count_73_io_out ? io_r_63_b : _GEN_14962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14964 = 8'h40 == r_count_73_io_out ? io_r_64_b : _GEN_14963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14965 = 8'h41 == r_count_73_io_out ? io_r_65_b : _GEN_14964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14966 = 8'h42 == r_count_73_io_out ? io_r_66_b : _GEN_14965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14967 = 8'h43 == r_count_73_io_out ? io_r_67_b : _GEN_14966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14968 = 8'h44 == r_count_73_io_out ? io_r_68_b : _GEN_14967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14969 = 8'h45 == r_count_73_io_out ? io_r_69_b : _GEN_14968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14970 = 8'h46 == r_count_73_io_out ? io_r_70_b : _GEN_14969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14971 = 8'h47 == r_count_73_io_out ? io_r_71_b : _GEN_14970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14972 = 8'h48 == r_count_73_io_out ? io_r_72_b : _GEN_14971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14973 = 8'h49 == r_count_73_io_out ? io_r_73_b : _GEN_14972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14974 = 8'h4a == r_count_73_io_out ? io_r_74_b : _GEN_14973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14975 = 8'h4b == r_count_73_io_out ? io_r_75_b : _GEN_14974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14976 = 8'h4c == r_count_73_io_out ? io_r_76_b : _GEN_14975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14977 = 8'h4d == r_count_73_io_out ? io_r_77_b : _GEN_14976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14978 = 8'h4e == r_count_73_io_out ? io_r_78_b : _GEN_14977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14979 = 8'h4f == r_count_73_io_out ? io_r_79_b : _GEN_14978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14980 = 8'h50 == r_count_73_io_out ? io_r_80_b : _GEN_14979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14981 = 8'h51 == r_count_73_io_out ? io_r_81_b : _GEN_14980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14982 = 8'h52 == r_count_73_io_out ? io_r_82_b : _GEN_14981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14983 = 8'h53 == r_count_73_io_out ? io_r_83_b : _GEN_14982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14984 = 8'h54 == r_count_73_io_out ? io_r_84_b : _GEN_14983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14985 = 8'h55 == r_count_73_io_out ? io_r_85_b : _GEN_14984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14986 = 8'h56 == r_count_73_io_out ? io_r_86_b : _GEN_14985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14987 = 8'h57 == r_count_73_io_out ? io_r_87_b : _GEN_14986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14988 = 8'h58 == r_count_73_io_out ? io_r_88_b : _GEN_14987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14989 = 8'h59 == r_count_73_io_out ? io_r_89_b : _GEN_14988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14990 = 8'h5a == r_count_73_io_out ? io_r_90_b : _GEN_14989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14991 = 8'h5b == r_count_73_io_out ? io_r_91_b : _GEN_14990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14992 = 8'h5c == r_count_73_io_out ? io_r_92_b : _GEN_14991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14993 = 8'h5d == r_count_73_io_out ? io_r_93_b : _GEN_14992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14994 = 8'h5e == r_count_73_io_out ? io_r_94_b : _GEN_14993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14995 = 8'h5f == r_count_73_io_out ? io_r_95_b : _GEN_14994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14996 = 8'h60 == r_count_73_io_out ? io_r_96_b : _GEN_14995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14997 = 8'h61 == r_count_73_io_out ? io_r_97_b : _GEN_14996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14998 = 8'h62 == r_count_73_io_out ? io_r_98_b : _GEN_14997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_14999 = 8'h63 == r_count_73_io_out ? io_r_99_b : _GEN_14998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15000 = 8'h64 == r_count_73_io_out ? io_r_100_b : _GEN_14999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15001 = 8'h65 == r_count_73_io_out ? io_r_101_b : _GEN_15000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15002 = 8'h66 == r_count_73_io_out ? io_r_102_b : _GEN_15001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15003 = 8'h67 == r_count_73_io_out ? io_r_103_b : _GEN_15002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15004 = 8'h68 == r_count_73_io_out ? io_r_104_b : _GEN_15003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15005 = 8'h69 == r_count_73_io_out ? io_r_105_b : _GEN_15004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15006 = 8'h6a == r_count_73_io_out ? io_r_106_b : _GEN_15005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15007 = 8'h6b == r_count_73_io_out ? io_r_107_b : _GEN_15006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15008 = 8'h6c == r_count_73_io_out ? io_r_108_b : _GEN_15007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15009 = 8'h6d == r_count_73_io_out ? io_r_109_b : _GEN_15008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15010 = 8'h6e == r_count_73_io_out ? io_r_110_b : _GEN_15009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15011 = 8'h6f == r_count_73_io_out ? io_r_111_b : _GEN_15010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15012 = 8'h70 == r_count_73_io_out ? io_r_112_b : _GEN_15011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15013 = 8'h71 == r_count_73_io_out ? io_r_113_b : _GEN_15012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15014 = 8'h72 == r_count_73_io_out ? io_r_114_b : _GEN_15013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15015 = 8'h73 == r_count_73_io_out ? io_r_115_b : _GEN_15014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15016 = 8'h74 == r_count_73_io_out ? io_r_116_b : _GEN_15015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15017 = 8'h75 == r_count_73_io_out ? io_r_117_b : _GEN_15016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15018 = 8'h76 == r_count_73_io_out ? io_r_118_b : _GEN_15017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15019 = 8'h77 == r_count_73_io_out ? io_r_119_b : _GEN_15018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15020 = 8'h78 == r_count_73_io_out ? io_r_120_b : _GEN_15019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15021 = 8'h79 == r_count_73_io_out ? io_r_121_b : _GEN_15020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15022 = 8'h7a == r_count_73_io_out ? io_r_122_b : _GEN_15021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15023 = 8'h7b == r_count_73_io_out ? io_r_123_b : _GEN_15022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15024 = 8'h7c == r_count_73_io_out ? io_r_124_b : _GEN_15023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15025 = 8'h7d == r_count_73_io_out ? io_r_125_b : _GEN_15024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15026 = 8'h7e == r_count_73_io_out ? io_r_126_b : _GEN_15025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15027 = 8'h7f == r_count_73_io_out ? io_r_127_b : _GEN_15026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15028 = 8'h80 == r_count_73_io_out ? io_r_128_b : _GEN_15027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15029 = 8'h81 == r_count_73_io_out ? io_r_129_b : _GEN_15028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15030 = 8'h82 == r_count_73_io_out ? io_r_130_b : _GEN_15029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15031 = 8'h83 == r_count_73_io_out ? io_r_131_b : _GEN_15030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15032 = 8'h84 == r_count_73_io_out ? io_r_132_b : _GEN_15031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15033 = 8'h85 == r_count_73_io_out ? io_r_133_b : _GEN_15032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15034 = 8'h86 == r_count_73_io_out ? io_r_134_b : _GEN_15033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15035 = 8'h87 == r_count_73_io_out ? io_r_135_b : _GEN_15034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15036 = 8'h88 == r_count_73_io_out ? io_r_136_b : _GEN_15035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15037 = 8'h89 == r_count_73_io_out ? io_r_137_b : _GEN_15036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15038 = 8'h8a == r_count_73_io_out ? io_r_138_b : _GEN_15037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15039 = 8'h8b == r_count_73_io_out ? io_r_139_b : _GEN_15038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15040 = 8'h8c == r_count_73_io_out ? io_r_140_b : _GEN_15039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15041 = 8'h8d == r_count_73_io_out ? io_r_141_b : _GEN_15040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15042 = 8'h8e == r_count_73_io_out ? io_r_142_b : _GEN_15041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15043 = 8'h8f == r_count_73_io_out ? io_r_143_b : _GEN_15042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15044 = 8'h90 == r_count_73_io_out ? io_r_144_b : _GEN_15043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15045 = 8'h91 == r_count_73_io_out ? io_r_145_b : _GEN_15044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15046 = 8'h92 == r_count_73_io_out ? io_r_146_b : _GEN_15045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15047 = 8'h93 == r_count_73_io_out ? io_r_147_b : _GEN_15046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15048 = 8'h94 == r_count_73_io_out ? io_r_148_b : _GEN_15047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15049 = 8'h95 == r_count_73_io_out ? io_r_149_b : _GEN_15048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15050 = 8'h96 == r_count_73_io_out ? io_r_150_b : _GEN_15049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15051 = 8'h97 == r_count_73_io_out ? io_r_151_b : _GEN_15050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15052 = 8'h98 == r_count_73_io_out ? io_r_152_b : _GEN_15051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15053 = 8'h99 == r_count_73_io_out ? io_r_153_b : _GEN_15052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15054 = 8'h9a == r_count_73_io_out ? io_r_154_b : _GEN_15053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15055 = 8'h9b == r_count_73_io_out ? io_r_155_b : _GEN_15054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15056 = 8'h9c == r_count_73_io_out ? io_r_156_b : _GEN_15055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15057 = 8'h9d == r_count_73_io_out ? io_r_157_b : _GEN_15056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15058 = 8'h9e == r_count_73_io_out ? io_r_158_b : _GEN_15057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15059 = 8'h9f == r_count_73_io_out ? io_r_159_b : _GEN_15058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15060 = 8'ha0 == r_count_73_io_out ? io_r_160_b : _GEN_15059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15061 = 8'ha1 == r_count_73_io_out ? io_r_161_b : _GEN_15060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15062 = 8'ha2 == r_count_73_io_out ? io_r_162_b : _GEN_15061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15063 = 8'ha3 == r_count_73_io_out ? io_r_163_b : _GEN_15062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15064 = 8'ha4 == r_count_73_io_out ? io_r_164_b : _GEN_15063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15065 = 8'ha5 == r_count_73_io_out ? io_r_165_b : _GEN_15064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15066 = 8'ha6 == r_count_73_io_out ? io_r_166_b : _GEN_15065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15067 = 8'ha7 == r_count_73_io_out ? io_r_167_b : _GEN_15066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15068 = 8'ha8 == r_count_73_io_out ? io_r_168_b : _GEN_15067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15069 = 8'ha9 == r_count_73_io_out ? io_r_169_b : _GEN_15068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15070 = 8'haa == r_count_73_io_out ? io_r_170_b : _GEN_15069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15071 = 8'hab == r_count_73_io_out ? io_r_171_b : _GEN_15070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15072 = 8'hac == r_count_73_io_out ? io_r_172_b : _GEN_15071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15073 = 8'had == r_count_73_io_out ? io_r_173_b : _GEN_15072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15074 = 8'hae == r_count_73_io_out ? io_r_174_b : _GEN_15073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15075 = 8'haf == r_count_73_io_out ? io_r_175_b : _GEN_15074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15076 = 8'hb0 == r_count_73_io_out ? io_r_176_b : _GEN_15075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15077 = 8'hb1 == r_count_73_io_out ? io_r_177_b : _GEN_15076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15078 = 8'hb2 == r_count_73_io_out ? io_r_178_b : _GEN_15077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15079 = 8'hb3 == r_count_73_io_out ? io_r_179_b : _GEN_15078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15080 = 8'hb4 == r_count_73_io_out ? io_r_180_b : _GEN_15079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15081 = 8'hb5 == r_count_73_io_out ? io_r_181_b : _GEN_15080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15082 = 8'hb6 == r_count_73_io_out ? io_r_182_b : _GEN_15081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15083 = 8'hb7 == r_count_73_io_out ? io_r_183_b : _GEN_15082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15084 = 8'hb8 == r_count_73_io_out ? io_r_184_b : _GEN_15083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15085 = 8'hb9 == r_count_73_io_out ? io_r_185_b : _GEN_15084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15086 = 8'hba == r_count_73_io_out ? io_r_186_b : _GEN_15085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15087 = 8'hbb == r_count_73_io_out ? io_r_187_b : _GEN_15086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15088 = 8'hbc == r_count_73_io_out ? io_r_188_b : _GEN_15087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15089 = 8'hbd == r_count_73_io_out ? io_r_189_b : _GEN_15088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15090 = 8'hbe == r_count_73_io_out ? io_r_190_b : _GEN_15089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15091 = 8'hbf == r_count_73_io_out ? io_r_191_b : _GEN_15090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15092 = 8'hc0 == r_count_73_io_out ? io_r_192_b : _GEN_15091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15093 = 8'hc1 == r_count_73_io_out ? io_r_193_b : _GEN_15092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15094 = 8'hc2 == r_count_73_io_out ? io_r_194_b : _GEN_15093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15095 = 8'hc3 == r_count_73_io_out ? io_r_195_b : _GEN_15094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15096 = 8'hc4 == r_count_73_io_out ? io_r_196_b : _GEN_15095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15097 = 8'hc5 == r_count_73_io_out ? io_r_197_b : _GEN_15096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15098 = 8'hc6 == r_count_73_io_out ? io_r_198_b : _GEN_15097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15101 = 8'h1 == r_count_74_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15102 = 8'h2 == r_count_74_io_out ? io_r_2_b : _GEN_15101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15103 = 8'h3 == r_count_74_io_out ? io_r_3_b : _GEN_15102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15104 = 8'h4 == r_count_74_io_out ? io_r_4_b : _GEN_15103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15105 = 8'h5 == r_count_74_io_out ? io_r_5_b : _GEN_15104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15106 = 8'h6 == r_count_74_io_out ? io_r_6_b : _GEN_15105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15107 = 8'h7 == r_count_74_io_out ? io_r_7_b : _GEN_15106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15108 = 8'h8 == r_count_74_io_out ? io_r_8_b : _GEN_15107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15109 = 8'h9 == r_count_74_io_out ? io_r_9_b : _GEN_15108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15110 = 8'ha == r_count_74_io_out ? io_r_10_b : _GEN_15109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15111 = 8'hb == r_count_74_io_out ? io_r_11_b : _GEN_15110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15112 = 8'hc == r_count_74_io_out ? io_r_12_b : _GEN_15111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15113 = 8'hd == r_count_74_io_out ? io_r_13_b : _GEN_15112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15114 = 8'he == r_count_74_io_out ? io_r_14_b : _GEN_15113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15115 = 8'hf == r_count_74_io_out ? io_r_15_b : _GEN_15114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15116 = 8'h10 == r_count_74_io_out ? io_r_16_b : _GEN_15115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15117 = 8'h11 == r_count_74_io_out ? io_r_17_b : _GEN_15116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15118 = 8'h12 == r_count_74_io_out ? io_r_18_b : _GEN_15117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15119 = 8'h13 == r_count_74_io_out ? io_r_19_b : _GEN_15118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15120 = 8'h14 == r_count_74_io_out ? io_r_20_b : _GEN_15119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15121 = 8'h15 == r_count_74_io_out ? io_r_21_b : _GEN_15120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15122 = 8'h16 == r_count_74_io_out ? io_r_22_b : _GEN_15121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15123 = 8'h17 == r_count_74_io_out ? io_r_23_b : _GEN_15122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15124 = 8'h18 == r_count_74_io_out ? io_r_24_b : _GEN_15123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15125 = 8'h19 == r_count_74_io_out ? io_r_25_b : _GEN_15124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15126 = 8'h1a == r_count_74_io_out ? io_r_26_b : _GEN_15125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15127 = 8'h1b == r_count_74_io_out ? io_r_27_b : _GEN_15126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15128 = 8'h1c == r_count_74_io_out ? io_r_28_b : _GEN_15127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15129 = 8'h1d == r_count_74_io_out ? io_r_29_b : _GEN_15128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15130 = 8'h1e == r_count_74_io_out ? io_r_30_b : _GEN_15129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15131 = 8'h1f == r_count_74_io_out ? io_r_31_b : _GEN_15130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15132 = 8'h20 == r_count_74_io_out ? io_r_32_b : _GEN_15131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15133 = 8'h21 == r_count_74_io_out ? io_r_33_b : _GEN_15132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15134 = 8'h22 == r_count_74_io_out ? io_r_34_b : _GEN_15133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15135 = 8'h23 == r_count_74_io_out ? io_r_35_b : _GEN_15134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15136 = 8'h24 == r_count_74_io_out ? io_r_36_b : _GEN_15135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15137 = 8'h25 == r_count_74_io_out ? io_r_37_b : _GEN_15136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15138 = 8'h26 == r_count_74_io_out ? io_r_38_b : _GEN_15137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15139 = 8'h27 == r_count_74_io_out ? io_r_39_b : _GEN_15138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15140 = 8'h28 == r_count_74_io_out ? io_r_40_b : _GEN_15139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15141 = 8'h29 == r_count_74_io_out ? io_r_41_b : _GEN_15140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15142 = 8'h2a == r_count_74_io_out ? io_r_42_b : _GEN_15141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15143 = 8'h2b == r_count_74_io_out ? io_r_43_b : _GEN_15142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15144 = 8'h2c == r_count_74_io_out ? io_r_44_b : _GEN_15143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15145 = 8'h2d == r_count_74_io_out ? io_r_45_b : _GEN_15144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15146 = 8'h2e == r_count_74_io_out ? io_r_46_b : _GEN_15145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15147 = 8'h2f == r_count_74_io_out ? io_r_47_b : _GEN_15146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15148 = 8'h30 == r_count_74_io_out ? io_r_48_b : _GEN_15147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15149 = 8'h31 == r_count_74_io_out ? io_r_49_b : _GEN_15148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15150 = 8'h32 == r_count_74_io_out ? io_r_50_b : _GEN_15149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15151 = 8'h33 == r_count_74_io_out ? io_r_51_b : _GEN_15150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15152 = 8'h34 == r_count_74_io_out ? io_r_52_b : _GEN_15151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15153 = 8'h35 == r_count_74_io_out ? io_r_53_b : _GEN_15152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15154 = 8'h36 == r_count_74_io_out ? io_r_54_b : _GEN_15153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15155 = 8'h37 == r_count_74_io_out ? io_r_55_b : _GEN_15154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15156 = 8'h38 == r_count_74_io_out ? io_r_56_b : _GEN_15155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15157 = 8'h39 == r_count_74_io_out ? io_r_57_b : _GEN_15156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15158 = 8'h3a == r_count_74_io_out ? io_r_58_b : _GEN_15157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15159 = 8'h3b == r_count_74_io_out ? io_r_59_b : _GEN_15158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15160 = 8'h3c == r_count_74_io_out ? io_r_60_b : _GEN_15159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15161 = 8'h3d == r_count_74_io_out ? io_r_61_b : _GEN_15160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15162 = 8'h3e == r_count_74_io_out ? io_r_62_b : _GEN_15161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15163 = 8'h3f == r_count_74_io_out ? io_r_63_b : _GEN_15162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15164 = 8'h40 == r_count_74_io_out ? io_r_64_b : _GEN_15163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15165 = 8'h41 == r_count_74_io_out ? io_r_65_b : _GEN_15164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15166 = 8'h42 == r_count_74_io_out ? io_r_66_b : _GEN_15165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15167 = 8'h43 == r_count_74_io_out ? io_r_67_b : _GEN_15166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15168 = 8'h44 == r_count_74_io_out ? io_r_68_b : _GEN_15167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15169 = 8'h45 == r_count_74_io_out ? io_r_69_b : _GEN_15168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15170 = 8'h46 == r_count_74_io_out ? io_r_70_b : _GEN_15169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15171 = 8'h47 == r_count_74_io_out ? io_r_71_b : _GEN_15170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15172 = 8'h48 == r_count_74_io_out ? io_r_72_b : _GEN_15171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15173 = 8'h49 == r_count_74_io_out ? io_r_73_b : _GEN_15172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15174 = 8'h4a == r_count_74_io_out ? io_r_74_b : _GEN_15173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15175 = 8'h4b == r_count_74_io_out ? io_r_75_b : _GEN_15174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15176 = 8'h4c == r_count_74_io_out ? io_r_76_b : _GEN_15175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15177 = 8'h4d == r_count_74_io_out ? io_r_77_b : _GEN_15176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15178 = 8'h4e == r_count_74_io_out ? io_r_78_b : _GEN_15177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15179 = 8'h4f == r_count_74_io_out ? io_r_79_b : _GEN_15178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15180 = 8'h50 == r_count_74_io_out ? io_r_80_b : _GEN_15179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15181 = 8'h51 == r_count_74_io_out ? io_r_81_b : _GEN_15180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15182 = 8'h52 == r_count_74_io_out ? io_r_82_b : _GEN_15181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15183 = 8'h53 == r_count_74_io_out ? io_r_83_b : _GEN_15182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15184 = 8'h54 == r_count_74_io_out ? io_r_84_b : _GEN_15183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15185 = 8'h55 == r_count_74_io_out ? io_r_85_b : _GEN_15184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15186 = 8'h56 == r_count_74_io_out ? io_r_86_b : _GEN_15185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15187 = 8'h57 == r_count_74_io_out ? io_r_87_b : _GEN_15186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15188 = 8'h58 == r_count_74_io_out ? io_r_88_b : _GEN_15187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15189 = 8'h59 == r_count_74_io_out ? io_r_89_b : _GEN_15188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15190 = 8'h5a == r_count_74_io_out ? io_r_90_b : _GEN_15189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15191 = 8'h5b == r_count_74_io_out ? io_r_91_b : _GEN_15190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15192 = 8'h5c == r_count_74_io_out ? io_r_92_b : _GEN_15191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15193 = 8'h5d == r_count_74_io_out ? io_r_93_b : _GEN_15192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15194 = 8'h5e == r_count_74_io_out ? io_r_94_b : _GEN_15193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15195 = 8'h5f == r_count_74_io_out ? io_r_95_b : _GEN_15194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15196 = 8'h60 == r_count_74_io_out ? io_r_96_b : _GEN_15195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15197 = 8'h61 == r_count_74_io_out ? io_r_97_b : _GEN_15196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15198 = 8'h62 == r_count_74_io_out ? io_r_98_b : _GEN_15197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15199 = 8'h63 == r_count_74_io_out ? io_r_99_b : _GEN_15198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15200 = 8'h64 == r_count_74_io_out ? io_r_100_b : _GEN_15199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15201 = 8'h65 == r_count_74_io_out ? io_r_101_b : _GEN_15200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15202 = 8'h66 == r_count_74_io_out ? io_r_102_b : _GEN_15201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15203 = 8'h67 == r_count_74_io_out ? io_r_103_b : _GEN_15202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15204 = 8'h68 == r_count_74_io_out ? io_r_104_b : _GEN_15203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15205 = 8'h69 == r_count_74_io_out ? io_r_105_b : _GEN_15204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15206 = 8'h6a == r_count_74_io_out ? io_r_106_b : _GEN_15205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15207 = 8'h6b == r_count_74_io_out ? io_r_107_b : _GEN_15206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15208 = 8'h6c == r_count_74_io_out ? io_r_108_b : _GEN_15207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15209 = 8'h6d == r_count_74_io_out ? io_r_109_b : _GEN_15208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15210 = 8'h6e == r_count_74_io_out ? io_r_110_b : _GEN_15209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15211 = 8'h6f == r_count_74_io_out ? io_r_111_b : _GEN_15210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15212 = 8'h70 == r_count_74_io_out ? io_r_112_b : _GEN_15211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15213 = 8'h71 == r_count_74_io_out ? io_r_113_b : _GEN_15212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15214 = 8'h72 == r_count_74_io_out ? io_r_114_b : _GEN_15213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15215 = 8'h73 == r_count_74_io_out ? io_r_115_b : _GEN_15214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15216 = 8'h74 == r_count_74_io_out ? io_r_116_b : _GEN_15215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15217 = 8'h75 == r_count_74_io_out ? io_r_117_b : _GEN_15216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15218 = 8'h76 == r_count_74_io_out ? io_r_118_b : _GEN_15217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15219 = 8'h77 == r_count_74_io_out ? io_r_119_b : _GEN_15218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15220 = 8'h78 == r_count_74_io_out ? io_r_120_b : _GEN_15219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15221 = 8'h79 == r_count_74_io_out ? io_r_121_b : _GEN_15220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15222 = 8'h7a == r_count_74_io_out ? io_r_122_b : _GEN_15221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15223 = 8'h7b == r_count_74_io_out ? io_r_123_b : _GEN_15222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15224 = 8'h7c == r_count_74_io_out ? io_r_124_b : _GEN_15223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15225 = 8'h7d == r_count_74_io_out ? io_r_125_b : _GEN_15224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15226 = 8'h7e == r_count_74_io_out ? io_r_126_b : _GEN_15225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15227 = 8'h7f == r_count_74_io_out ? io_r_127_b : _GEN_15226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15228 = 8'h80 == r_count_74_io_out ? io_r_128_b : _GEN_15227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15229 = 8'h81 == r_count_74_io_out ? io_r_129_b : _GEN_15228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15230 = 8'h82 == r_count_74_io_out ? io_r_130_b : _GEN_15229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15231 = 8'h83 == r_count_74_io_out ? io_r_131_b : _GEN_15230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15232 = 8'h84 == r_count_74_io_out ? io_r_132_b : _GEN_15231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15233 = 8'h85 == r_count_74_io_out ? io_r_133_b : _GEN_15232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15234 = 8'h86 == r_count_74_io_out ? io_r_134_b : _GEN_15233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15235 = 8'h87 == r_count_74_io_out ? io_r_135_b : _GEN_15234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15236 = 8'h88 == r_count_74_io_out ? io_r_136_b : _GEN_15235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15237 = 8'h89 == r_count_74_io_out ? io_r_137_b : _GEN_15236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15238 = 8'h8a == r_count_74_io_out ? io_r_138_b : _GEN_15237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15239 = 8'h8b == r_count_74_io_out ? io_r_139_b : _GEN_15238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15240 = 8'h8c == r_count_74_io_out ? io_r_140_b : _GEN_15239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15241 = 8'h8d == r_count_74_io_out ? io_r_141_b : _GEN_15240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15242 = 8'h8e == r_count_74_io_out ? io_r_142_b : _GEN_15241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15243 = 8'h8f == r_count_74_io_out ? io_r_143_b : _GEN_15242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15244 = 8'h90 == r_count_74_io_out ? io_r_144_b : _GEN_15243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15245 = 8'h91 == r_count_74_io_out ? io_r_145_b : _GEN_15244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15246 = 8'h92 == r_count_74_io_out ? io_r_146_b : _GEN_15245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15247 = 8'h93 == r_count_74_io_out ? io_r_147_b : _GEN_15246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15248 = 8'h94 == r_count_74_io_out ? io_r_148_b : _GEN_15247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15249 = 8'h95 == r_count_74_io_out ? io_r_149_b : _GEN_15248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15250 = 8'h96 == r_count_74_io_out ? io_r_150_b : _GEN_15249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15251 = 8'h97 == r_count_74_io_out ? io_r_151_b : _GEN_15250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15252 = 8'h98 == r_count_74_io_out ? io_r_152_b : _GEN_15251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15253 = 8'h99 == r_count_74_io_out ? io_r_153_b : _GEN_15252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15254 = 8'h9a == r_count_74_io_out ? io_r_154_b : _GEN_15253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15255 = 8'h9b == r_count_74_io_out ? io_r_155_b : _GEN_15254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15256 = 8'h9c == r_count_74_io_out ? io_r_156_b : _GEN_15255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15257 = 8'h9d == r_count_74_io_out ? io_r_157_b : _GEN_15256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15258 = 8'h9e == r_count_74_io_out ? io_r_158_b : _GEN_15257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15259 = 8'h9f == r_count_74_io_out ? io_r_159_b : _GEN_15258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15260 = 8'ha0 == r_count_74_io_out ? io_r_160_b : _GEN_15259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15261 = 8'ha1 == r_count_74_io_out ? io_r_161_b : _GEN_15260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15262 = 8'ha2 == r_count_74_io_out ? io_r_162_b : _GEN_15261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15263 = 8'ha3 == r_count_74_io_out ? io_r_163_b : _GEN_15262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15264 = 8'ha4 == r_count_74_io_out ? io_r_164_b : _GEN_15263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15265 = 8'ha5 == r_count_74_io_out ? io_r_165_b : _GEN_15264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15266 = 8'ha6 == r_count_74_io_out ? io_r_166_b : _GEN_15265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15267 = 8'ha7 == r_count_74_io_out ? io_r_167_b : _GEN_15266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15268 = 8'ha8 == r_count_74_io_out ? io_r_168_b : _GEN_15267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15269 = 8'ha9 == r_count_74_io_out ? io_r_169_b : _GEN_15268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15270 = 8'haa == r_count_74_io_out ? io_r_170_b : _GEN_15269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15271 = 8'hab == r_count_74_io_out ? io_r_171_b : _GEN_15270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15272 = 8'hac == r_count_74_io_out ? io_r_172_b : _GEN_15271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15273 = 8'had == r_count_74_io_out ? io_r_173_b : _GEN_15272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15274 = 8'hae == r_count_74_io_out ? io_r_174_b : _GEN_15273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15275 = 8'haf == r_count_74_io_out ? io_r_175_b : _GEN_15274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15276 = 8'hb0 == r_count_74_io_out ? io_r_176_b : _GEN_15275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15277 = 8'hb1 == r_count_74_io_out ? io_r_177_b : _GEN_15276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15278 = 8'hb2 == r_count_74_io_out ? io_r_178_b : _GEN_15277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15279 = 8'hb3 == r_count_74_io_out ? io_r_179_b : _GEN_15278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15280 = 8'hb4 == r_count_74_io_out ? io_r_180_b : _GEN_15279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15281 = 8'hb5 == r_count_74_io_out ? io_r_181_b : _GEN_15280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15282 = 8'hb6 == r_count_74_io_out ? io_r_182_b : _GEN_15281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15283 = 8'hb7 == r_count_74_io_out ? io_r_183_b : _GEN_15282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15284 = 8'hb8 == r_count_74_io_out ? io_r_184_b : _GEN_15283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15285 = 8'hb9 == r_count_74_io_out ? io_r_185_b : _GEN_15284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15286 = 8'hba == r_count_74_io_out ? io_r_186_b : _GEN_15285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15287 = 8'hbb == r_count_74_io_out ? io_r_187_b : _GEN_15286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15288 = 8'hbc == r_count_74_io_out ? io_r_188_b : _GEN_15287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15289 = 8'hbd == r_count_74_io_out ? io_r_189_b : _GEN_15288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15290 = 8'hbe == r_count_74_io_out ? io_r_190_b : _GEN_15289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15291 = 8'hbf == r_count_74_io_out ? io_r_191_b : _GEN_15290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15292 = 8'hc0 == r_count_74_io_out ? io_r_192_b : _GEN_15291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15293 = 8'hc1 == r_count_74_io_out ? io_r_193_b : _GEN_15292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15294 = 8'hc2 == r_count_74_io_out ? io_r_194_b : _GEN_15293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15295 = 8'hc3 == r_count_74_io_out ? io_r_195_b : _GEN_15294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15296 = 8'hc4 == r_count_74_io_out ? io_r_196_b : _GEN_15295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15297 = 8'hc5 == r_count_74_io_out ? io_r_197_b : _GEN_15296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15298 = 8'hc6 == r_count_74_io_out ? io_r_198_b : _GEN_15297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15301 = 8'h1 == r_count_75_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15302 = 8'h2 == r_count_75_io_out ? io_r_2_b : _GEN_15301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15303 = 8'h3 == r_count_75_io_out ? io_r_3_b : _GEN_15302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15304 = 8'h4 == r_count_75_io_out ? io_r_4_b : _GEN_15303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15305 = 8'h5 == r_count_75_io_out ? io_r_5_b : _GEN_15304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15306 = 8'h6 == r_count_75_io_out ? io_r_6_b : _GEN_15305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15307 = 8'h7 == r_count_75_io_out ? io_r_7_b : _GEN_15306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15308 = 8'h8 == r_count_75_io_out ? io_r_8_b : _GEN_15307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15309 = 8'h9 == r_count_75_io_out ? io_r_9_b : _GEN_15308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15310 = 8'ha == r_count_75_io_out ? io_r_10_b : _GEN_15309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15311 = 8'hb == r_count_75_io_out ? io_r_11_b : _GEN_15310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15312 = 8'hc == r_count_75_io_out ? io_r_12_b : _GEN_15311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15313 = 8'hd == r_count_75_io_out ? io_r_13_b : _GEN_15312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15314 = 8'he == r_count_75_io_out ? io_r_14_b : _GEN_15313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15315 = 8'hf == r_count_75_io_out ? io_r_15_b : _GEN_15314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15316 = 8'h10 == r_count_75_io_out ? io_r_16_b : _GEN_15315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15317 = 8'h11 == r_count_75_io_out ? io_r_17_b : _GEN_15316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15318 = 8'h12 == r_count_75_io_out ? io_r_18_b : _GEN_15317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15319 = 8'h13 == r_count_75_io_out ? io_r_19_b : _GEN_15318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15320 = 8'h14 == r_count_75_io_out ? io_r_20_b : _GEN_15319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15321 = 8'h15 == r_count_75_io_out ? io_r_21_b : _GEN_15320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15322 = 8'h16 == r_count_75_io_out ? io_r_22_b : _GEN_15321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15323 = 8'h17 == r_count_75_io_out ? io_r_23_b : _GEN_15322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15324 = 8'h18 == r_count_75_io_out ? io_r_24_b : _GEN_15323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15325 = 8'h19 == r_count_75_io_out ? io_r_25_b : _GEN_15324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15326 = 8'h1a == r_count_75_io_out ? io_r_26_b : _GEN_15325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15327 = 8'h1b == r_count_75_io_out ? io_r_27_b : _GEN_15326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15328 = 8'h1c == r_count_75_io_out ? io_r_28_b : _GEN_15327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15329 = 8'h1d == r_count_75_io_out ? io_r_29_b : _GEN_15328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15330 = 8'h1e == r_count_75_io_out ? io_r_30_b : _GEN_15329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15331 = 8'h1f == r_count_75_io_out ? io_r_31_b : _GEN_15330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15332 = 8'h20 == r_count_75_io_out ? io_r_32_b : _GEN_15331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15333 = 8'h21 == r_count_75_io_out ? io_r_33_b : _GEN_15332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15334 = 8'h22 == r_count_75_io_out ? io_r_34_b : _GEN_15333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15335 = 8'h23 == r_count_75_io_out ? io_r_35_b : _GEN_15334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15336 = 8'h24 == r_count_75_io_out ? io_r_36_b : _GEN_15335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15337 = 8'h25 == r_count_75_io_out ? io_r_37_b : _GEN_15336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15338 = 8'h26 == r_count_75_io_out ? io_r_38_b : _GEN_15337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15339 = 8'h27 == r_count_75_io_out ? io_r_39_b : _GEN_15338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15340 = 8'h28 == r_count_75_io_out ? io_r_40_b : _GEN_15339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15341 = 8'h29 == r_count_75_io_out ? io_r_41_b : _GEN_15340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15342 = 8'h2a == r_count_75_io_out ? io_r_42_b : _GEN_15341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15343 = 8'h2b == r_count_75_io_out ? io_r_43_b : _GEN_15342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15344 = 8'h2c == r_count_75_io_out ? io_r_44_b : _GEN_15343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15345 = 8'h2d == r_count_75_io_out ? io_r_45_b : _GEN_15344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15346 = 8'h2e == r_count_75_io_out ? io_r_46_b : _GEN_15345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15347 = 8'h2f == r_count_75_io_out ? io_r_47_b : _GEN_15346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15348 = 8'h30 == r_count_75_io_out ? io_r_48_b : _GEN_15347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15349 = 8'h31 == r_count_75_io_out ? io_r_49_b : _GEN_15348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15350 = 8'h32 == r_count_75_io_out ? io_r_50_b : _GEN_15349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15351 = 8'h33 == r_count_75_io_out ? io_r_51_b : _GEN_15350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15352 = 8'h34 == r_count_75_io_out ? io_r_52_b : _GEN_15351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15353 = 8'h35 == r_count_75_io_out ? io_r_53_b : _GEN_15352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15354 = 8'h36 == r_count_75_io_out ? io_r_54_b : _GEN_15353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15355 = 8'h37 == r_count_75_io_out ? io_r_55_b : _GEN_15354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15356 = 8'h38 == r_count_75_io_out ? io_r_56_b : _GEN_15355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15357 = 8'h39 == r_count_75_io_out ? io_r_57_b : _GEN_15356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15358 = 8'h3a == r_count_75_io_out ? io_r_58_b : _GEN_15357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15359 = 8'h3b == r_count_75_io_out ? io_r_59_b : _GEN_15358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15360 = 8'h3c == r_count_75_io_out ? io_r_60_b : _GEN_15359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15361 = 8'h3d == r_count_75_io_out ? io_r_61_b : _GEN_15360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15362 = 8'h3e == r_count_75_io_out ? io_r_62_b : _GEN_15361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15363 = 8'h3f == r_count_75_io_out ? io_r_63_b : _GEN_15362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15364 = 8'h40 == r_count_75_io_out ? io_r_64_b : _GEN_15363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15365 = 8'h41 == r_count_75_io_out ? io_r_65_b : _GEN_15364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15366 = 8'h42 == r_count_75_io_out ? io_r_66_b : _GEN_15365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15367 = 8'h43 == r_count_75_io_out ? io_r_67_b : _GEN_15366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15368 = 8'h44 == r_count_75_io_out ? io_r_68_b : _GEN_15367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15369 = 8'h45 == r_count_75_io_out ? io_r_69_b : _GEN_15368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15370 = 8'h46 == r_count_75_io_out ? io_r_70_b : _GEN_15369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15371 = 8'h47 == r_count_75_io_out ? io_r_71_b : _GEN_15370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15372 = 8'h48 == r_count_75_io_out ? io_r_72_b : _GEN_15371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15373 = 8'h49 == r_count_75_io_out ? io_r_73_b : _GEN_15372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15374 = 8'h4a == r_count_75_io_out ? io_r_74_b : _GEN_15373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15375 = 8'h4b == r_count_75_io_out ? io_r_75_b : _GEN_15374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15376 = 8'h4c == r_count_75_io_out ? io_r_76_b : _GEN_15375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15377 = 8'h4d == r_count_75_io_out ? io_r_77_b : _GEN_15376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15378 = 8'h4e == r_count_75_io_out ? io_r_78_b : _GEN_15377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15379 = 8'h4f == r_count_75_io_out ? io_r_79_b : _GEN_15378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15380 = 8'h50 == r_count_75_io_out ? io_r_80_b : _GEN_15379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15381 = 8'h51 == r_count_75_io_out ? io_r_81_b : _GEN_15380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15382 = 8'h52 == r_count_75_io_out ? io_r_82_b : _GEN_15381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15383 = 8'h53 == r_count_75_io_out ? io_r_83_b : _GEN_15382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15384 = 8'h54 == r_count_75_io_out ? io_r_84_b : _GEN_15383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15385 = 8'h55 == r_count_75_io_out ? io_r_85_b : _GEN_15384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15386 = 8'h56 == r_count_75_io_out ? io_r_86_b : _GEN_15385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15387 = 8'h57 == r_count_75_io_out ? io_r_87_b : _GEN_15386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15388 = 8'h58 == r_count_75_io_out ? io_r_88_b : _GEN_15387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15389 = 8'h59 == r_count_75_io_out ? io_r_89_b : _GEN_15388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15390 = 8'h5a == r_count_75_io_out ? io_r_90_b : _GEN_15389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15391 = 8'h5b == r_count_75_io_out ? io_r_91_b : _GEN_15390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15392 = 8'h5c == r_count_75_io_out ? io_r_92_b : _GEN_15391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15393 = 8'h5d == r_count_75_io_out ? io_r_93_b : _GEN_15392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15394 = 8'h5e == r_count_75_io_out ? io_r_94_b : _GEN_15393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15395 = 8'h5f == r_count_75_io_out ? io_r_95_b : _GEN_15394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15396 = 8'h60 == r_count_75_io_out ? io_r_96_b : _GEN_15395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15397 = 8'h61 == r_count_75_io_out ? io_r_97_b : _GEN_15396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15398 = 8'h62 == r_count_75_io_out ? io_r_98_b : _GEN_15397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15399 = 8'h63 == r_count_75_io_out ? io_r_99_b : _GEN_15398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15400 = 8'h64 == r_count_75_io_out ? io_r_100_b : _GEN_15399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15401 = 8'h65 == r_count_75_io_out ? io_r_101_b : _GEN_15400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15402 = 8'h66 == r_count_75_io_out ? io_r_102_b : _GEN_15401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15403 = 8'h67 == r_count_75_io_out ? io_r_103_b : _GEN_15402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15404 = 8'h68 == r_count_75_io_out ? io_r_104_b : _GEN_15403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15405 = 8'h69 == r_count_75_io_out ? io_r_105_b : _GEN_15404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15406 = 8'h6a == r_count_75_io_out ? io_r_106_b : _GEN_15405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15407 = 8'h6b == r_count_75_io_out ? io_r_107_b : _GEN_15406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15408 = 8'h6c == r_count_75_io_out ? io_r_108_b : _GEN_15407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15409 = 8'h6d == r_count_75_io_out ? io_r_109_b : _GEN_15408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15410 = 8'h6e == r_count_75_io_out ? io_r_110_b : _GEN_15409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15411 = 8'h6f == r_count_75_io_out ? io_r_111_b : _GEN_15410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15412 = 8'h70 == r_count_75_io_out ? io_r_112_b : _GEN_15411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15413 = 8'h71 == r_count_75_io_out ? io_r_113_b : _GEN_15412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15414 = 8'h72 == r_count_75_io_out ? io_r_114_b : _GEN_15413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15415 = 8'h73 == r_count_75_io_out ? io_r_115_b : _GEN_15414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15416 = 8'h74 == r_count_75_io_out ? io_r_116_b : _GEN_15415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15417 = 8'h75 == r_count_75_io_out ? io_r_117_b : _GEN_15416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15418 = 8'h76 == r_count_75_io_out ? io_r_118_b : _GEN_15417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15419 = 8'h77 == r_count_75_io_out ? io_r_119_b : _GEN_15418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15420 = 8'h78 == r_count_75_io_out ? io_r_120_b : _GEN_15419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15421 = 8'h79 == r_count_75_io_out ? io_r_121_b : _GEN_15420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15422 = 8'h7a == r_count_75_io_out ? io_r_122_b : _GEN_15421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15423 = 8'h7b == r_count_75_io_out ? io_r_123_b : _GEN_15422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15424 = 8'h7c == r_count_75_io_out ? io_r_124_b : _GEN_15423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15425 = 8'h7d == r_count_75_io_out ? io_r_125_b : _GEN_15424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15426 = 8'h7e == r_count_75_io_out ? io_r_126_b : _GEN_15425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15427 = 8'h7f == r_count_75_io_out ? io_r_127_b : _GEN_15426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15428 = 8'h80 == r_count_75_io_out ? io_r_128_b : _GEN_15427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15429 = 8'h81 == r_count_75_io_out ? io_r_129_b : _GEN_15428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15430 = 8'h82 == r_count_75_io_out ? io_r_130_b : _GEN_15429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15431 = 8'h83 == r_count_75_io_out ? io_r_131_b : _GEN_15430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15432 = 8'h84 == r_count_75_io_out ? io_r_132_b : _GEN_15431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15433 = 8'h85 == r_count_75_io_out ? io_r_133_b : _GEN_15432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15434 = 8'h86 == r_count_75_io_out ? io_r_134_b : _GEN_15433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15435 = 8'h87 == r_count_75_io_out ? io_r_135_b : _GEN_15434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15436 = 8'h88 == r_count_75_io_out ? io_r_136_b : _GEN_15435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15437 = 8'h89 == r_count_75_io_out ? io_r_137_b : _GEN_15436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15438 = 8'h8a == r_count_75_io_out ? io_r_138_b : _GEN_15437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15439 = 8'h8b == r_count_75_io_out ? io_r_139_b : _GEN_15438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15440 = 8'h8c == r_count_75_io_out ? io_r_140_b : _GEN_15439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15441 = 8'h8d == r_count_75_io_out ? io_r_141_b : _GEN_15440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15442 = 8'h8e == r_count_75_io_out ? io_r_142_b : _GEN_15441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15443 = 8'h8f == r_count_75_io_out ? io_r_143_b : _GEN_15442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15444 = 8'h90 == r_count_75_io_out ? io_r_144_b : _GEN_15443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15445 = 8'h91 == r_count_75_io_out ? io_r_145_b : _GEN_15444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15446 = 8'h92 == r_count_75_io_out ? io_r_146_b : _GEN_15445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15447 = 8'h93 == r_count_75_io_out ? io_r_147_b : _GEN_15446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15448 = 8'h94 == r_count_75_io_out ? io_r_148_b : _GEN_15447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15449 = 8'h95 == r_count_75_io_out ? io_r_149_b : _GEN_15448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15450 = 8'h96 == r_count_75_io_out ? io_r_150_b : _GEN_15449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15451 = 8'h97 == r_count_75_io_out ? io_r_151_b : _GEN_15450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15452 = 8'h98 == r_count_75_io_out ? io_r_152_b : _GEN_15451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15453 = 8'h99 == r_count_75_io_out ? io_r_153_b : _GEN_15452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15454 = 8'h9a == r_count_75_io_out ? io_r_154_b : _GEN_15453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15455 = 8'h9b == r_count_75_io_out ? io_r_155_b : _GEN_15454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15456 = 8'h9c == r_count_75_io_out ? io_r_156_b : _GEN_15455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15457 = 8'h9d == r_count_75_io_out ? io_r_157_b : _GEN_15456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15458 = 8'h9e == r_count_75_io_out ? io_r_158_b : _GEN_15457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15459 = 8'h9f == r_count_75_io_out ? io_r_159_b : _GEN_15458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15460 = 8'ha0 == r_count_75_io_out ? io_r_160_b : _GEN_15459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15461 = 8'ha1 == r_count_75_io_out ? io_r_161_b : _GEN_15460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15462 = 8'ha2 == r_count_75_io_out ? io_r_162_b : _GEN_15461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15463 = 8'ha3 == r_count_75_io_out ? io_r_163_b : _GEN_15462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15464 = 8'ha4 == r_count_75_io_out ? io_r_164_b : _GEN_15463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15465 = 8'ha5 == r_count_75_io_out ? io_r_165_b : _GEN_15464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15466 = 8'ha6 == r_count_75_io_out ? io_r_166_b : _GEN_15465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15467 = 8'ha7 == r_count_75_io_out ? io_r_167_b : _GEN_15466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15468 = 8'ha8 == r_count_75_io_out ? io_r_168_b : _GEN_15467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15469 = 8'ha9 == r_count_75_io_out ? io_r_169_b : _GEN_15468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15470 = 8'haa == r_count_75_io_out ? io_r_170_b : _GEN_15469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15471 = 8'hab == r_count_75_io_out ? io_r_171_b : _GEN_15470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15472 = 8'hac == r_count_75_io_out ? io_r_172_b : _GEN_15471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15473 = 8'had == r_count_75_io_out ? io_r_173_b : _GEN_15472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15474 = 8'hae == r_count_75_io_out ? io_r_174_b : _GEN_15473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15475 = 8'haf == r_count_75_io_out ? io_r_175_b : _GEN_15474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15476 = 8'hb0 == r_count_75_io_out ? io_r_176_b : _GEN_15475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15477 = 8'hb1 == r_count_75_io_out ? io_r_177_b : _GEN_15476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15478 = 8'hb2 == r_count_75_io_out ? io_r_178_b : _GEN_15477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15479 = 8'hb3 == r_count_75_io_out ? io_r_179_b : _GEN_15478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15480 = 8'hb4 == r_count_75_io_out ? io_r_180_b : _GEN_15479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15481 = 8'hb5 == r_count_75_io_out ? io_r_181_b : _GEN_15480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15482 = 8'hb6 == r_count_75_io_out ? io_r_182_b : _GEN_15481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15483 = 8'hb7 == r_count_75_io_out ? io_r_183_b : _GEN_15482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15484 = 8'hb8 == r_count_75_io_out ? io_r_184_b : _GEN_15483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15485 = 8'hb9 == r_count_75_io_out ? io_r_185_b : _GEN_15484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15486 = 8'hba == r_count_75_io_out ? io_r_186_b : _GEN_15485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15487 = 8'hbb == r_count_75_io_out ? io_r_187_b : _GEN_15486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15488 = 8'hbc == r_count_75_io_out ? io_r_188_b : _GEN_15487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15489 = 8'hbd == r_count_75_io_out ? io_r_189_b : _GEN_15488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15490 = 8'hbe == r_count_75_io_out ? io_r_190_b : _GEN_15489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15491 = 8'hbf == r_count_75_io_out ? io_r_191_b : _GEN_15490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15492 = 8'hc0 == r_count_75_io_out ? io_r_192_b : _GEN_15491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15493 = 8'hc1 == r_count_75_io_out ? io_r_193_b : _GEN_15492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15494 = 8'hc2 == r_count_75_io_out ? io_r_194_b : _GEN_15493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15495 = 8'hc3 == r_count_75_io_out ? io_r_195_b : _GEN_15494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15496 = 8'hc4 == r_count_75_io_out ? io_r_196_b : _GEN_15495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15497 = 8'hc5 == r_count_75_io_out ? io_r_197_b : _GEN_15496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15498 = 8'hc6 == r_count_75_io_out ? io_r_198_b : _GEN_15497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15501 = 8'h1 == r_count_76_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15502 = 8'h2 == r_count_76_io_out ? io_r_2_b : _GEN_15501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15503 = 8'h3 == r_count_76_io_out ? io_r_3_b : _GEN_15502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15504 = 8'h4 == r_count_76_io_out ? io_r_4_b : _GEN_15503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15505 = 8'h5 == r_count_76_io_out ? io_r_5_b : _GEN_15504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15506 = 8'h6 == r_count_76_io_out ? io_r_6_b : _GEN_15505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15507 = 8'h7 == r_count_76_io_out ? io_r_7_b : _GEN_15506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15508 = 8'h8 == r_count_76_io_out ? io_r_8_b : _GEN_15507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15509 = 8'h9 == r_count_76_io_out ? io_r_9_b : _GEN_15508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15510 = 8'ha == r_count_76_io_out ? io_r_10_b : _GEN_15509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15511 = 8'hb == r_count_76_io_out ? io_r_11_b : _GEN_15510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15512 = 8'hc == r_count_76_io_out ? io_r_12_b : _GEN_15511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15513 = 8'hd == r_count_76_io_out ? io_r_13_b : _GEN_15512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15514 = 8'he == r_count_76_io_out ? io_r_14_b : _GEN_15513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15515 = 8'hf == r_count_76_io_out ? io_r_15_b : _GEN_15514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15516 = 8'h10 == r_count_76_io_out ? io_r_16_b : _GEN_15515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15517 = 8'h11 == r_count_76_io_out ? io_r_17_b : _GEN_15516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15518 = 8'h12 == r_count_76_io_out ? io_r_18_b : _GEN_15517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15519 = 8'h13 == r_count_76_io_out ? io_r_19_b : _GEN_15518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15520 = 8'h14 == r_count_76_io_out ? io_r_20_b : _GEN_15519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15521 = 8'h15 == r_count_76_io_out ? io_r_21_b : _GEN_15520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15522 = 8'h16 == r_count_76_io_out ? io_r_22_b : _GEN_15521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15523 = 8'h17 == r_count_76_io_out ? io_r_23_b : _GEN_15522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15524 = 8'h18 == r_count_76_io_out ? io_r_24_b : _GEN_15523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15525 = 8'h19 == r_count_76_io_out ? io_r_25_b : _GEN_15524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15526 = 8'h1a == r_count_76_io_out ? io_r_26_b : _GEN_15525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15527 = 8'h1b == r_count_76_io_out ? io_r_27_b : _GEN_15526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15528 = 8'h1c == r_count_76_io_out ? io_r_28_b : _GEN_15527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15529 = 8'h1d == r_count_76_io_out ? io_r_29_b : _GEN_15528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15530 = 8'h1e == r_count_76_io_out ? io_r_30_b : _GEN_15529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15531 = 8'h1f == r_count_76_io_out ? io_r_31_b : _GEN_15530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15532 = 8'h20 == r_count_76_io_out ? io_r_32_b : _GEN_15531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15533 = 8'h21 == r_count_76_io_out ? io_r_33_b : _GEN_15532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15534 = 8'h22 == r_count_76_io_out ? io_r_34_b : _GEN_15533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15535 = 8'h23 == r_count_76_io_out ? io_r_35_b : _GEN_15534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15536 = 8'h24 == r_count_76_io_out ? io_r_36_b : _GEN_15535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15537 = 8'h25 == r_count_76_io_out ? io_r_37_b : _GEN_15536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15538 = 8'h26 == r_count_76_io_out ? io_r_38_b : _GEN_15537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15539 = 8'h27 == r_count_76_io_out ? io_r_39_b : _GEN_15538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15540 = 8'h28 == r_count_76_io_out ? io_r_40_b : _GEN_15539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15541 = 8'h29 == r_count_76_io_out ? io_r_41_b : _GEN_15540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15542 = 8'h2a == r_count_76_io_out ? io_r_42_b : _GEN_15541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15543 = 8'h2b == r_count_76_io_out ? io_r_43_b : _GEN_15542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15544 = 8'h2c == r_count_76_io_out ? io_r_44_b : _GEN_15543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15545 = 8'h2d == r_count_76_io_out ? io_r_45_b : _GEN_15544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15546 = 8'h2e == r_count_76_io_out ? io_r_46_b : _GEN_15545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15547 = 8'h2f == r_count_76_io_out ? io_r_47_b : _GEN_15546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15548 = 8'h30 == r_count_76_io_out ? io_r_48_b : _GEN_15547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15549 = 8'h31 == r_count_76_io_out ? io_r_49_b : _GEN_15548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15550 = 8'h32 == r_count_76_io_out ? io_r_50_b : _GEN_15549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15551 = 8'h33 == r_count_76_io_out ? io_r_51_b : _GEN_15550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15552 = 8'h34 == r_count_76_io_out ? io_r_52_b : _GEN_15551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15553 = 8'h35 == r_count_76_io_out ? io_r_53_b : _GEN_15552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15554 = 8'h36 == r_count_76_io_out ? io_r_54_b : _GEN_15553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15555 = 8'h37 == r_count_76_io_out ? io_r_55_b : _GEN_15554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15556 = 8'h38 == r_count_76_io_out ? io_r_56_b : _GEN_15555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15557 = 8'h39 == r_count_76_io_out ? io_r_57_b : _GEN_15556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15558 = 8'h3a == r_count_76_io_out ? io_r_58_b : _GEN_15557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15559 = 8'h3b == r_count_76_io_out ? io_r_59_b : _GEN_15558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15560 = 8'h3c == r_count_76_io_out ? io_r_60_b : _GEN_15559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15561 = 8'h3d == r_count_76_io_out ? io_r_61_b : _GEN_15560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15562 = 8'h3e == r_count_76_io_out ? io_r_62_b : _GEN_15561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15563 = 8'h3f == r_count_76_io_out ? io_r_63_b : _GEN_15562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15564 = 8'h40 == r_count_76_io_out ? io_r_64_b : _GEN_15563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15565 = 8'h41 == r_count_76_io_out ? io_r_65_b : _GEN_15564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15566 = 8'h42 == r_count_76_io_out ? io_r_66_b : _GEN_15565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15567 = 8'h43 == r_count_76_io_out ? io_r_67_b : _GEN_15566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15568 = 8'h44 == r_count_76_io_out ? io_r_68_b : _GEN_15567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15569 = 8'h45 == r_count_76_io_out ? io_r_69_b : _GEN_15568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15570 = 8'h46 == r_count_76_io_out ? io_r_70_b : _GEN_15569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15571 = 8'h47 == r_count_76_io_out ? io_r_71_b : _GEN_15570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15572 = 8'h48 == r_count_76_io_out ? io_r_72_b : _GEN_15571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15573 = 8'h49 == r_count_76_io_out ? io_r_73_b : _GEN_15572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15574 = 8'h4a == r_count_76_io_out ? io_r_74_b : _GEN_15573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15575 = 8'h4b == r_count_76_io_out ? io_r_75_b : _GEN_15574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15576 = 8'h4c == r_count_76_io_out ? io_r_76_b : _GEN_15575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15577 = 8'h4d == r_count_76_io_out ? io_r_77_b : _GEN_15576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15578 = 8'h4e == r_count_76_io_out ? io_r_78_b : _GEN_15577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15579 = 8'h4f == r_count_76_io_out ? io_r_79_b : _GEN_15578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15580 = 8'h50 == r_count_76_io_out ? io_r_80_b : _GEN_15579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15581 = 8'h51 == r_count_76_io_out ? io_r_81_b : _GEN_15580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15582 = 8'h52 == r_count_76_io_out ? io_r_82_b : _GEN_15581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15583 = 8'h53 == r_count_76_io_out ? io_r_83_b : _GEN_15582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15584 = 8'h54 == r_count_76_io_out ? io_r_84_b : _GEN_15583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15585 = 8'h55 == r_count_76_io_out ? io_r_85_b : _GEN_15584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15586 = 8'h56 == r_count_76_io_out ? io_r_86_b : _GEN_15585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15587 = 8'h57 == r_count_76_io_out ? io_r_87_b : _GEN_15586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15588 = 8'h58 == r_count_76_io_out ? io_r_88_b : _GEN_15587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15589 = 8'h59 == r_count_76_io_out ? io_r_89_b : _GEN_15588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15590 = 8'h5a == r_count_76_io_out ? io_r_90_b : _GEN_15589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15591 = 8'h5b == r_count_76_io_out ? io_r_91_b : _GEN_15590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15592 = 8'h5c == r_count_76_io_out ? io_r_92_b : _GEN_15591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15593 = 8'h5d == r_count_76_io_out ? io_r_93_b : _GEN_15592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15594 = 8'h5e == r_count_76_io_out ? io_r_94_b : _GEN_15593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15595 = 8'h5f == r_count_76_io_out ? io_r_95_b : _GEN_15594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15596 = 8'h60 == r_count_76_io_out ? io_r_96_b : _GEN_15595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15597 = 8'h61 == r_count_76_io_out ? io_r_97_b : _GEN_15596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15598 = 8'h62 == r_count_76_io_out ? io_r_98_b : _GEN_15597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15599 = 8'h63 == r_count_76_io_out ? io_r_99_b : _GEN_15598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15600 = 8'h64 == r_count_76_io_out ? io_r_100_b : _GEN_15599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15601 = 8'h65 == r_count_76_io_out ? io_r_101_b : _GEN_15600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15602 = 8'h66 == r_count_76_io_out ? io_r_102_b : _GEN_15601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15603 = 8'h67 == r_count_76_io_out ? io_r_103_b : _GEN_15602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15604 = 8'h68 == r_count_76_io_out ? io_r_104_b : _GEN_15603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15605 = 8'h69 == r_count_76_io_out ? io_r_105_b : _GEN_15604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15606 = 8'h6a == r_count_76_io_out ? io_r_106_b : _GEN_15605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15607 = 8'h6b == r_count_76_io_out ? io_r_107_b : _GEN_15606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15608 = 8'h6c == r_count_76_io_out ? io_r_108_b : _GEN_15607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15609 = 8'h6d == r_count_76_io_out ? io_r_109_b : _GEN_15608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15610 = 8'h6e == r_count_76_io_out ? io_r_110_b : _GEN_15609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15611 = 8'h6f == r_count_76_io_out ? io_r_111_b : _GEN_15610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15612 = 8'h70 == r_count_76_io_out ? io_r_112_b : _GEN_15611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15613 = 8'h71 == r_count_76_io_out ? io_r_113_b : _GEN_15612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15614 = 8'h72 == r_count_76_io_out ? io_r_114_b : _GEN_15613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15615 = 8'h73 == r_count_76_io_out ? io_r_115_b : _GEN_15614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15616 = 8'h74 == r_count_76_io_out ? io_r_116_b : _GEN_15615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15617 = 8'h75 == r_count_76_io_out ? io_r_117_b : _GEN_15616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15618 = 8'h76 == r_count_76_io_out ? io_r_118_b : _GEN_15617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15619 = 8'h77 == r_count_76_io_out ? io_r_119_b : _GEN_15618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15620 = 8'h78 == r_count_76_io_out ? io_r_120_b : _GEN_15619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15621 = 8'h79 == r_count_76_io_out ? io_r_121_b : _GEN_15620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15622 = 8'h7a == r_count_76_io_out ? io_r_122_b : _GEN_15621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15623 = 8'h7b == r_count_76_io_out ? io_r_123_b : _GEN_15622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15624 = 8'h7c == r_count_76_io_out ? io_r_124_b : _GEN_15623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15625 = 8'h7d == r_count_76_io_out ? io_r_125_b : _GEN_15624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15626 = 8'h7e == r_count_76_io_out ? io_r_126_b : _GEN_15625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15627 = 8'h7f == r_count_76_io_out ? io_r_127_b : _GEN_15626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15628 = 8'h80 == r_count_76_io_out ? io_r_128_b : _GEN_15627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15629 = 8'h81 == r_count_76_io_out ? io_r_129_b : _GEN_15628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15630 = 8'h82 == r_count_76_io_out ? io_r_130_b : _GEN_15629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15631 = 8'h83 == r_count_76_io_out ? io_r_131_b : _GEN_15630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15632 = 8'h84 == r_count_76_io_out ? io_r_132_b : _GEN_15631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15633 = 8'h85 == r_count_76_io_out ? io_r_133_b : _GEN_15632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15634 = 8'h86 == r_count_76_io_out ? io_r_134_b : _GEN_15633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15635 = 8'h87 == r_count_76_io_out ? io_r_135_b : _GEN_15634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15636 = 8'h88 == r_count_76_io_out ? io_r_136_b : _GEN_15635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15637 = 8'h89 == r_count_76_io_out ? io_r_137_b : _GEN_15636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15638 = 8'h8a == r_count_76_io_out ? io_r_138_b : _GEN_15637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15639 = 8'h8b == r_count_76_io_out ? io_r_139_b : _GEN_15638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15640 = 8'h8c == r_count_76_io_out ? io_r_140_b : _GEN_15639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15641 = 8'h8d == r_count_76_io_out ? io_r_141_b : _GEN_15640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15642 = 8'h8e == r_count_76_io_out ? io_r_142_b : _GEN_15641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15643 = 8'h8f == r_count_76_io_out ? io_r_143_b : _GEN_15642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15644 = 8'h90 == r_count_76_io_out ? io_r_144_b : _GEN_15643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15645 = 8'h91 == r_count_76_io_out ? io_r_145_b : _GEN_15644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15646 = 8'h92 == r_count_76_io_out ? io_r_146_b : _GEN_15645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15647 = 8'h93 == r_count_76_io_out ? io_r_147_b : _GEN_15646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15648 = 8'h94 == r_count_76_io_out ? io_r_148_b : _GEN_15647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15649 = 8'h95 == r_count_76_io_out ? io_r_149_b : _GEN_15648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15650 = 8'h96 == r_count_76_io_out ? io_r_150_b : _GEN_15649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15651 = 8'h97 == r_count_76_io_out ? io_r_151_b : _GEN_15650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15652 = 8'h98 == r_count_76_io_out ? io_r_152_b : _GEN_15651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15653 = 8'h99 == r_count_76_io_out ? io_r_153_b : _GEN_15652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15654 = 8'h9a == r_count_76_io_out ? io_r_154_b : _GEN_15653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15655 = 8'h9b == r_count_76_io_out ? io_r_155_b : _GEN_15654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15656 = 8'h9c == r_count_76_io_out ? io_r_156_b : _GEN_15655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15657 = 8'h9d == r_count_76_io_out ? io_r_157_b : _GEN_15656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15658 = 8'h9e == r_count_76_io_out ? io_r_158_b : _GEN_15657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15659 = 8'h9f == r_count_76_io_out ? io_r_159_b : _GEN_15658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15660 = 8'ha0 == r_count_76_io_out ? io_r_160_b : _GEN_15659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15661 = 8'ha1 == r_count_76_io_out ? io_r_161_b : _GEN_15660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15662 = 8'ha2 == r_count_76_io_out ? io_r_162_b : _GEN_15661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15663 = 8'ha3 == r_count_76_io_out ? io_r_163_b : _GEN_15662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15664 = 8'ha4 == r_count_76_io_out ? io_r_164_b : _GEN_15663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15665 = 8'ha5 == r_count_76_io_out ? io_r_165_b : _GEN_15664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15666 = 8'ha6 == r_count_76_io_out ? io_r_166_b : _GEN_15665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15667 = 8'ha7 == r_count_76_io_out ? io_r_167_b : _GEN_15666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15668 = 8'ha8 == r_count_76_io_out ? io_r_168_b : _GEN_15667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15669 = 8'ha9 == r_count_76_io_out ? io_r_169_b : _GEN_15668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15670 = 8'haa == r_count_76_io_out ? io_r_170_b : _GEN_15669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15671 = 8'hab == r_count_76_io_out ? io_r_171_b : _GEN_15670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15672 = 8'hac == r_count_76_io_out ? io_r_172_b : _GEN_15671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15673 = 8'had == r_count_76_io_out ? io_r_173_b : _GEN_15672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15674 = 8'hae == r_count_76_io_out ? io_r_174_b : _GEN_15673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15675 = 8'haf == r_count_76_io_out ? io_r_175_b : _GEN_15674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15676 = 8'hb0 == r_count_76_io_out ? io_r_176_b : _GEN_15675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15677 = 8'hb1 == r_count_76_io_out ? io_r_177_b : _GEN_15676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15678 = 8'hb2 == r_count_76_io_out ? io_r_178_b : _GEN_15677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15679 = 8'hb3 == r_count_76_io_out ? io_r_179_b : _GEN_15678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15680 = 8'hb4 == r_count_76_io_out ? io_r_180_b : _GEN_15679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15681 = 8'hb5 == r_count_76_io_out ? io_r_181_b : _GEN_15680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15682 = 8'hb6 == r_count_76_io_out ? io_r_182_b : _GEN_15681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15683 = 8'hb7 == r_count_76_io_out ? io_r_183_b : _GEN_15682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15684 = 8'hb8 == r_count_76_io_out ? io_r_184_b : _GEN_15683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15685 = 8'hb9 == r_count_76_io_out ? io_r_185_b : _GEN_15684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15686 = 8'hba == r_count_76_io_out ? io_r_186_b : _GEN_15685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15687 = 8'hbb == r_count_76_io_out ? io_r_187_b : _GEN_15686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15688 = 8'hbc == r_count_76_io_out ? io_r_188_b : _GEN_15687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15689 = 8'hbd == r_count_76_io_out ? io_r_189_b : _GEN_15688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15690 = 8'hbe == r_count_76_io_out ? io_r_190_b : _GEN_15689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15691 = 8'hbf == r_count_76_io_out ? io_r_191_b : _GEN_15690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15692 = 8'hc0 == r_count_76_io_out ? io_r_192_b : _GEN_15691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15693 = 8'hc1 == r_count_76_io_out ? io_r_193_b : _GEN_15692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15694 = 8'hc2 == r_count_76_io_out ? io_r_194_b : _GEN_15693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15695 = 8'hc3 == r_count_76_io_out ? io_r_195_b : _GEN_15694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15696 = 8'hc4 == r_count_76_io_out ? io_r_196_b : _GEN_15695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15697 = 8'hc5 == r_count_76_io_out ? io_r_197_b : _GEN_15696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15698 = 8'hc6 == r_count_76_io_out ? io_r_198_b : _GEN_15697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15701 = 8'h1 == r_count_77_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15702 = 8'h2 == r_count_77_io_out ? io_r_2_b : _GEN_15701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15703 = 8'h3 == r_count_77_io_out ? io_r_3_b : _GEN_15702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15704 = 8'h4 == r_count_77_io_out ? io_r_4_b : _GEN_15703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15705 = 8'h5 == r_count_77_io_out ? io_r_5_b : _GEN_15704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15706 = 8'h6 == r_count_77_io_out ? io_r_6_b : _GEN_15705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15707 = 8'h7 == r_count_77_io_out ? io_r_7_b : _GEN_15706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15708 = 8'h8 == r_count_77_io_out ? io_r_8_b : _GEN_15707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15709 = 8'h9 == r_count_77_io_out ? io_r_9_b : _GEN_15708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15710 = 8'ha == r_count_77_io_out ? io_r_10_b : _GEN_15709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15711 = 8'hb == r_count_77_io_out ? io_r_11_b : _GEN_15710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15712 = 8'hc == r_count_77_io_out ? io_r_12_b : _GEN_15711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15713 = 8'hd == r_count_77_io_out ? io_r_13_b : _GEN_15712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15714 = 8'he == r_count_77_io_out ? io_r_14_b : _GEN_15713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15715 = 8'hf == r_count_77_io_out ? io_r_15_b : _GEN_15714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15716 = 8'h10 == r_count_77_io_out ? io_r_16_b : _GEN_15715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15717 = 8'h11 == r_count_77_io_out ? io_r_17_b : _GEN_15716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15718 = 8'h12 == r_count_77_io_out ? io_r_18_b : _GEN_15717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15719 = 8'h13 == r_count_77_io_out ? io_r_19_b : _GEN_15718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15720 = 8'h14 == r_count_77_io_out ? io_r_20_b : _GEN_15719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15721 = 8'h15 == r_count_77_io_out ? io_r_21_b : _GEN_15720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15722 = 8'h16 == r_count_77_io_out ? io_r_22_b : _GEN_15721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15723 = 8'h17 == r_count_77_io_out ? io_r_23_b : _GEN_15722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15724 = 8'h18 == r_count_77_io_out ? io_r_24_b : _GEN_15723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15725 = 8'h19 == r_count_77_io_out ? io_r_25_b : _GEN_15724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15726 = 8'h1a == r_count_77_io_out ? io_r_26_b : _GEN_15725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15727 = 8'h1b == r_count_77_io_out ? io_r_27_b : _GEN_15726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15728 = 8'h1c == r_count_77_io_out ? io_r_28_b : _GEN_15727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15729 = 8'h1d == r_count_77_io_out ? io_r_29_b : _GEN_15728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15730 = 8'h1e == r_count_77_io_out ? io_r_30_b : _GEN_15729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15731 = 8'h1f == r_count_77_io_out ? io_r_31_b : _GEN_15730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15732 = 8'h20 == r_count_77_io_out ? io_r_32_b : _GEN_15731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15733 = 8'h21 == r_count_77_io_out ? io_r_33_b : _GEN_15732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15734 = 8'h22 == r_count_77_io_out ? io_r_34_b : _GEN_15733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15735 = 8'h23 == r_count_77_io_out ? io_r_35_b : _GEN_15734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15736 = 8'h24 == r_count_77_io_out ? io_r_36_b : _GEN_15735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15737 = 8'h25 == r_count_77_io_out ? io_r_37_b : _GEN_15736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15738 = 8'h26 == r_count_77_io_out ? io_r_38_b : _GEN_15737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15739 = 8'h27 == r_count_77_io_out ? io_r_39_b : _GEN_15738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15740 = 8'h28 == r_count_77_io_out ? io_r_40_b : _GEN_15739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15741 = 8'h29 == r_count_77_io_out ? io_r_41_b : _GEN_15740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15742 = 8'h2a == r_count_77_io_out ? io_r_42_b : _GEN_15741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15743 = 8'h2b == r_count_77_io_out ? io_r_43_b : _GEN_15742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15744 = 8'h2c == r_count_77_io_out ? io_r_44_b : _GEN_15743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15745 = 8'h2d == r_count_77_io_out ? io_r_45_b : _GEN_15744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15746 = 8'h2e == r_count_77_io_out ? io_r_46_b : _GEN_15745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15747 = 8'h2f == r_count_77_io_out ? io_r_47_b : _GEN_15746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15748 = 8'h30 == r_count_77_io_out ? io_r_48_b : _GEN_15747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15749 = 8'h31 == r_count_77_io_out ? io_r_49_b : _GEN_15748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15750 = 8'h32 == r_count_77_io_out ? io_r_50_b : _GEN_15749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15751 = 8'h33 == r_count_77_io_out ? io_r_51_b : _GEN_15750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15752 = 8'h34 == r_count_77_io_out ? io_r_52_b : _GEN_15751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15753 = 8'h35 == r_count_77_io_out ? io_r_53_b : _GEN_15752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15754 = 8'h36 == r_count_77_io_out ? io_r_54_b : _GEN_15753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15755 = 8'h37 == r_count_77_io_out ? io_r_55_b : _GEN_15754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15756 = 8'h38 == r_count_77_io_out ? io_r_56_b : _GEN_15755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15757 = 8'h39 == r_count_77_io_out ? io_r_57_b : _GEN_15756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15758 = 8'h3a == r_count_77_io_out ? io_r_58_b : _GEN_15757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15759 = 8'h3b == r_count_77_io_out ? io_r_59_b : _GEN_15758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15760 = 8'h3c == r_count_77_io_out ? io_r_60_b : _GEN_15759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15761 = 8'h3d == r_count_77_io_out ? io_r_61_b : _GEN_15760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15762 = 8'h3e == r_count_77_io_out ? io_r_62_b : _GEN_15761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15763 = 8'h3f == r_count_77_io_out ? io_r_63_b : _GEN_15762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15764 = 8'h40 == r_count_77_io_out ? io_r_64_b : _GEN_15763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15765 = 8'h41 == r_count_77_io_out ? io_r_65_b : _GEN_15764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15766 = 8'h42 == r_count_77_io_out ? io_r_66_b : _GEN_15765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15767 = 8'h43 == r_count_77_io_out ? io_r_67_b : _GEN_15766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15768 = 8'h44 == r_count_77_io_out ? io_r_68_b : _GEN_15767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15769 = 8'h45 == r_count_77_io_out ? io_r_69_b : _GEN_15768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15770 = 8'h46 == r_count_77_io_out ? io_r_70_b : _GEN_15769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15771 = 8'h47 == r_count_77_io_out ? io_r_71_b : _GEN_15770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15772 = 8'h48 == r_count_77_io_out ? io_r_72_b : _GEN_15771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15773 = 8'h49 == r_count_77_io_out ? io_r_73_b : _GEN_15772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15774 = 8'h4a == r_count_77_io_out ? io_r_74_b : _GEN_15773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15775 = 8'h4b == r_count_77_io_out ? io_r_75_b : _GEN_15774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15776 = 8'h4c == r_count_77_io_out ? io_r_76_b : _GEN_15775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15777 = 8'h4d == r_count_77_io_out ? io_r_77_b : _GEN_15776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15778 = 8'h4e == r_count_77_io_out ? io_r_78_b : _GEN_15777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15779 = 8'h4f == r_count_77_io_out ? io_r_79_b : _GEN_15778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15780 = 8'h50 == r_count_77_io_out ? io_r_80_b : _GEN_15779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15781 = 8'h51 == r_count_77_io_out ? io_r_81_b : _GEN_15780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15782 = 8'h52 == r_count_77_io_out ? io_r_82_b : _GEN_15781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15783 = 8'h53 == r_count_77_io_out ? io_r_83_b : _GEN_15782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15784 = 8'h54 == r_count_77_io_out ? io_r_84_b : _GEN_15783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15785 = 8'h55 == r_count_77_io_out ? io_r_85_b : _GEN_15784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15786 = 8'h56 == r_count_77_io_out ? io_r_86_b : _GEN_15785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15787 = 8'h57 == r_count_77_io_out ? io_r_87_b : _GEN_15786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15788 = 8'h58 == r_count_77_io_out ? io_r_88_b : _GEN_15787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15789 = 8'h59 == r_count_77_io_out ? io_r_89_b : _GEN_15788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15790 = 8'h5a == r_count_77_io_out ? io_r_90_b : _GEN_15789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15791 = 8'h5b == r_count_77_io_out ? io_r_91_b : _GEN_15790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15792 = 8'h5c == r_count_77_io_out ? io_r_92_b : _GEN_15791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15793 = 8'h5d == r_count_77_io_out ? io_r_93_b : _GEN_15792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15794 = 8'h5e == r_count_77_io_out ? io_r_94_b : _GEN_15793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15795 = 8'h5f == r_count_77_io_out ? io_r_95_b : _GEN_15794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15796 = 8'h60 == r_count_77_io_out ? io_r_96_b : _GEN_15795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15797 = 8'h61 == r_count_77_io_out ? io_r_97_b : _GEN_15796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15798 = 8'h62 == r_count_77_io_out ? io_r_98_b : _GEN_15797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15799 = 8'h63 == r_count_77_io_out ? io_r_99_b : _GEN_15798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15800 = 8'h64 == r_count_77_io_out ? io_r_100_b : _GEN_15799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15801 = 8'h65 == r_count_77_io_out ? io_r_101_b : _GEN_15800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15802 = 8'h66 == r_count_77_io_out ? io_r_102_b : _GEN_15801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15803 = 8'h67 == r_count_77_io_out ? io_r_103_b : _GEN_15802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15804 = 8'h68 == r_count_77_io_out ? io_r_104_b : _GEN_15803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15805 = 8'h69 == r_count_77_io_out ? io_r_105_b : _GEN_15804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15806 = 8'h6a == r_count_77_io_out ? io_r_106_b : _GEN_15805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15807 = 8'h6b == r_count_77_io_out ? io_r_107_b : _GEN_15806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15808 = 8'h6c == r_count_77_io_out ? io_r_108_b : _GEN_15807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15809 = 8'h6d == r_count_77_io_out ? io_r_109_b : _GEN_15808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15810 = 8'h6e == r_count_77_io_out ? io_r_110_b : _GEN_15809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15811 = 8'h6f == r_count_77_io_out ? io_r_111_b : _GEN_15810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15812 = 8'h70 == r_count_77_io_out ? io_r_112_b : _GEN_15811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15813 = 8'h71 == r_count_77_io_out ? io_r_113_b : _GEN_15812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15814 = 8'h72 == r_count_77_io_out ? io_r_114_b : _GEN_15813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15815 = 8'h73 == r_count_77_io_out ? io_r_115_b : _GEN_15814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15816 = 8'h74 == r_count_77_io_out ? io_r_116_b : _GEN_15815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15817 = 8'h75 == r_count_77_io_out ? io_r_117_b : _GEN_15816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15818 = 8'h76 == r_count_77_io_out ? io_r_118_b : _GEN_15817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15819 = 8'h77 == r_count_77_io_out ? io_r_119_b : _GEN_15818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15820 = 8'h78 == r_count_77_io_out ? io_r_120_b : _GEN_15819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15821 = 8'h79 == r_count_77_io_out ? io_r_121_b : _GEN_15820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15822 = 8'h7a == r_count_77_io_out ? io_r_122_b : _GEN_15821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15823 = 8'h7b == r_count_77_io_out ? io_r_123_b : _GEN_15822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15824 = 8'h7c == r_count_77_io_out ? io_r_124_b : _GEN_15823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15825 = 8'h7d == r_count_77_io_out ? io_r_125_b : _GEN_15824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15826 = 8'h7e == r_count_77_io_out ? io_r_126_b : _GEN_15825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15827 = 8'h7f == r_count_77_io_out ? io_r_127_b : _GEN_15826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15828 = 8'h80 == r_count_77_io_out ? io_r_128_b : _GEN_15827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15829 = 8'h81 == r_count_77_io_out ? io_r_129_b : _GEN_15828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15830 = 8'h82 == r_count_77_io_out ? io_r_130_b : _GEN_15829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15831 = 8'h83 == r_count_77_io_out ? io_r_131_b : _GEN_15830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15832 = 8'h84 == r_count_77_io_out ? io_r_132_b : _GEN_15831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15833 = 8'h85 == r_count_77_io_out ? io_r_133_b : _GEN_15832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15834 = 8'h86 == r_count_77_io_out ? io_r_134_b : _GEN_15833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15835 = 8'h87 == r_count_77_io_out ? io_r_135_b : _GEN_15834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15836 = 8'h88 == r_count_77_io_out ? io_r_136_b : _GEN_15835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15837 = 8'h89 == r_count_77_io_out ? io_r_137_b : _GEN_15836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15838 = 8'h8a == r_count_77_io_out ? io_r_138_b : _GEN_15837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15839 = 8'h8b == r_count_77_io_out ? io_r_139_b : _GEN_15838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15840 = 8'h8c == r_count_77_io_out ? io_r_140_b : _GEN_15839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15841 = 8'h8d == r_count_77_io_out ? io_r_141_b : _GEN_15840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15842 = 8'h8e == r_count_77_io_out ? io_r_142_b : _GEN_15841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15843 = 8'h8f == r_count_77_io_out ? io_r_143_b : _GEN_15842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15844 = 8'h90 == r_count_77_io_out ? io_r_144_b : _GEN_15843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15845 = 8'h91 == r_count_77_io_out ? io_r_145_b : _GEN_15844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15846 = 8'h92 == r_count_77_io_out ? io_r_146_b : _GEN_15845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15847 = 8'h93 == r_count_77_io_out ? io_r_147_b : _GEN_15846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15848 = 8'h94 == r_count_77_io_out ? io_r_148_b : _GEN_15847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15849 = 8'h95 == r_count_77_io_out ? io_r_149_b : _GEN_15848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15850 = 8'h96 == r_count_77_io_out ? io_r_150_b : _GEN_15849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15851 = 8'h97 == r_count_77_io_out ? io_r_151_b : _GEN_15850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15852 = 8'h98 == r_count_77_io_out ? io_r_152_b : _GEN_15851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15853 = 8'h99 == r_count_77_io_out ? io_r_153_b : _GEN_15852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15854 = 8'h9a == r_count_77_io_out ? io_r_154_b : _GEN_15853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15855 = 8'h9b == r_count_77_io_out ? io_r_155_b : _GEN_15854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15856 = 8'h9c == r_count_77_io_out ? io_r_156_b : _GEN_15855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15857 = 8'h9d == r_count_77_io_out ? io_r_157_b : _GEN_15856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15858 = 8'h9e == r_count_77_io_out ? io_r_158_b : _GEN_15857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15859 = 8'h9f == r_count_77_io_out ? io_r_159_b : _GEN_15858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15860 = 8'ha0 == r_count_77_io_out ? io_r_160_b : _GEN_15859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15861 = 8'ha1 == r_count_77_io_out ? io_r_161_b : _GEN_15860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15862 = 8'ha2 == r_count_77_io_out ? io_r_162_b : _GEN_15861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15863 = 8'ha3 == r_count_77_io_out ? io_r_163_b : _GEN_15862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15864 = 8'ha4 == r_count_77_io_out ? io_r_164_b : _GEN_15863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15865 = 8'ha5 == r_count_77_io_out ? io_r_165_b : _GEN_15864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15866 = 8'ha6 == r_count_77_io_out ? io_r_166_b : _GEN_15865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15867 = 8'ha7 == r_count_77_io_out ? io_r_167_b : _GEN_15866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15868 = 8'ha8 == r_count_77_io_out ? io_r_168_b : _GEN_15867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15869 = 8'ha9 == r_count_77_io_out ? io_r_169_b : _GEN_15868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15870 = 8'haa == r_count_77_io_out ? io_r_170_b : _GEN_15869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15871 = 8'hab == r_count_77_io_out ? io_r_171_b : _GEN_15870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15872 = 8'hac == r_count_77_io_out ? io_r_172_b : _GEN_15871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15873 = 8'had == r_count_77_io_out ? io_r_173_b : _GEN_15872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15874 = 8'hae == r_count_77_io_out ? io_r_174_b : _GEN_15873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15875 = 8'haf == r_count_77_io_out ? io_r_175_b : _GEN_15874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15876 = 8'hb0 == r_count_77_io_out ? io_r_176_b : _GEN_15875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15877 = 8'hb1 == r_count_77_io_out ? io_r_177_b : _GEN_15876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15878 = 8'hb2 == r_count_77_io_out ? io_r_178_b : _GEN_15877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15879 = 8'hb3 == r_count_77_io_out ? io_r_179_b : _GEN_15878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15880 = 8'hb4 == r_count_77_io_out ? io_r_180_b : _GEN_15879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15881 = 8'hb5 == r_count_77_io_out ? io_r_181_b : _GEN_15880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15882 = 8'hb6 == r_count_77_io_out ? io_r_182_b : _GEN_15881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15883 = 8'hb7 == r_count_77_io_out ? io_r_183_b : _GEN_15882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15884 = 8'hb8 == r_count_77_io_out ? io_r_184_b : _GEN_15883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15885 = 8'hb9 == r_count_77_io_out ? io_r_185_b : _GEN_15884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15886 = 8'hba == r_count_77_io_out ? io_r_186_b : _GEN_15885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15887 = 8'hbb == r_count_77_io_out ? io_r_187_b : _GEN_15886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15888 = 8'hbc == r_count_77_io_out ? io_r_188_b : _GEN_15887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15889 = 8'hbd == r_count_77_io_out ? io_r_189_b : _GEN_15888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15890 = 8'hbe == r_count_77_io_out ? io_r_190_b : _GEN_15889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15891 = 8'hbf == r_count_77_io_out ? io_r_191_b : _GEN_15890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15892 = 8'hc0 == r_count_77_io_out ? io_r_192_b : _GEN_15891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15893 = 8'hc1 == r_count_77_io_out ? io_r_193_b : _GEN_15892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15894 = 8'hc2 == r_count_77_io_out ? io_r_194_b : _GEN_15893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15895 = 8'hc3 == r_count_77_io_out ? io_r_195_b : _GEN_15894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15896 = 8'hc4 == r_count_77_io_out ? io_r_196_b : _GEN_15895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15897 = 8'hc5 == r_count_77_io_out ? io_r_197_b : _GEN_15896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15898 = 8'hc6 == r_count_77_io_out ? io_r_198_b : _GEN_15897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15901 = 8'h1 == r_count_78_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15902 = 8'h2 == r_count_78_io_out ? io_r_2_b : _GEN_15901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15903 = 8'h3 == r_count_78_io_out ? io_r_3_b : _GEN_15902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15904 = 8'h4 == r_count_78_io_out ? io_r_4_b : _GEN_15903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15905 = 8'h5 == r_count_78_io_out ? io_r_5_b : _GEN_15904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15906 = 8'h6 == r_count_78_io_out ? io_r_6_b : _GEN_15905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15907 = 8'h7 == r_count_78_io_out ? io_r_7_b : _GEN_15906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15908 = 8'h8 == r_count_78_io_out ? io_r_8_b : _GEN_15907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15909 = 8'h9 == r_count_78_io_out ? io_r_9_b : _GEN_15908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15910 = 8'ha == r_count_78_io_out ? io_r_10_b : _GEN_15909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15911 = 8'hb == r_count_78_io_out ? io_r_11_b : _GEN_15910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15912 = 8'hc == r_count_78_io_out ? io_r_12_b : _GEN_15911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15913 = 8'hd == r_count_78_io_out ? io_r_13_b : _GEN_15912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15914 = 8'he == r_count_78_io_out ? io_r_14_b : _GEN_15913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15915 = 8'hf == r_count_78_io_out ? io_r_15_b : _GEN_15914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15916 = 8'h10 == r_count_78_io_out ? io_r_16_b : _GEN_15915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15917 = 8'h11 == r_count_78_io_out ? io_r_17_b : _GEN_15916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15918 = 8'h12 == r_count_78_io_out ? io_r_18_b : _GEN_15917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15919 = 8'h13 == r_count_78_io_out ? io_r_19_b : _GEN_15918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15920 = 8'h14 == r_count_78_io_out ? io_r_20_b : _GEN_15919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15921 = 8'h15 == r_count_78_io_out ? io_r_21_b : _GEN_15920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15922 = 8'h16 == r_count_78_io_out ? io_r_22_b : _GEN_15921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15923 = 8'h17 == r_count_78_io_out ? io_r_23_b : _GEN_15922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15924 = 8'h18 == r_count_78_io_out ? io_r_24_b : _GEN_15923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15925 = 8'h19 == r_count_78_io_out ? io_r_25_b : _GEN_15924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15926 = 8'h1a == r_count_78_io_out ? io_r_26_b : _GEN_15925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15927 = 8'h1b == r_count_78_io_out ? io_r_27_b : _GEN_15926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15928 = 8'h1c == r_count_78_io_out ? io_r_28_b : _GEN_15927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15929 = 8'h1d == r_count_78_io_out ? io_r_29_b : _GEN_15928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15930 = 8'h1e == r_count_78_io_out ? io_r_30_b : _GEN_15929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15931 = 8'h1f == r_count_78_io_out ? io_r_31_b : _GEN_15930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15932 = 8'h20 == r_count_78_io_out ? io_r_32_b : _GEN_15931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15933 = 8'h21 == r_count_78_io_out ? io_r_33_b : _GEN_15932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15934 = 8'h22 == r_count_78_io_out ? io_r_34_b : _GEN_15933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15935 = 8'h23 == r_count_78_io_out ? io_r_35_b : _GEN_15934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15936 = 8'h24 == r_count_78_io_out ? io_r_36_b : _GEN_15935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15937 = 8'h25 == r_count_78_io_out ? io_r_37_b : _GEN_15936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15938 = 8'h26 == r_count_78_io_out ? io_r_38_b : _GEN_15937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15939 = 8'h27 == r_count_78_io_out ? io_r_39_b : _GEN_15938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15940 = 8'h28 == r_count_78_io_out ? io_r_40_b : _GEN_15939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15941 = 8'h29 == r_count_78_io_out ? io_r_41_b : _GEN_15940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15942 = 8'h2a == r_count_78_io_out ? io_r_42_b : _GEN_15941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15943 = 8'h2b == r_count_78_io_out ? io_r_43_b : _GEN_15942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15944 = 8'h2c == r_count_78_io_out ? io_r_44_b : _GEN_15943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15945 = 8'h2d == r_count_78_io_out ? io_r_45_b : _GEN_15944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15946 = 8'h2e == r_count_78_io_out ? io_r_46_b : _GEN_15945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15947 = 8'h2f == r_count_78_io_out ? io_r_47_b : _GEN_15946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15948 = 8'h30 == r_count_78_io_out ? io_r_48_b : _GEN_15947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15949 = 8'h31 == r_count_78_io_out ? io_r_49_b : _GEN_15948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15950 = 8'h32 == r_count_78_io_out ? io_r_50_b : _GEN_15949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15951 = 8'h33 == r_count_78_io_out ? io_r_51_b : _GEN_15950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15952 = 8'h34 == r_count_78_io_out ? io_r_52_b : _GEN_15951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15953 = 8'h35 == r_count_78_io_out ? io_r_53_b : _GEN_15952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15954 = 8'h36 == r_count_78_io_out ? io_r_54_b : _GEN_15953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15955 = 8'h37 == r_count_78_io_out ? io_r_55_b : _GEN_15954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15956 = 8'h38 == r_count_78_io_out ? io_r_56_b : _GEN_15955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15957 = 8'h39 == r_count_78_io_out ? io_r_57_b : _GEN_15956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15958 = 8'h3a == r_count_78_io_out ? io_r_58_b : _GEN_15957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15959 = 8'h3b == r_count_78_io_out ? io_r_59_b : _GEN_15958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15960 = 8'h3c == r_count_78_io_out ? io_r_60_b : _GEN_15959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15961 = 8'h3d == r_count_78_io_out ? io_r_61_b : _GEN_15960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15962 = 8'h3e == r_count_78_io_out ? io_r_62_b : _GEN_15961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15963 = 8'h3f == r_count_78_io_out ? io_r_63_b : _GEN_15962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15964 = 8'h40 == r_count_78_io_out ? io_r_64_b : _GEN_15963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15965 = 8'h41 == r_count_78_io_out ? io_r_65_b : _GEN_15964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15966 = 8'h42 == r_count_78_io_out ? io_r_66_b : _GEN_15965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15967 = 8'h43 == r_count_78_io_out ? io_r_67_b : _GEN_15966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15968 = 8'h44 == r_count_78_io_out ? io_r_68_b : _GEN_15967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15969 = 8'h45 == r_count_78_io_out ? io_r_69_b : _GEN_15968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15970 = 8'h46 == r_count_78_io_out ? io_r_70_b : _GEN_15969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15971 = 8'h47 == r_count_78_io_out ? io_r_71_b : _GEN_15970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15972 = 8'h48 == r_count_78_io_out ? io_r_72_b : _GEN_15971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15973 = 8'h49 == r_count_78_io_out ? io_r_73_b : _GEN_15972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15974 = 8'h4a == r_count_78_io_out ? io_r_74_b : _GEN_15973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15975 = 8'h4b == r_count_78_io_out ? io_r_75_b : _GEN_15974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15976 = 8'h4c == r_count_78_io_out ? io_r_76_b : _GEN_15975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15977 = 8'h4d == r_count_78_io_out ? io_r_77_b : _GEN_15976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15978 = 8'h4e == r_count_78_io_out ? io_r_78_b : _GEN_15977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15979 = 8'h4f == r_count_78_io_out ? io_r_79_b : _GEN_15978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15980 = 8'h50 == r_count_78_io_out ? io_r_80_b : _GEN_15979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15981 = 8'h51 == r_count_78_io_out ? io_r_81_b : _GEN_15980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15982 = 8'h52 == r_count_78_io_out ? io_r_82_b : _GEN_15981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15983 = 8'h53 == r_count_78_io_out ? io_r_83_b : _GEN_15982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15984 = 8'h54 == r_count_78_io_out ? io_r_84_b : _GEN_15983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15985 = 8'h55 == r_count_78_io_out ? io_r_85_b : _GEN_15984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15986 = 8'h56 == r_count_78_io_out ? io_r_86_b : _GEN_15985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15987 = 8'h57 == r_count_78_io_out ? io_r_87_b : _GEN_15986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15988 = 8'h58 == r_count_78_io_out ? io_r_88_b : _GEN_15987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15989 = 8'h59 == r_count_78_io_out ? io_r_89_b : _GEN_15988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15990 = 8'h5a == r_count_78_io_out ? io_r_90_b : _GEN_15989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15991 = 8'h5b == r_count_78_io_out ? io_r_91_b : _GEN_15990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15992 = 8'h5c == r_count_78_io_out ? io_r_92_b : _GEN_15991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15993 = 8'h5d == r_count_78_io_out ? io_r_93_b : _GEN_15992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15994 = 8'h5e == r_count_78_io_out ? io_r_94_b : _GEN_15993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15995 = 8'h5f == r_count_78_io_out ? io_r_95_b : _GEN_15994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15996 = 8'h60 == r_count_78_io_out ? io_r_96_b : _GEN_15995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15997 = 8'h61 == r_count_78_io_out ? io_r_97_b : _GEN_15996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15998 = 8'h62 == r_count_78_io_out ? io_r_98_b : _GEN_15997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_15999 = 8'h63 == r_count_78_io_out ? io_r_99_b : _GEN_15998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16000 = 8'h64 == r_count_78_io_out ? io_r_100_b : _GEN_15999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16001 = 8'h65 == r_count_78_io_out ? io_r_101_b : _GEN_16000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16002 = 8'h66 == r_count_78_io_out ? io_r_102_b : _GEN_16001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16003 = 8'h67 == r_count_78_io_out ? io_r_103_b : _GEN_16002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16004 = 8'h68 == r_count_78_io_out ? io_r_104_b : _GEN_16003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16005 = 8'h69 == r_count_78_io_out ? io_r_105_b : _GEN_16004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16006 = 8'h6a == r_count_78_io_out ? io_r_106_b : _GEN_16005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16007 = 8'h6b == r_count_78_io_out ? io_r_107_b : _GEN_16006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16008 = 8'h6c == r_count_78_io_out ? io_r_108_b : _GEN_16007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16009 = 8'h6d == r_count_78_io_out ? io_r_109_b : _GEN_16008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16010 = 8'h6e == r_count_78_io_out ? io_r_110_b : _GEN_16009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16011 = 8'h6f == r_count_78_io_out ? io_r_111_b : _GEN_16010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16012 = 8'h70 == r_count_78_io_out ? io_r_112_b : _GEN_16011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16013 = 8'h71 == r_count_78_io_out ? io_r_113_b : _GEN_16012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16014 = 8'h72 == r_count_78_io_out ? io_r_114_b : _GEN_16013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16015 = 8'h73 == r_count_78_io_out ? io_r_115_b : _GEN_16014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16016 = 8'h74 == r_count_78_io_out ? io_r_116_b : _GEN_16015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16017 = 8'h75 == r_count_78_io_out ? io_r_117_b : _GEN_16016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16018 = 8'h76 == r_count_78_io_out ? io_r_118_b : _GEN_16017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16019 = 8'h77 == r_count_78_io_out ? io_r_119_b : _GEN_16018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16020 = 8'h78 == r_count_78_io_out ? io_r_120_b : _GEN_16019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16021 = 8'h79 == r_count_78_io_out ? io_r_121_b : _GEN_16020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16022 = 8'h7a == r_count_78_io_out ? io_r_122_b : _GEN_16021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16023 = 8'h7b == r_count_78_io_out ? io_r_123_b : _GEN_16022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16024 = 8'h7c == r_count_78_io_out ? io_r_124_b : _GEN_16023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16025 = 8'h7d == r_count_78_io_out ? io_r_125_b : _GEN_16024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16026 = 8'h7e == r_count_78_io_out ? io_r_126_b : _GEN_16025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16027 = 8'h7f == r_count_78_io_out ? io_r_127_b : _GEN_16026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16028 = 8'h80 == r_count_78_io_out ? io_r_128_b : _GEN_16027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16029 = 8'h81 == r_count_78_io_out ? io_r_129_b : _GEN_16028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16030 = 8'h82 == r_count_78_io_out ? io_r_130_b : _GEN_16029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16031 = 8'h83 == r_count_78_io_out ? io_r_131_b : _GEN_16030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16032 = 8'h84 == r_count_78_io_out ? io_r_132_b : _GEN_16031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16033 = 8'h85 == r_count_78_io_out ? io_r_133_b : _GEN_16032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16034 = 8'h86 == r_count_78_io_out ? io_r_134_b : _GEN_16033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16035 = 8'h87 == r_count_78_io_out ? io_r_135_b : _GEN_16034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16036 = 8'h88 == r_count_78_io_out ? io_r_136_b : _GEN_16035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16037 = 8'h89 == r_count_78_io_out ? io_r_137_b : _GEN_16036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16038 = 8'h8a == r_count_78_io_out ? io_r_138_b : _GEN_16037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16039 = 8'h8b == r_count_78_io_out ? io_r_139_b : _GEN_16038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16040 = 8'h8c == r_count_78_io_out ? io_r_140_b : _GEN_16039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16041 = 8'h8d == r_count_78_io_out ? io_r_141_b : _GEN_16040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16042 = 8'h8e == r_count_78_io_out ? io_r_142_b : _GEN_16041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16043 = 8'h8f == r_count_78_io_out ? io_r_143_b : _GEN_16042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16044 = 8'h90 == r_count_78_io_out ? io_r_144_b : _GEN_16043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16045 = 8'h91 == r_count_78_io_out ? io_r_145_b : _GEN_16044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16046 = 8'h92 == r_count_78_io_out ? io_r_146_b : _GEN_16045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16047 = 8'h93 == r_count_78_io_out ? io_r_147_b : _GEN_16046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16048 = 8'h94 == r_count_78_io_out ? io_r_148_b : _GEN_16047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16049 = 8'h95 == r_count_78_io_out ? io_r_149_b : _GEN_16048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16050 = 8'h96 == r_count_78_io_out ? io_r_150_b : _GEN_16049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16051 = 8'h97 == r_count_78_io_out ? io_r_151_b : _GEN_16050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16052 = 8'h98 == r_count_78_io_out ? io_r_152_b : _GEN_16051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16053 = 8'h99 == r_count_78_io_out ? io_r_153_b : _GEN_16052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16054 = 8'h9a == r_count_78_io_out ? io_r_154_b : _GEN_16053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16055 = 8'h9b == r_count_78_io_out ? io_r_155_b : _GEN_16054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16056 = 8'h9c == r_count_78_io_out ? io_r_156_b : _GEN_16055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16057 = 8'h9d == r_count_78_io_out ? io_r_157_b : _GEN_16056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16058 = 8'h9e == r_count_78_io_out ? io_r_158_b : _GEN_16057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16059 = 8'h9f == r_count_78_io_out ? io_r_159_b : _GEN_16058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16060 = 8'ha0 == r_count_78_io_out ? io_r_160_b : _GEN_16059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16061 = 8'ha1 == r_count_78_io_out ? io_r_161_b : _GEN_16060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16062 = 8'ha2 == r_count_78_io_out ? io_r_162_b : _GEN_16061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16063 = 8'ha3 == r_count_78_io_out ? io_r_163_b : _GEN_16062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16064 = 8'ha4 == r_count_78_io_out ? io_r_164_b : _GEN_16063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16065 = 8'ha5 == r_count_78_io_out ? io_r_165_b : _GEN_16064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16066 = 8'ha6 == r_count_78_io_out ? io_r_166_b : _GEN_16065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16067 = 8'ha7 == r_count_78_io_out ? io_r_167_b : _GEN_16066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16068 = 8'ha8 == r_count_78_io_out ? io_r_168_b : _GEN_16067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16069 = 8'ha9 == r_count_78_io_out ? io_r_169_b : _GEN_16068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16070 = 8'haa == r_count_78_io_out ? io_r_170_b : _GEN_16069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16071 = 8'hab == r_count_78_io_out ? io_r_171_b : _GEN_16070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16072 = 8'hac == r_count_78_io_out ? io_r_172_b : _GEN_16071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16073 = 8'had == r_count_78_io_out ? io_r_173_b : _GEN_16072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16074 = 8'hae == r_count_78_io_out ? io_r_174_b : _GEN_16073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16075 = 8'haf == r_count_78_io_out ? io_r_175_b : _GEN_16074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16076 = 8'hb0 == r_count_78_io_out ? io_r_176_b : _GEN_16075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16077 = 8'hb1 == r_count_78_io_out ? io_r_177_b : _GEN_16076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16078 = 8'hb2 == r_count_78_io_out ? io_r_178_b : _GEN_16077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16079 = 8'hb3 == r_count_78_io_out ? io_r_179_b : _GEN_16078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16080 = 8'hb4 == r_count_78_io_out ? io_r_180_b : _GEN_16079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16081 = 8'hb5 == r_count_78_io_out ? io_r_181_b : _GEN_16080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16082 = 8'hb6 == r_count_78_io_out ? io_r_182_b : _GEN_16081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16083 = 8'hb7 == r_count_78_io_out ? io_r_183_b : _GEN_16082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16084 = 8'hb8 == r_count_78_io_out ? io_r_184_b : _GEN_16083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16085 = 8'hb9 == r_count_78_io_out ? io_r_185_b : _GEN_16084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16086 = 8'hba == r_count_78_io_out ? io_r_186_b : _GEN_16085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16087 = 8'hbb == r_count_78_io_out ? io_r_187_b : _GEN_16086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16088 = 8'hbc == r_count_78_io_out ? io_r_188_b : _GEN_16087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16089 = 8'hbd == r_count_78_io_out ? io_r_189_b : _GEN_16088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16090 = 8'hbe == r_count_78_io_out ? io_r_190_b : _GEN_16089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16091 = 8'hbf == r_count_78_io_out ? io_r_191_b : _GEN_16090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16092 = 8'hc0 == r_count_78_io_out ? io_r_192_b : _GEN_16091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16093 = 8'hc1 == r_count_78_io_out ? io_r_193_b : _GEN_16092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16094 = 8'hc2 == r_count_78_io_out ? io_r_194_b : _GEN_16093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16095 = 8'hc3 == r_count_78_io_out ? io_r_195_b : _GEN_16094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16096 = 8'hc4 == r_count_78_io_out ? io_r_196_b : _GEN_16095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16097 = 8'hc5 == r_count_78_io_out ? io_r_197_b : _GEN_16096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16098 = 8'hc6 == r_count_78_io_out ? io_r_198_b : _GEN_16097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16101 = 8'h1 == r_count_79_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16102 = 8'h2 == r_count_79_io_out ? io_r_2_b : _GEN_16101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16103 = 8'h3 == r_count_79_io_out ? io_r_3_b : _GEN_16102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16104 = 8'h4 == r_count_79_io_out ? io_r_4_b : _GEN_16103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16105 = 8'h5 == r_count_79_io_out ? io_r_5_b : _GEN_16104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16106 = 8'h6 == r_count_79_io_out ? io_r_6_b : _GEN_16105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16107 = 8'h7 == r_count_79_io_out ? io_r_7_b : _GEN_16106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16108 = 8'h8 == r_count_79_io_out ? io_r_8_b : _GEN_16107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16109 = 8'h9 == r_count_79_io_out ? io_r_9_b : _GEN_16108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16110 = 8'ha == r_count_79_io_out ? io_r_10_b : _GEN_16109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16111 = 8'hb == r_count_79_io_out ? io_r_11_b : _GEN_16110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16112 = 8'hc == r_count_79_io_out ? io_r_12_b : _GEN_16111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16113 = 8'hd == r_count_79_io_out ? io_r_13_b : _GEN_16112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16114 = 8'he == r_count_79_io_out ? io_r_14_b : _GEN_16113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16115 = 8'hf == r_count_79_io_out ? io_r_15_b : _GEN_16114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16116 = 8'h10 == r_count_79_io_out ? io_r_16_b : _GEN_16115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16117 = 8'h11 == r_count_79_io_out ? io_r_17_b : _GEN_16116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16118 = 8'h12 == r_count_79_io_out ? io_r_18_b : _GEN_16117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16119 = 8'h13 == r_count_79_io_out ? io_r_19_b : _GEN_16118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16120 = 8'h14 == r_count_79_io_out ? io_r_20_b : _GEN_16119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16121 = 8'h15 == r_count_79_io_out ? io_r_21_b : _GEN_16120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16122 = 8'h16 == r_count_79_io_out ? io_r_22_b : _GEN_16121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16123 = 8'h17 == r_count_79_io_out ? io_r_23_b : _GEN_16122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16124 = 8'h18 == r_count_79_io_out ? io_r_24_b : _GEN_16123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16125 = 8'h19 == r_count_79_io_out ? io_r_25_b : _GEN_16124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16126 = 8'h1a == r_count_79_io_out ? io_r_26_b : _GEN_16125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16127 = 8'h1b == r_count_79_io_out ? io_r_27_b : _GEN_16126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16128 = 8'h1c == r_count_79_io_out ? io_r_28_b : _GEN_16127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16129 = 8'h1d == r_count_79_io_out ? io_r_29_b : _GEN_16128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16130 = 8'h1e == r_count_79_io_out ? io_r_30_b : _GEN_16129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16131 = 8'h1f == r_count_79_io_out ? io_r_31_b : _GEN_16130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16132 = 8'h20 == r_count_79_io_out ? io_r_32_b : _GEN_16131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16133 = 8'h21 == r_count_79_io_out ? io_r_33_b : _GEN_16132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16134 = 8'h22 == r_count_79_io_out ? io_r_34_b : _GEN_16133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16135 = 8'h23 == r_count_79_io_out ? io_r_35_b : _GEN_16134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16136 = 8'h24 == r_count_79_io_out ? io_r_36_b : _GEN_16135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16137 = 8'h25 == r_count_79_io_out ? io_r_37_b : _GEN_16136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16138 = 8'h26 == r_count_79_io_out ? io_r_38_b : _GEN_16137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16139 = 8'h27 == r_count_79_io_out ? io_r_39_b : _GEN_16138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16140 = 8'h28 == r_count_79_io_out ? io_r_40_b : _GEN_16139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16141 = 8'h29 == r_count_79_io_out ? io_r_41_b : _GEN_16140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16142 = 8'h2a == r_count_79_io_out ? io_r_42_b : _GEN_16141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16143 = 8'h2b == r_count_79_io_out ? io_r_43_b : _GEN_16142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16144 = 8'h2c == r_count_79_io_out ? io_r_44_b : _GEN_16143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16145 = 8'h2d == r_count_79_io_out ? io_r_45_b : _GEN_16144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16146 = 8'h2e == r_count_79_io_out ? io_r_46_b : _GEN_16145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16147 = 8'h2f == r_count_79_io_out ? io_r_47_b : _GEN_16146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16148 = 8'h30 == r_count_79_io_out ? io_r_48_b : _GEN_16147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16149 = 8'h31 == r_count_79_io_out ? io_r_49_b : _GEN_16148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16150 = 8'h32 == r_count_79_io_out ? io_r_50_b : _GEN_16149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16151 = 8'h33 == r_count_79_io_out ? io_r_51_b : _GEN_16150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16152 = 8'h34 == r_count_79_io_out ? io_r_52_b : _GEN_16151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16153 = 8'h35 == r_count_79_io_out ? io_r_53_b : _GEN_16152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16154 = 8'h36 == r_count_79_io_out ? io_r_54_b : _GEN_16153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16155 = 8'h37 == r_count_79_io_out ? io_r_55_b : _GEN_16154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16156 = 8'h38 == r_count_79_io_out ? io_r_56_b : _GEN_16155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16157 = 8'h39 == r_count_79_io_out ? io_r_57_b : _GEN_16156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16158 = 8'h3a == r_count_79_io_out ? io_r_58_b : _GEN_16157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16159 = 8'h3b == r_count_79_io_out ? io_r_59_b : _GEN_16158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16160 = 8'h3c == r_count_79_io_out ? io_r_60_b : _GEN_16159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16161 = 8'h3d == r_count_79_io_out ? io_r_61_b : _GEN_16160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16162 = 8'h3e == r_count_79_io_out ? io_r_62_b : _GEN_16161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16163 = 8'h3f == r_count_79_io_out ? io_r_63_b : _GEN_16162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16164 = 8'h40 == r_count_79_io_out ? io_r_64_b : _GEN_16163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16165 = 8'h41 == r_count_79_io_out ? io_r_65_b : _GEN_16164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16166 = 8'h42 == r_count_79_io_out ? io_r_66_b : _GEN_16165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16167 = 8'h43 == r_count_79_io_out ? io_r_67_b : _GEN_16166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16168 = 8'h44 == r_count_79_io_out ? io_r_68_b : _GEN_16167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16169 = 8'h45 == r_count_79_io_out ? io_r_69_b : _GEN_16168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16170 = 8'h46 == r_count_79_io_out ? io_r_70_b : _GEN_16169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16171 = 8'h47 == r_count_79_io_out ? io_r_71_b : _GEN_16170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16172 = 8'h48 == r_count_79_io_out ? io_r_72_b : _GEN_16171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16173 = 8'h49 == r_count_79_io_out ? io_r_73_b : _GEN_16172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16174 = 8'h4a == r_count_79_io_out ? io_r_74_b : _GEN_16173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16175 = 8'h4b == r_count_79_io_out ? io_r_75_b : _GEN_16174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16176 = 8'h4c == r_count_79_io_out ? io_r_76_b : _GEN_16175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16177 = 8'h4d == r_count_79_io_out ? io_r_77_b : _GEN_16176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16178 = 8'h4e == r_count_79_io_out ? io_r_78_b : _GEN_16177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16179 = 8'h4f == r_count_79_io_out ? io_r_79_b : _GEN_16178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16180 = 8'h50 == r_count_79_io_out ? io_r_80_b : _GEN_16179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16181 = 8'h51 == r_count_79_io_out ? io_r_81_b : _GEN_16180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16182 = 8'h52 == r_count_79_io_out ? io_r_82_b : _GEN_16181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16183 = 8'h53 == r_count_79_io_out ? io_r_83_b : _GEN_16182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16184 = 8'h54 == r_count_79_io_out ? io_r_84_b : _GEN_16183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16185 = 8'h55 == r_count_79_io_out ? io_r_85_b : _GEN_16184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16186 = 8'h56 == r_count_79_io_out ? io_r_86_b : _GEN_16185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16187 = 8'h57 == r_count_79_io_out ? io_r_87_b : _GEN_16186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16188 = 8'h58 == r_count_79_io_out ? io_r_88_b : _GEN_16187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16189 = 8'h59 == r_count_79_io_out ? io_r_89_b : _GEN_16188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16190 = 8'h5a == r_count_79_io_out ? io_r_90_b : _GEN_16189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16191 = 8'h5b == r_count_79_io_out ? io_r_91_b : _GEN_16190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16192 = 8'h5c == r_count_79_io_out ? io_r_92_b : _GEN_16191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16193 = 8'h5d == r_count_79_io_out ? io_r_93_b : _GEN_16192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16194 = 8'h5e == r_count_79_io_out ? io_r_94_b : _GEN_16193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16195 = 8'h5f == r_count_79_io_out ? io_r_95_b : _GEN_16194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16196 = 8'h60 == r_count_79_io_out ? io_r_96_b : _GEN_16195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16197 = 8'h61 == r_count_79_io_out ? io_r_97_b : _GEN_16196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16198 = 8'h62 == r_count_79_io_out ? io_r_98_b : _GEN_16197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16199 = 8'h63 == r_count_79_io_out ? io_r_99_b : _GEN_16198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16200 = 8'h64 == r_count_79_io_out ? io_r_100_b : _GEN_16199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16201 = 8'h65 == r_count_79_io_out ? io_r_101_b : _GEN_16200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16202 = 8'h66 == r_count_79_io_out ? io_r_102_b : _GEN_16201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16203 = 8'h67 == r_count_79_io_out ? io_r_103_b : _GEN_16202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16204 = 8'h68 == r_count_79_io_out ? io_r_104_b : _GEN_16203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16205 = 8'h69 == r_count_79_io_out ? io_r_105_b : _GEN_16204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16206 = 8'h6a == r_count_79_io_out ? io_r_106_b : _GEN_16205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16207 = 8'h6b == r_count_79_io_out ? io_r_107_b : _GEN_16206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16208 = 8'h6c == r_count_79_io_out ? io_r_108_b : _GEN_16207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16209 = 8'h6d == r_count_79_io_out ? io_r_109_b : _GEN_16208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16210 = 8'h6e == r_count_79_io_out ? io_r_110_b : _GEN_16209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16211 = 8'h6f == r_count_79_io_out ? io_r_111_b : _GEN_16210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16212 = 8'h70 == r_count_79_io_out ? io_r_112_b : _GEN_16211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16213 = 8'h71 == r_count_79_io_out ? io_r_113_b : _GEN_16212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16214 = 8'h72 == r_count_79_io_out ? io_r_114_b : _GEN_16213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16215 = 8'h73 == r_count_79_io_out ? io_r_115_b : _GEN_16214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16216 = 8'h74 == r_count_79_io_out ? io_r_116_b : _GEN_16215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16217 = 8'h75 == r_count_79_io_out ? io_r_117_b : _GEN_16216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16218 = 8'h76 == r_count_79_io_out ? io_r_118_b : _GEN_16217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16219 = 8'h77 == r_count_79_io_out ? io_r_119_b : _GEN_16218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16220 = 8'h78 == r_count_79_io_out ? io_r_120_b : _GEN_16219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16221 = 8'h79 == r_count_79_io_out ? io_r_121_b : _GEN_16220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16222 = 8'h7a == r_count_79_io_out ? io_r_122_b : _GEN_16221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16223 = 8'h7b == r_count_79_io_out ? io_r_123_b : _GEN_16222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16224 = 8'h7c == r_count_79_io_out ? io_r_124_b : _GEN_16223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16225 = 8'h7d == r_count_79_io_out ? io_r_125_b : _GEN_16224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16226 = 8'h7e == r_count_79_io_out ? io_r_126_b : _GEN_16225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16227 = 8'h7f == r_count_79_io_out ? io_r_127_b : _GEN_16226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16228 = 8'h80 == r_count_79_io_out ? io_r_128_b : _GEN_16227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16229 = 8'h81 == r_count_79_io_out ? io_r_129_b : _GEN_16228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16230 = 8'h82 == r_count_79_io_out ? io_r_130_b : _GEN_16229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16231 = 8'h83 == r_count_79_io_out ? io_r_131_b : _GEN_16230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16232 = 8'h84 == r_count_79_io_out ? io_r_132_b : _GEN_16231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16233 = 8'h85 == r_count_79_io_out ? io_r_133_b : _GEN_16232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16234 = 8'h86 == r_count_79_io_out ? io_r_134_b : _GEN_16233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16235 = 8'h87 == r_count_79_io_out ? io_r_135_b : _GEN_16234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16236 = 8'h88 == r_count_79_io_out ? io_r_136_b : _GEN_16235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16237 = 8'h89 == r_count_79_io_out ? io_r_137_b : _GEN_16236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16238 = 8'h8a == r_count_79_io_out ? io_r_138_b : _GEN_16237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16239 = 8'h8b == r_count_79_io_out ? io_r_139_b : _GEN_16238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16240 = 8'h8c == r_count_79_io_out ? io_r_140_b : _GEN_16239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16241 = 8'h8d == r_count_79_io_out ? io_r_141_b : _GEN_16240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16242 = 8'h8e == r_count_79_io_out ? io_r_142_b : _GEN_16241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16243 = 8'h8f == r_count_79_io_out ? io_r_143_b : _GEN_16242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16244 = 8'h90 == r_count_79_io_out ? io_r_144_b : _GEN_16243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16245 = 8'h91 == r_count_79_io_out ? io_r_145_b : _GEN_16244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16246 = 8'h92 == r_count_79_io_out ? io_r_146_b : _GEN_16245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16247 = 8'h93 == r_count_79_io_out ? io_r_147_b : _GEN_16246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16248 = 8'h94 == r_count_79_io_out ? io_r_148_b : _GEN_16247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16249 = 8'h95 == r_count_79_io_out ? io_r_149_b : _GEN_16248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16250 = 8'h96 == r_count_79_io_out ? io_r_150_b : _GEN_16249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16251 = 8'h97 == r_count_79_io_out ? io_r_151_b : _GEN_16250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16252 = 8'h98 == r_count_79_io_out ? io_r_152_b : _GEN_16251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16253 = 8'h99 == r_count_79_io_out ? io_r_153_b : _GEN_16252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16254 = 8'h9a == r_count_79_io_out ? io_r_154_b : _GEN_16253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16255 = 8'h9b == r_count_79_io_out ? io_r_155_b : _GEN_16254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16256 = 8'h9c == r_count_79_io_out ? io_r_156_b : _GEN_16255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16257 = 8'h9d == r_count_79_io_out ? io_r_157_b : _GEN_16256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16258 = 8'h9e == r_count_79_io_out ? io_r_158_b : _GEN_16257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16259 = 8'h9f == r_count_79_io_out ? io_r_159_b : _GEN_16258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16260 = 8'ha0 == r_count_79_io_out ? io_r_160_b : _GEN_16259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16261 = 8'ha1 == r_count_79_io_out ? io_r_161_b : _GEN_16260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16262 = 8'ha2 == r_count_79_io_out ? io_r_162_b : _GEN_16261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16263 = 8'ha3 == r_count_79_io_out ? io_r_163_b : _GEN_16262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16264 = 8'ha4 == r_count_79_io_out ? io_r_164_b : _GEN_16263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16265 = 8'ha5 == r_count_79_io_out ? io_r_165_b : _GEN_16264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16266 = 8'ha6 == r_count_79_io_out ? io_r_166_b : _GEN_16265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16267 = 8'ha7 == r_count_79_io_out ? io_r_167_b : _GEN_16266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16268 = 8'ha8 == r_count_79_io_out ? io_r_168_b : _GEN_16267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16269 = 8'ha9 == r_count_79_io_out ? io_r_169_b : _GEN_16268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16270 = 8'haa == r_count_79_io_out ? io_r_170_b : _GEN_16269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16271 = 8'hab == r_count_79_io_out ? io_r_171_b : _GEN_16270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16272 = 8'hac == r_count_79_io_out ? io_r_172_b : _GEN_16271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16273 = 8'had == r_count_79_io_out ? io_r_173_b : _GEN_16272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16274 = 8'hae == r_count_79_io_out ? io_r_174_b : _GEN_16273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16275 = 8'haf == r_count_79_io_out ? io_r_175_b : _GEN_16274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16276 = 8'hb0 == r_count_79_io_out ? io_r_176_b : _GEN_16275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16277 = 8'hb1 == r_count_79_io_out ? io_r_177_b : _GEN_16276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16278 = 8'hb2 == r_count_79_io_out ? io_r_178_b : _GEN_16277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16279 = 8'hb3 == r_count_79_io_out ? io_r_179_b : _GEN_16278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16280 = 8'hb4 == r_count_79_io_out ? io_r_180_b : _GEN_16279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16281 = 8'hb5 == r_count_79_io_out ? io_r_181_b : _GEN_16280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16282 = 8'hb6 == r_count_79_io_out ? io_r_182_b : _GEN_16281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16283 = 8'hb7 == r_count_79_io_out ? io_r_183_b : _GEN_16282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16284 = 8'hb8 == r_count_79_io_out ? io_r_184_b : _GEN_16283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16285 = 8'hb9 == r_count_79_io_out ? io_r_185_b : _GEN_16284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16286 = 8'hba == r_count_79_io_out ? io_r_186_b : _GEN_16285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16287 = 8'hbb == r_count_79_io_out ? io_r_187_b : _GEN_16286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16288 = 8'hbc == r_count_79_io_out ? io_r_188_b : _GEN_16287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16289 = 8'hbd == r_count_79_io_out ? io_r_189_b : _GEN_16288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16290 = 8'hbe == r_count_79_io_out ? io_r_190_b : _GEN_16289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16291 = 8'hbf == r_count_79_io_out ? io_r_191_b : _GEN_16290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16292 = 8'hc0 == r_count_79_io_out ? io_r_192_b : _GEN_16291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16293 = 8'hc1 == r_count_79_io_out ? io_r_193_b : _GEN_16292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16294 = 8'hc2 == r_count_79_io_out ? io_r_194_b : _GEN_16293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16295 = 8'hc3 == r_count_79_io_out ? io_r_195_b : _GEN_16294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16296 = 8'hc4 == r_count_79_io_out ? io_r_196_b : _GEN_16295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16297 = 8'hc5 == r_count_79_io_out ? io_r_197_b : _GEN_16296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16298 = 8'hc6 == r_count_79_io_out ? io_r_198_b : _GEN_16297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16301 = 8'h1 == r_count_80_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16302 = 8'h2 == r_count_80_io_out ? io_r_2_b : _GEN_16301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16303 = 8'h3 == r_count_80_io_out ? io_r_3_b : _GEN_16302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16304 = 8'h4 == r_count_80_io_out ? io_r_4_b : _GEN_16303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16305 = 8'h5 == r_count_80_io_out ? io_r_5_b : _GEN_16304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16306 = 8'h6 == r_count_80_io_out ? io_r_6_b : _GEN_16305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16307 = 8'h7 == r_count_80_io_out ? io_r_7_b : _GEN_16306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16308 = 8'h8 == r_count_80_io_out ? io_r_8_b : _GEN_16307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16309 = 8'h9 == r_count_80_io_out ? io_r_9_b : _GEN_16308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16310 = 8'ha == r_count_80_io_out ? io_r_10_b : _GEN_16309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16311 = 8'hb == r_count_80_io_out ? io_r_11_b : _GEN_16310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16312 = 8'hc == r_count_80_io_out ? io_r_12_b : _GEN_16311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16313 = 8'hd == r_count_80_io_out ? io_r_13_b : _GEN_16312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16314 = 8'he == r_count_80_io_out ? io_r_14_b : _GEN_16313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16315 = 8'hf == r_count_80_io_out ? io_r_15_b : _GEN_16314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16316 = 8'h10 == r_count_80_io_out ? io_r_16_b : _GEN_16315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16317 = 8'h11 == r_count_80_io_out ? io_r_17_b : _GEN_16316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16318 = 8'h12 == r_count_80_io_out ? io_r_18_b : _GEN_16317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16319 = 8'h13 == r_count_80_io_out ? io_r_19_b : _GEN_16318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16320 = 8'h14 == r_count_80_io_out ? io_r_20_b : _GEN_16319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16321 = 8'h15 == r_count_80_io_out ? io_r_21_b : _GEN_16320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16322 = 8'h16 == r_count_80_io_out ? io_r_22_b : _GEN_16321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16323 = 8'h17 == r_count_80_io_out ? io_r_23_b : _GEN_16322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16324 = 8'h18 == r_count_80_io_out ? io_r_24_b : _GEN_16323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16325 = 8'h19 == r_count_80_io_out ? io_r_25_b : _GEN_16324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16326 = 8'h1a == r_count_80_io_out ? io_r_26_b : _GEN_16325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16327 = 8'h1b == r_count_80_io_out ? io_r_27_b : _GEN_16326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16328 = 8'h1c == r_count_80_io_out ? io_r_28_b : _GEN_16327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16329 = 8'h1d == r_count_80_io_out ? io_r_29_b : _GEN_16328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16330 = 8'h1e == r_count_80_io_out ? io_r_30_b : _GEN_16329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16331 = 8'h1f == r_count_80_io_out ? io_r_31_b : _GEN_16330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16332 = 8'h20 == r_count_80_io_out ? io_r_32_b : _GEN_16331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16333 = 8'h21 == r_count_80_io_out ? io_r_33_b : _GEN_16332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16334 = 8'h22 == r_count_80_io_out ? io_r_34_b : _GEN_16333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16335 = 8'h23 == r_count_80_io_out ? io_r_35_b : _GEN_16334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16336 = 8'h24 == r_count_80_io_out ? io_r_36_b : _GEN_16335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16337 = 8'h25 == r_count_80_io_out ? io_r_37_b : _GEN_16336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16338 = 8'h26 == r_count_80_io_out ? io_r_38_b : _GEN_16337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16339 = 8'h27 == r_count_80_io_out ? io_r_39_b : _GEN_16338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16340 = 8'h28 == r_count_80_io_out ? io_r_40_b : _GEN_16339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16341 = 8'h29 == r_count_80_io_out ? io_r_41_b : _GEN_16340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16342 = 8'h2a == r_count_80_io_out ? io_r_42_b : _GEN_16341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16343 = 8'h2b == r_count_80_io_out ? io_r_43_b : _GEN_16342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16344 = 8'h2c == r_count_80_io_out ? io_r_44_b : _GEN_16343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16345 = 8'h2d == r_count_80_io_out ? io_r_45_b : _GEN_16344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16346 = 8'h2e == r_count_80_io_out ? io_r_46_b : _GEN_16345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16347 = 8'h2f == r_count_80_io_out ? io_r_47_b : _GEN_16346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16348 = 8'h30 == r_count_80_io_out ? io_r_48_b : _GEN_16347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16349 = 8'h31 == r_count_80_io_out ? io_r_49_b : _GEN_16348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16350 = 8'h32 == r_count_80_io_out ? io_r_50_b : _GEN_16349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16351 = 8'h33 == r_count_80_io_out ? io_r_51_b : _GEN_16350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16352 = 8'h34 == r_count_80_io_out ? io_r_52_b : _GEN_16351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16353 = 8'h35 == r_count_80_io_out ? io_r_53_b : _GEN_16352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16354 = 8'h36 == r_count_80_io_out ? io_r_54_b : _GEN_16353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16355 = 8'h37 == r_count_80_io_out ? io_r_55_b : _GEN_16354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16356 = 8'h38 == r_count_80_io_out ? io_r_56_b : _GEN_16355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16357 = 8'h39 == r_count_80_io_out ? io_r_57_b : _GEN_16356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16358 = 8'h3a == r_count_80_io_out ? io_r_58_b : _GEN_16357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16359 = 8'h3b == r_count_80_io_out ? io_r_59_b : _GEN_16358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16360 = 8'h3c == r_count_80_io_out ? io_r_60_b : _GEN_16359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16361 = 8'h3d == r_count_80_io_out ? io_r_61_b : _GEN_16360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16362 = 8'h3e == r_count_80_io_out ? io_r_62_b : _GEN_16361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16363 = 8'h3f == r_count_80_io_out ? io_r_63_b : _GEN_16362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16364 = 8'h40 == r_count_80_io_out ? io_r_64_b : _GEN_16363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16365 = 8'h41 == r_count_80_io_out ? io_r_65_b : _GEN_16364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16366 = 8'h42 == r_count_80_io_out ? io_r_66_b : _GEN_16365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16367 = 8'h43 == r_count_80_io_out ? io_r_67_b : _GEN_16366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16368 = 8'h44 == r_count_80_io_out ? io_r_68_b : _GEN_16367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16369 = 8'h45 == r_count_80_io_out ? io_r_69_b : _GEN_16368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16370 = 8'h46 == r_count_80_io_out ? io_r_70_b : _GEN_16369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16371 = 8'h47 == r_count_80_io_out ? io_r_71_b : _GEN_16370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16372 = 8'h48 == r_count_80_io_out ? io_r_72_b : _GEN_16371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16373 = 8'h49 == r_count_80_io_out ? io_r_73_b : _GEN_16372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16374 = 8'h4a == r_count_80_io_out ? io_r_74_b : _GEN_16373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16375 = 8'h4b == r_count_80_io_out ? io_r_75_b : _GEN_16374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16376 = 8'h4c == r_count_80_io_out ? io_r_76_b : _GEN_16375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16377 = 8'h4d == r_count_80_io_out ? io_r_77_b : _GEN_16376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16378 = 8'h4e == r_count_80_io_out ? io_r_78_b : _GEN_16377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16379 = 8'h4f == r_count_80_io_out ? io_r_79_b : _GEN_16378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16380 = 8'h50 == r_count_80_io_out ? io_r_80_b : _GEN_16379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16381 = 8'h51 == r_count_80_io_out ? io_r_81_b : _GEN_16380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16382 = 8'h52 == r_count_80_io_out ? io_r_82_b : _GEN_16381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16383 = 8'h53 == r_count_80_io_out ? io_r_83_b : _GEN_16382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16384 = 8'h54 == r_count_80_io_out ? io_r_84_b : _GEN_16383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16385 = 8'h55 == r_count_80_io_out ? io_r_85_b : _GEN_16384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16386 = 8'h56 == r_count_80_io_out ? io_r_86_b : _GEN_16385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16387 = 8'h57 == r_count_80_io_out ? io_r_87_b : _GEN_16386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16388 = 8'h58 == r_count_80_io_out ? io_r_88_b : _GEN_16387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16389 = 8'h59 == r_count_80_io_out ? io_r_89_b : _GEN_16388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16390 = 8'h5a == r_count_80_io_out ? io_r_90_b : _GEN_16389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16391 = 8'h5b == r_count_80_io_out ? io_r_91_b : _GEN_16390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16392 = 8'h5c == r_count_80_io_out ? io_r_92_b : _GEN_16391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16393 = 8'h5d == r_count_80_io_out ? io_r_93_b : _GEN_16392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16394 = 8'h5e == r_count_80_io_out ? io_r_94_b : _GEN_16393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16395 = 8'h5f == r_count_80_io_out ? io_r_95_b : _GEN_16394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16396 = 8'h60 == r_count_80_io_out ? io_r_96_b : _GEN_16395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16397 = 8'h61 == r_count_80_io_out ? io_r_97_b : _GEN_16396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16398 = 8'h62 == r_count_80_io_out ? io_r_98_b : _GEN_16397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16399 = 8'h63 == r_count_80_io_out ? io_r_99_b : _GEN_16398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16400 = 8'h64 == r_count_80_io_out ? io_r_100_b : _GEN_16399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16401 = 8'h65 == r_count_80_io_out ? io_r_101_b : _GEN_16400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16402 = 8'h66 == r_count_80_io_out ? io_r_102_b : _GEN_16401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16403 = 8'h67 == r_count_80_io_out ? io_r_103_b : _GEN_16402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16404 = 8'h68 == r_count_80_io_out ? io_r_104_b : _GEN_16403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16405 = 8'h69 == r_count_80_io_out ? io_r_105_b : _GEN_16404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16406 = 8'h6a == r_count_80_io_out ? io_r_106_b : _GEN_16405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16407 = 8'h6b == r_count_80_io_out ? io_r_107_b : _GEN_16406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16408 = 8'h6c == r_count_80_io_out ? io_r_108_b : _GEN_16407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16409 = 8'h6d == r_count_80_io_out ? io_r_109_b : _GEN_16408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16410 = 8'h6e == r_count_80_io_out ? io_r_110_b : _GEN_16409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16411 = 8'h6f == r_count_80_io_out ? io_r_111_b : _GEN_16410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16412 = 8'h70 == r_count_80_io_out ? io_r_112_b : _GEN_16411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16413 = 8'h71 == r_count_80_io_out ? io_r_113_b : _GEN_16412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16414 = 8'h72 == r_count_80_io_out ? io_r_114_b : _GEN_16413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16415 = 8'h73 == r_count_80_io_out ? io_r_115_b : _GEN_16414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16416 = 8'h74 == r_count_80_io_out ? io_r_116_b : _GEN_16415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16417 = 8'h75 == r_count_80_io_out ? io_r_117_b : _GEN_16416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16418 = 8'h76 == r_count_80_io_out ? io_r_118_b : _GEN_16417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16419 = 8'h77 == r_count_80_io_out ? io_r_119_b : _GEN_16418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16420 = 8'h78 == r_count_80_io_out ? io_r_120_b : _GEN_16419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16421 = 8'h79 == r_count_80_io_out ? io_r_121_b : _GEN_16420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16422 = 8'h7a == r_count_80_io_out ? io_r_122_b : _GEN_16421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16423 = 8'h7b == r_count_80_io_out ? io_r_123_b : _GEN_16422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16424 = 8'h7c == r_count_80_io_out ? io_r_124_b : _GEN_16423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16425 = 8'h7d == r_count_80_io_out ? io_r_125_b : _GEN_16424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16426 = 8'h7e == r_count_80_io_out ? io_r_126_b : _GEN_16425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16427 = 8'h7f == r_count_80_io_out ? io_r_127_b : _GEN_16426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16428 = 8'h80 == r_count_80_io_out ? io_r_128_b : _GEN_16427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16429 = 8'h81 == r_count_80_io_out ? io_r_129_b : _GEN_16428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16430 = 8'h82 == r_count_80_io_out ? io_r_130_b : _GEN_16429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16431 = 8'h83 == r_count_80_io_out ? io_r_131_b : _GEN_16430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16432 = 8'h84 == r_count_80_io_out ? io_r_132_b : _GEN_16431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16433 = 8'h85 == r_count_80_io_out ? io_r_133_b : _GEN_16432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16434 = 8'h86 == r_count_80_io_out ? io_r_134_b : _GEN_16433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16435 = 8'h87 == r_count_80_io_out ? io_r_135_b : _GEN_16434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16436 = 8'h88 == r_count_80_io_out ? io_r_136_b : _GEN_16435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16437 = 8'h89 == r_count_80_io_out ? io_r_137_b : _GEN_16436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16438 = 8'h8a == r_count_80_io_out ? io_r_138_b : _GEN_16437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16439 = 8'h8b == r_count_80_io_out ? io_r_139_b : _GEN_16438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16440 = 8'h8c == r_count_80_io_out ? io_r_140_b : _GEN_16439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16441 = 8'h8d == r_count_80_io_out ? io_r_141_b : _GEN_16440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16442 = 8'h8e == r_count_80_io_out ? io_r_142_b : _GEN_16441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16443 = 8'h8f == r_count_80_io_out ? io_r_143_b : _GEN_16442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16444 = 8'h90 == r_count_80_io_out ? io_r_144_b : _GEN_16443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16445 = 8'h91 == r_count_80_io_out ? io_r_145_b : _GEN_16444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16446 = 8'h92 == r_count_80_io_out ? io_r_146_b : _GEN_16445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16447 = 8'h93 == r_count_80_io_out ? io_r_147_b : _GEN_16446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16448 = 8'h94 == r_count_80_io_out ? io_r_148_b : _GEN_16447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16449 = 8'h95 == r_count_80_io_out ? io_r_149_b : _GEN_16448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16450 = 8'h96 == r_count_80_io_out ? io_r_150_b : _GEN_16449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16451 = 8'h97 == r_count_80_io_out ? io_r_151_b : _GEN_16450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16452 = 8'h98 == r_count_80_io_out ? io_r_152_b : _GEN_16451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16453 = 8'h99 == r_count_80_io_out ? io_r_153_b : _GEN_16452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16454 = 8'h9a == r_count_80_io_out ? io_r_154_b : _GEN_16453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16455 = 8'h9b == r_count_80_io_out ? io_r_155_b : _GEN_16454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16456 = 8'h9c == r_count_80_io_out ? io_r_156_b : _GEN_16455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16457 = 8'h9d == r_count_80_io_out ? io_r_157_b : _GEN_16456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16458 = 8'h9e == r_count_80_io_out ? io_r_158_b : _GEN_16457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16459 = 8'h9f == r_count_80_io_out ? io_r_159_b : _GEN_16458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16460 = 8'ha0 == r_count_80_io_out ? io_r_160_b : _GEN_16459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16461 = 8'ha1 == r_count_80_io_out ? io_r_161_b : _GEN_16460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16462 = 8'ha2 == r_count_80_io_out ? io_r_162_b : _GEN_16461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16463 = 8'ha3 == r_count_80_io_out ? io_r_163_b : _GEN_16462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16464 = 8'ha4 == r_count_80_io_out ? io_r_164_b : _GEN_16463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16465 = 8'ha5 == r_count_80_io_out ? io_r_165_b : _GEN_16464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16466 = 8'ha6 == r_count_80_io_out ? io_r_166_b : _GEN_16465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16467 = 8'ha7 == r_count_80_io_out ? io_r_167_b : _GEN_16466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16468 = 8'ha8 == r_count_80_io_out ? io_r_168_b : _GEN_16467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16469 = 8'ha9 == r_count_80_io_out ? io_r_169_b : _GEN_16468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16470 = 8'haa == r_count_80_io_out ? io_r_170_b : _GEN_16469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16471 = 8'hab == r_count_80_io_out ? io_r_171_b : _GEN_16470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16472 = 8'hac == r_count_80_io_out ? io_r_172_b : _GEN_16471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16473 = 8'had == r_count_80_io_out ? io_r_173_b : _GEN_16472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16474 = 8'hae == r_count_80_io_out ? io_r_174_b : _GEN_16473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16475 = 8'haf == r_count_80_io_out ? io_r_175_b : _GEN_16474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16476 = 8'hb0 == r_count_80_io_out ? io_r_176_b : _GEN_16475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16477 = 8'hb1 == r_count_80_io_out ? io_r_177_b : _GEN_16476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16478 = 8'hb2 == r_count_80_io_out ? io_r_178_b : _GEN_16477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16479 = 8'hb3 == r_count_80_io_out ? io_r_179_b : _GEN_16478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16480 = 8'hb4 == r_count_80_io_out ? io_r_180_b : _GEN_16479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16481 = 8'hb5 == r_count_80_io_out ? io_r_181_b : _GEN_16480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16482 = 8'hb6 == r_count_80_io_out ? io_r_182_b : _GEN_16481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16483 = 8'hb7 == r_count_80_io_out ? io_r_183_b : _GEN_16482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16484 = 8'hb8 == r_count_80_io_out ? io_r_184_b : _GEN_16483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16485 = 8'hb9 == r_count_80_io_out ? io_r_185_b : _GEN_16484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16486 = 8'hba == r_count_80_io_out ? io_r_186_b : _GEN_16485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16487 = 8'hbb == r_count_80_io_out ? io_r_187_b : _GEN_16486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16488 = 8'hbc == r_count_80_io_out ? io_r_188_b : _GEN_16487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16489 = 8'hbd == r_count_80_io_out ? io_r_189_b : _GEN_16488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16490 = 8'hbe == r_count_80_io_out ? io_r_190_b : _GEN_16489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16491 = 8'hbf == r_count_80_io_out ? io_r_191_b : _GEN_16490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16492 = 8'hc0 == r_count_80_io_out ? io_r_192_b : _GEN_16491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16493 = 8'hc1 == r_count_80_io_out ? io_r_193_b : _GEN_16492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16494 = 8'hc2 == r_count_80_io_out ? io_r_194_b : _GEN_16493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16495 = 8'hc3 == r_count_80_io_out ? io_r_195_b : _GEN_16494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16496 = 8'hc4 == r_count_80_io_out ? io_r_196_b : _GEN_16495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16497 = 8'hc5 == r_count_80_io_out ? io_r_197_b : _GEN_16496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16498 = 8'hc6 == r_count_80_io_out ? io_r_198_b : _GEN_16497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16501 = 8'h1 == r_count_81_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16502 = 8'h2 == r_count_81_io_out ? io_r_2_b : _GEN_16501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16503 = 8'h3 == r_count_81_io_out ? io_r_3_b : _GEN_16502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16504 = 8'h4 == r_count_81_io_out ? io_r_4_b : _GEN_16503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16505 = 8'h5 == r_count_81_io_out ? io_r_5_b : _GEN_16504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16506 = 8'h6 == r_count_81_io_out ? io_r_6_b : _GEN_16505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16507 = 8'h7 == r_count_81_io_out ? io_r_7_b : _GEN_16506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16508 = 8'h8 == r_count_81_io_out ? io_r_8_b : _GEN_16507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16509 = 8'h9 == r_count_81_io_out ? io_r_9_b : _GEN_16508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16510 = 8'ha == r_count_81_io_out ? io_r_10_b : _GEN_16509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16511 = 8'hb == r_count_81_io_out ? io_r_11_b : _GEN_16510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16512 = 8'hc == r_count_81_io_out ? io_r_12_b : _GEN_16511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16513 = 8'hd == r_count_81_io_out ? io_r_13_b : _GEN_16512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16514 = 8'he == r_count_81_io_out ? io_r_14_b : _GEN_16513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16515 = 8'hf == r_count_81_io_out ? io_r_15_b : _GEN_16514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16516 = 8'h10 == r_count_81_io_out ? io_r_16_b : _GEN_16515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16517 = 8'h11 == r_count_81_io_out ? io_r_17_b : _GEN_16516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16518 = 8'h12 == r_count_81_io_out ? io_r_18_b : _GEN_16517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16519 = 8'h13 == r_count_81_io_out ? io_r_19_b : _GEN_16518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16520 = 8'h14 == r_count_81_io_out ? io_r_20_b : _GEN_16519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16521 = 8'h15 == r_count_81_io_out ? io_r_21_b : _GEN_16520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16522 = 8'h16 == r_count_81_io_out ? io_r_22_b : _GEN_16521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16523 = 8'h17 == r_count_81_io_out ? io_r_23_b : _GEN_16522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16524 = 8'h18 == r_count_81_io_out ? io_r_24_b : _GEN_16523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16525 = 8'h19 == r_count_81_io_out ? io_r_25_b : _GEN_16524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16526 = 8'h1a == r_count_81_io_out ? io_r_26_b : _GEN_16525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16527 = 8'h1b == r_count_81_io_out ? io_r_27_b : _GEN_16526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16528 = 8'h1c == r_count_81_io_out ? io_r_28_b : _GEN_16527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16529 = 8'h1d == r_count_81_io_out ? io_r_29_b : _GEN_16528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16530 = 8'h1e == r_count_81_io_out ? io_r_30_b : _GEN_16529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16531 = 8'h1f == r_count_81_io_out ? io_r_31_b : _GEN_16530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16532 = 8'h20 == r_count_81_io_out ? io_r_32_b : _GEN_16531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16533 = 8'h21 == r_count_81_io_out ? io_r_33_b : _GEN_16532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16534 = 8'h22 == r_count_81_io_out ? io_r_34_b : _GEN_16533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16535 = 8'h23 == r_count_81_io_out ? io_r_35_b : _GEN_16534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16536 = 8'h24 == r_count_81_io_out ? io_r_36_b : _GEN_16535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16537 = 8'h25 == r_count_81_io_out ? io_r_37_b : _GEN_16536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16538 = 8'h26 == r_count_81_io_out ? io_r_38_b : _GEN_16537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16539 = 8'h27 == r_count_81_io_out ? io_r_39_b : _GEN_16538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16540 = 8'h28 == r_count_81_io_out ? io_r_40_b : _GEN_16539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16541 = 8'h29 == r_count_81_io_out ? io_r_41_b : _GEN_16540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16542 = 8'h2a == r_count_81_io_out ? io_r_42_b : _GEN_16541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16543 = 8'h2b == r_count_81_io_out ? io_r_43_b : _GEN_16542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16544 = 8'h2c == r_count_81_io_out ? io_r_44_b : _GEN_16543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16545 = 8'h2d == r_count_81_io_out ? io_r_45_b : _GEN_16544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16546 = 8'h2e == r_count_81_io_out ? io_r_46_b : _GEN_16545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16547 = 8'h2f == r_count_81_io_out ? io_r_47_b : _GEN_16546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16548 = 8'h30 == r_count_81_io_out ? io_r_48_b : _GEN_16547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16549 = 8'h31 == r_count_81_io_out ? io_r_49_b : _GEN_16548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16550 = 8'h32 == r_count_81_io_out ? io_r_50_b : _GEN_16549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16551 = 8'h33 == r_count_81_io_out ? io_r_51_b : _GEN_16550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16552 = 8'h34 == r_count_81_io_out ? io_r_52_b : _GEN_16551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16553 = 8'h35 == r_count_81_io_out ? io_r_53_b : _GEN_16552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16554 = 8'h36 == r_count_81_io_out ? io_r_54_b : _GEN_16553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16555 = 8'h37 == r_count_81_io_out ? io_r_55_b : _GEN_16554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16556 = 8'h38 == r_count_81_io_out ? io_r_56_b : _GEN_16555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16557 = 8'h39 == r_count_81_io_out ? io_r_57_b : _GEN_16556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16558 = 8'h3a == r_count_81_io_out ? io_r_58_b : _GEN_16557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16559 = 8'h3b == r_count_81_io_out ? io_r_59_b : _GEN_16558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16560 = 8'h3c == r_count_81_io_out ? io_r_60_b : _GEN_16559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16561 = 8'h3d == r_count_81_io_out ? io_r_61_b : _GEN_16560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16562 = 8'h3e == r_count_81_io_out ? io_r_62_b : _GEN_16561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16563 = 8'h3f == r_count_81_io_out ? io_r_63_b : _GEN_16562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16564 = 8'h40 == r_count_81_io_out ? io_r_64_b : _GEN_16563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16565 = 8'h41 == r_count_81_io_out ? io_r_65_b : _GEN_16564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16566 = 8'h42 == r_count_81_io_out ? io_r_66_b : _GEN_16565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16567 = 8'h43 == r_count_81_io_out ? io_r_67_b : _GEN_16566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16568 = 8'h44 == r_count_81_io_out ? io_r_68_b : _GEN_16567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16569 = 8'h45 == r_count_81_io_out ? io_r_69_b : _GEN_16568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16570 = 8'h46 == r_count_81_io_out ? io_r_70_b : _GEN_16569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16571 = 8'h47 == r_count_81_io_out ? io_r_71_b : _GEN_16570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16572 = 8'h48 == r_count_81_io_out ? io_r_72_b : _GEN_16571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16573 = 8'h49 == r_count_81_io_out ? io_r_73_b : _GEN_16572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16574 = 8'h4a == r_count_81_io_out ? io_r_74_b : _GEN_16573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16575 = 8'h4b == r_count_81_io_out ? io_r_75_b : _GEN_16574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16576 = 8'h4c == r_count_81_io_out ? io_r_76_b : _GEN_16575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16577 = 8'h4d == r_count_81_io_out ? io_r_77_b : _GEN_16576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16578 = 8'h4e == r_count_81_io_out ? io_r_78_b : _GEN_16577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16579 = 8'h4f == r_count_81_io_out ? io_r_79_b : _GEN_16578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16580 = 8'h50 == r_count_81_io_out ? io_r_80_b : _GEN_16579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16581 = 8'h51 == r_count_81_io_out ? io_r_81_b : _GEN_16580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16582 = 8'h52 == r_count_81_io_out ? io_r_82_b : _GEN_16581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16583 = 8'h53 == r_count_81_io_out ? io_r_83_b : _GEN_16582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16584 = 8'h54 == r_count_81_io_out ? io_r_84_b : _GEN_16583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16585 = 8'h55 == r_count_81_io_out ? io_r_85_b : _GEN_16584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16586 = 8'h56 == r_count_81_io_out ? io_r_86_b : _GEN_16585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16587 = 8'h57 == r_count_81_io_out ? io_r_87_b : _GEN_16586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16588 = 8'h58 == r_count_81_io_out ? io_r_88_b : _GEN_16587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16589 = 8'h59 == r_count_81_io_out ? io_r_89_b : _GEN_16588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16590 = 8'h5a == r_count_81_io_out ? io_r_90_b : _GEN_16589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16591 = 8'h5b == r_count_81_io_out ? io_r_91_b : _GEN_16590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16592 = 8'h5c == r_count_81_io_out ? io_r_92_b : _GEN_16591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16593 = 8'h5d == r_count_81_io_out ? io_r_93_b : _GEN_16592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16594 = 8'h5e == r_count_81_io_out ? io_r_94_b : _GEN_16593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16595 = 8'h5f == r_count_81_io_out ? io_r_95_b : _GEN_16594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16596 = 8'h60 == r_count_81_io_out ? io_r_96_b : _GEN_16595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16597 = 8'h61 == r_count_81_io_out ? io_r_97_b : _GEN_16596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16598 = 8'h62 == r_count_81_io_out ? io_r_98_b : _GEN_16597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16599 = 8'h63 == r_count_81_io_out ? io_r_99_b : _GEN_16598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16600 = 8'h64 == r_count_81_io_out ? io_r_100_b : _GEN_16599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16601 = 8'h65 == r_count_81_io_out ? io_r_101_b : _GEN_16600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16602 = 8'h66 == r_count_81_io_out ? io_r_102_b : _GEN_16601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16603 = 8'h67 == r_count_81_io_out ? io_r_103_b : _GEN_16602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16604 = 8'h68 == r_count_81_io_out ? io_r_104_b : _GEN_16603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16605 = 8'h69 == r_count_81_io_out ? io_r_105_b : _GEN_16604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16606 = 8'h6a == r_count_81_io_out ? io_r_106_b : _GEN_16605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16607 = 8'h6b == r_count_81_io_out ? io_r_107_b : _GEN_16606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16608 = 8'h6c == r_count_81_io_out ? io_r_108_b : _GEN_16607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16609 = 8'h6d == r_count_81_io_out ? io_r_109_b : _GEN_16608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16610 = 8'h6e == r_count_81_io_out ? io_r_110_b : _GEN_16609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16611 = 8'h6f == r_count_81_io_out ? io_r_111_b : _GEN_16610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16612 = 8'h70 == r_count_81_io_out ? io_r_112_b : _GEN_16611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16613 = 8'h71 == r_count_81_io_out ? io_r_113_b : _GEN_16612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16614 = 8'h72 == r_count_81_io_out ? io_r_114_b : _GEN_16613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16615 = 8'h73 == r_count_81_io_out ? io_r_115_b : _GEN_16614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16616 = 8'h74 == r_count_81_io_out ? io_r_116_b : _GEN_16615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16617 = 8'h75 == r_count_81_io_out ? io_r_117_b : _GEN_16616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16618 = 8'h76 == r_count_81_io_out ? io_r_118_b : _GEN_16617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16619 = 8'h77 == r_count_81_io_out ? io_r_119_b : _GEN_16618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16620 = 8'h78 == r_count_81_io_out ? io_r_120_b : _GEN_16619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16621 = 8'h79 == r_count_81_io_out ? io_r_121_b : _GEN_16620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16622 = 8'h7a == r_count_81_io_out ? io_r_122_b : _GEN_16621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16623 = 8'h7b == r_count_81_io_out ? io_r_123_b : _GEN_16622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16624 = 8'h7c == r_count_81_io_out ? io_r_124_b : _GEN_16623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16625 = 8'h7d == r_count_81_io_out ? io_r_125_b : _GEN_16624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16626 = 8'h7e == r_count_81_io_out ? io_r_126_b : _GEN_16625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16627 = 8'h7f == r_count_81_io_out ? io_r_127_b : _GEN_16626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16628 = 8'h80 == r_count_81_io_out ? io_r_128_b : _GEN_16627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16629 = 8'h81 == r_count_81_io_out ? io_r_129_b : _GEN_16628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16630 = 8'h82 == r_count_81_io_out ? io_r_130_b : _GEN_16629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16631 = 8'h83 == r_count_81_io_out ? io_r_131_b : _GEN_16630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16632 = 8'h84 == r_count_81_io_out ? io_r_132_b : _GEN_16631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16633 = 8'h85 == r_count_81_io_out ? io_r_133_b : _GEN_16632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16634 = 8'h86 == r_count_81_io_out ? io_r_134_b : _GEN_16633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16635 = 8'h87 == r_count_81_io_out ? io_r_135_b : _GEN_16634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16636 = 8'h88 == r_count_81_io_out ? io_r_136_b : _GEN_16635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16637 = 8'h89 == r_count_81_io_out ? io_r_137_b : _GEN_16636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16638 = 8'h8a == r_count_81_io_out ? io_r_138_b : _GEN_16637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16639 = 8'h8b == r_count_81_io_out ? io_r_139_b : _GEN_16638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16640 = 8'h8c == r_count_81_io_out ? io_r_140_b : _GEN_16639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16641 = 8'h8d == r_count_81_io_out ? io_r_141_b : _GEN_16640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16642 = 8'h8e == r_count_81_io_out ? io_r_142_b : _GEN_16641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16643 = 8'h8f == r_count_81_io_out ? io_r_143_b : _GEN_16642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16644 = 8'h90 == r_count_81_io_out ? io_r_144_b : _GEN_16643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16645 = 8'h91 == r_count_81_io_out ? io_r_145_b : _GEN_16644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16646 = 8'h92 == r_count_81_io_out ? io_r_146_b : _GEN_16645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16647 = 8'h93 == r_count_81_io_out ? io_r_147_b : _GEN_16646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16648 = 8'h94 == r_count_81_io_out ? io_r_148_b : _GEN_16647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16649 = 8'h95 == r_count_81_io_out ? io_r_149_b : _GEN_16648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16650 = 8'h96 == r_count_81_io_out ? io_r_150_b : _GEN_16649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16651 = 8'h97 == r_count_81_io_out ? io_r_151_b : _GEN_16650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16652 = 8'h98 == r_count_81_io_out ? io_r_152_b : _GEN_16651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16653 = 8'h99 == r_count_81_io_out ? io_r_153_b : _GEN_16652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16654 = 8'h9a == r_count_81_io_out ? io_r_154_b : _GEN_16653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16655 = 8'h9b == r_count_81_io_out ? io_r_155_b : _GEN_16654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16656 = 8'h9c == r_count_81_io_out ? io_r_156_b : _GEN_16655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16657 = 8'h9d == r_count_81_io_out ? io_r_157_b : _GEN_16656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16658 = 8'h9e == r_count_81_io_out ? io_r_158_b : _GEN_16657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16659 = 8'h9f == r_count_81_io_out ? io_r_159_b : _GEN_16658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16660 = 8'ha0 == r_count_81_io_out ? io_r_160_b : _GEN_16659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16661 = 8'ha1 == r_count_81_io_out ? io_r_161_b : _GEN_16660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16662 = 8'ha2 == r_count_81_io_out ? io_r_162_b : _GEN_16661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16663 = 8'ha3 == r_count_81_io_out ? io_r_163_b : _GEN_16662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16664 = 8'ha4 == r_count_81_io_out ? io_r_164_b : _GEN_16663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16665 = 8'ha5 == r_count_81_io_out ? io_r_165_b : _GEN_16664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16666 = 8'ha6 == r_count_81_io_out ? io_r_166_b : _GEN_16665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16667 = 8'ha7 == r_count_81_io_out ? io_r_167_b : _GEN_16666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16668 = 8'ha8 == r_count_81_io_out ? io_r_168_b : _GEN_16667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16669 = 8'ha9 == r_count_81_io_out ? io_r_169_b : _GEN_16668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16670 = 8'haa == r_count_81_io_out ? io_r_170_b : _GEN_16669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16671 = 8'hab == r_count_81_io_out ? io_r_171_b : _GEN_16670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16672 = 8'hac == r_count_81_io_out ? io_r_172_b : _GEN_16671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16673 = 8'had == r_count_81_io_out ? io_r_173_b : _GEN_16672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16674 = 8'hae == r_count_81_io_out ? io_r_174_b : _GEN_16673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16675 = 8'haf == r_count_81_io_out ? io_r_175_b : _GEN_16674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16676 = 8'hb0 == r_count_81_io_out ? io_r_176_b : _GEN_16675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16677 = 8'hb1 == r_count_81_io_out ? io_r_177_b : _GEN_16676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16678 = 8'hb2 == r_count_81_io_out ? io_r_178_b : _GEN_16677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16679 = 8'hb3 == r_count_81_io_out ? io_r_179_b : _GEN_16678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16680 = 8'hb4 == r_count_81_io_out ? io_r_180_b : _GEN_16679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16681 = 8'hb5 == r_count_81_io_out ? io_r_181_b : _GEN_16680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16682 = 8'hb6 == r_count_81_io_out ? io_r_182_b : _GEN_16681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16683 = 8'hb7 == r_count_81_io_out ? io_r_183_b : _GEN_16682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16684 = 8'hb8 == r_count_81_io_out ? io_r_184_b : _GEN_16683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16685 = 8'hb9 == r_count_81_io_out ? io_r_185_b : _GEN_16684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16686 = 8'hba == r_count_81_io_out ? io_r_186_b : _GEN_16685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16687 = 8'hbb == r_count_81_io_out ? io_r_187_b : _GEN_16686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16688 = 8'hbc == r_count_81_io_out ? io_r_188_b : _GEN_16687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16689 = 8'hbd == r_count_81_io_out ? io_r_189_b : _GEN_16688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16690 = 8'hbe == r_count_81_io_out ? io_r_190_b : _GEN_16689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16691 = 8'hbf == r_count_81_io_out ? io_r_191_b : _GEN_16690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16692 = 8'hc0 == r_count_81_io_out ? io_r_192_b : _GEN_16691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16693 = 8'hc1 == r_count_81_io_out ? io_r_193_b : _GEN_16692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16694 = 8'hc2 == r_count_81_io_out ? io_r_194_b : _GEN_16693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16695 = 8'hc3 == r_count_81_io_out ? io_r_195_b : _GEN_16694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16696 = 8'hc4 == r_count_81_io_out ? io_r_196_b : _GEN_16695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16697 = 8'hc5 == r_count_81_io_out ? io_r_197_b : _GEN_16696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16698 = 8'hc6 == r_count_81_io_out ? io_r_198_b : _GEN_16697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16701 = 8'h1 == r_count_82_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16702 = 8'h2 == r_count_82_io_out ? io_r_2_b : _GEN_16701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16703 = 8'h3 == r_count_82_io_out ? io_r_3_b : _GEN_16702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16704 = 8'h4 == r_count_82_io_out ? io_r_4_b : _GEN_16703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16705 = 8'h5 == r_count_82_io_out ? io_r_5_b : _GEN_16704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16706 = 8'h6 == r_count_82_io_out ? io_r_6_b : _GEN_16705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16707 = 8'h7 == r_count_82_io_out ? io_r_7_b : _GEN_16706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16708 = 8'h8 == r_count_82_io_out ? io_r_8_b : _GEN_16707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16709 = 8'h9 == r_count_82_io_out ? io_r_9_b : _GEN_16708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16710 = 8'ha == r_count_82_io_out ? io_r_10_b : _GEN_16709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16711 = 8'hb == r_count_82_io_out ? io_r_11_b : _GEN_16710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16712 = 8'hc == r_count_82_io_out ? io_r_12_b : _GEN_16711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16713 = 8'hd == r_count_82_io_out ? io_r_13_b : _GEN_16712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16714 = 8'he == r_count_82_io_out ? io_r_14_b : _GEN_16713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16715 = 8'hf == r_count_82_io_out ? io_r_15_b : _GEN_16714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16716 = 8'h10 == r_count_82_io_out ? io_r_16_b : _GEN_16715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16717 = 8'h11 == r_count_82_io_out ? io_r_17_b : _GEN_16716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16718 = 8'h12 == r_count_82_io_out ? io_r_18_b : _GEN_16717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16719 = 8'h13 == r_count_82_io_out ? io_r_19_b : _GEN_16718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16720 = 8'h14 == r_count_82_io_out ? io_r_20_b : _GEN_16719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16721 = 8'h15 == r_count_82_io_out ? io_r_21_b : _GEN_16720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16722 = 8'h16 == r_count_82_io_out ? io_r_22_b : _GEN_16721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16723 = 8'h17 == r_count_82_io_out ? io_r_23_b : _GEN_16722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16724 = 8'h18 == r_count_82_io_out ? io_r_24_b : _GEN_16723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16725 = 8'h19 == r_count_82_io_out ? io_r_25_b : _GEN_16724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16726 = 8'h1a == r_count_82_io_out ? io_r_26_b : _GEN_16725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16727 = 8'h1b == r_count_82_io_out ? io_r_27_b : _GEN_16726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16728 = 8'h1c == r_count_82_io_out ? io_r_28_b : _GEN_16727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16729 = 8'h1d == r_count_82_io_out ? io_r_29_b : _GEN_16728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16730 = 8'h1e == r_count_82_io_out ? io_r_30_b : _GEN_16729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16731 = 8'h1f == r_count_82_io_out ? io_r_31_b : _GEN_16730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16732 = 8'h20 == r_count_82_io_out ? io_r_32_b : _GEN_16731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16733 = 8'h21 == r_count_82_io_out ? io_r_33_b : _GEN_16732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16734 = 8'h22 == r_count_82_io_out ? io_r_34_b : _GEN_16733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16735 = 8'h23 == r_count_82_io_out ? io_r_35_b : _GEN_16734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16736 = 8'h24 == r_count_82_io_out ? io_r_36_b : _GEN_16735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16737 = 8'h25 == r_count_82_io_out ? io_r_37_b : _GEN_16736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16738 = 8'h26 == r_count_82_io_out ? io_r_38_b : _GEN_16737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16739 = 8'h27 == r_count_82_io_out ? io_r_39_b : _GEN_16738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16740 = 8'h28 == r_count_82_io_out ? io_r_40_b : _GEN_16739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16741 = 8'h29 == r_count_82_io_out ? io_r_41_b : _GEN_16740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16742 = 8'h2a == r_count_82_io_out ? io_r_42_b : _GEN_16741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16743 = 8'h2b == r_count_82_io_out ? io_r_43_b : _GEN_16742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16744 = 8'h2c == r_count_82_io_out ? io_r_44_b : _GEN_16743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16745 = 8'h2d == r_count_82_io_out ? io_r_45_b : _GEN_16744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16746 = 8'h2e == r_count_82_io_out ? io_r_46_b : _GEN_16745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16747 = 8'h2f == r_count_82_io_out ? io_r_47_b : _GEN_16746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16748 = 8'h30 == r_count_82_io_out ? io_r_48_b : _GEN_16747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16749 = 8'h31 == r_count_82_io_out ? io_r_49_b : _GEN_16748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16750 = 8'h32 == r_count_82_io_out ? io_r_50_b : _GEN_16749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16751 = 8'h33 == r_count_82_io_out ? io_r_51_b : _GEN_16750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16752 = 8'h34 == r_count_82_io_out ? io_r_52_b : _GEN_16751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16753 = 8'h35 == r_count_82_io_out ? io_r_53_b : _GEN_16752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16754 = 8'h36 == r_count_82_io_out ? io_r_54_b : _GEN_16753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16755 = 8'h37 == r_count_82_io_out ? io_r_55_b : _GEN_16754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16756 = 8'h38 == r_count_82_io_out ? io_r_56_b : _GEN_16755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16757 = 8'h39 == r_count_82_io_out ? io_r_57_b : _GEN_16756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16758 = 8'h3a == r_count_82_io_out ? io_r_58_b : _GEN_16757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16759 = 8'h3b == r_count_82_io_out ? io_r_59_b : _GEN_16758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16760 = 8'h3c == r_count_82_io_out ? io_r_60_b : _GEN_16759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16761 = 8'h3d == r_count_82_io_out ? io_r_61_b : _GEN_16760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16762 = 8'h3e == r_count_82_io_out ? io_r_62_b : _GEN_16761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16763 = 8'h3f == r_count_82_io_out ? io_r_63_b : _GEN_16762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16764 = 8'h40 == r_count_82_io_out ? io_r_64_b : _GEN_16763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16765 = 8'h41 == r_count_82_io_out ? io_r_65_b : _GEN_16764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16766 = 8'h42 == r_count_82_io_out ? io_r_66_b : _GEN_16765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16767 = 8'h43 == r_count_82_io_out ? io_r_67_b : _GEN_16766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16768 = 8'h44 == r_count_82_io_out ? io_r_68_b : _GEN_16767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16769 = 8'h45 == r_count_82_io_out ? io_r_69_b : _GEN_16768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16770 = 8'h46 == r_count_82_io_out ? io_r_70_b : _GEN_16769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16771 = 8'h47 == r_count_82_io_out ? io_r_71_b : _GEN_16770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16772 = 8'h48 == r_count_82_io_out ? io_r_72_b : _GEN_16771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16773 = 8'h49 == r_count_82_io_out ? io_r_73_b : _GEN_16772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16774 = 8'h4a == r_count_82_io_out ? io_r_74_b : _GEN_16773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16775 = 8'h4b == r_count_82_io_out ? io_r_75_b : _GEN_16774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16776 = 8'h4c == r_count_82_io_out ? io_r_76_b : _GEN_16775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16777 = 8'h4d == r_count_82_io_out ? io_r_77_b : _GEN_16776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16778 = 8'h4e == r_count_82_io_out ? io_r_78_b : _GEN_16777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16779 = 8'h4f == r_count_82_io_out ? io_r_79_b : _GEN_16778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16780 = 8'h50 == r_count_82_io_out ? io_r_80_b : _GEN_16779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16781 = 8'h51 == r_count_82_io_out ? io_r_81_b : _GEN_16780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16782 = 8'h52 == r_count_82_io_out ? io_r_82_b : _GEN_16781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16783 = 8'h53 == r_count_82_io_out ? io_r_83_b : _GEN_16782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16784 = 8'h54 == r_count_82_io_out ? io_r_84_b : _GEN_16783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16785 = 8'h55 == r_count_82_io_out ? io_r_85_b : _GEN_16784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16786 = 8'h56 == r_count_82_io_out ? io_r_86_b : _GEN_16785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16787 = 8'h57 == r_count_82_io_out ? io_r_87_b : _GEN_16786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16788 = 8'h58 == r_count_82_io_out ? io_r_88_b : _GEN_16787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16789 = 8'h59 == r_count_82_io_out ? io_r_89_b : _GEN_16788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16790 = 8'h5a == r_count_82_io_out ? io_r_90_b : _GEN_16789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16791 = 8'h5b == r_count_82_io_out ? io_r_91_b : _GEN_16790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16792 = 8'h5c == r_count_82_io_out ? io_r_92_b : _GEN_16791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16793 = 8'h5d == r_count_82_io_out ? io_r_93_b : _GEN_16792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16794 = 8'h5e == r_count_82_io_out ? io_r_94_b : _GEN_16793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16795 = 8'h5f == r_count_82_io_out ? io_r_95_b : _GEN_16794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16796 = 8'h60 == r_count_82_io_out ? io_r_96_b : _GEN_16795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16797 = 8'h61 == r_count_82_io_out ? io_r_97_b : _GEN_16796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16798 = 8'h62 == r_count_82_io_out ? io_r_98_b : _GEN_16797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16799 = 8'h63 == r_count_82_io_out ? io_r_99_b : _GEN_16798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16800 = 8'h64 == r_count_82_io_out ? io_r_100_b : _GEN_16799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16801 = 8'h65 == r_count_82_io_out ? io_r_101_b : _GEN_16800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16802 = 8'h66 == r_count_82_io_out ? io_r_102_b : _GEN_16801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16803 = 8'h67 == r_count_82_io_out ? io_r_103_b : _GEN_16802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16804 = 8'h68 == r_count_82_io_out ? io_r_104_b : _GEN_16803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16805 = 8'h69 == r_count_82_io_out ? io_r_105_b : _GEN_16804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16806 = 8'h6a == r_count_82_io_out ? io_r_106_b : _GEN_16805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16807 = 8'h6b == r_count_82_io_out ? io_r_107_b : _GEN_16806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16808 = 8'h6c == r_count_82_io_out ? io_r_108_b : _GEN_16807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16809 = 8'h6d == r_count_82_io_out ? io_r_109_b : _GEN_16808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16810 = 8'h6e == r_count_82_io_out ? io_r_110_b : _GEN_16809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16811 = 8'h6f == r_count_82_io_out ? io_r_111_b : _GEN_16810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16812 = 8'h70 == r_count_82_io_out ? io_r_112_b : _GEN_16811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16813 = 8'h71 == r_count_82_io_out ? io_r_113_b : _GEN_16812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16814 = 8'h72 == r_count_82_io_out ? io_r_114_b : _GEN_16813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16815 = 8'h73 == r_count_82_io_out ? io_r_115_b : _GEN_16814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16816 = 8'h74 == r_count_82_io_out ? io_r_116_b : _GEN_16815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16817 = 8'h75 == r_count_82_io_out ? io_r_117_b : _GEN_16816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16818 = 8'h76 == r_count_82_io_out ? io_r_118_b : _GEN_16817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16819 = 8'h77 == r_count_82_io_out ? io_r_119_b : _GEN_16818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16820 = 8'h78 == r_count_82_io_out ? io_r_120_b : _GEN_16819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16821 = 8'h79 == r_count_82_io_out ? io_r_121_b : _GEN_16820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16822 = 8'h7a == r_count_82_io_out ? io_r_122_b : _GEN_16821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16823 = 8'h7b == r_count_82_io_out ? io_r_123_b : _GEN_16822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16824 = 8'h7c == r_count_82_io_out ? io_r_124_b : _GEN_16823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16825 = 8'h7d == r_count_82_io_out ? io_r_125_b : _GEN_16824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16826 = 8'h7e == r_count_82_io_out ? io_r_126_b : _GEN_16825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16827 = 8'h7f == r_count_82_io_out ? io_r_127_b : _GEN_16826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16828 = 8'h80 == r_count_82_io_out ? io_r_128_b : _GEN_16827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16829 = 8'h81 == r_count_82_io_out ? io_r_129_b : _GEN_16828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16830 = 8'h82 == r_count_82_io_out ? io_r_130_b : _GEN_16829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16831 = 8'h83 == r_count_82_io_out ? io_r_131_b : _GEN_16830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16832 = 8'h84 == r_count_82_io_out ? io_r_132_b : _GEN_16831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16833 = 8'h85 == r_count_82_io_out ? io_r_133_b : _GEN_16832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16834 = 8'h86 == r_count_82_io_out ? io_r_134_b : _GEN_16833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16835 = 8'h87 == r_count_82_io_out ? io_r_135_b : _GEN_16834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16836 = 8'h88 == r_count_82_io_out ? io_r_136_b : _GEN_16835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16837 = 8'h89 == r_count_82_io_out ? io_r_137_b : _GEN_16836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16838 = 8'h8a == r_count_82_io_out ? io_r_138_b : _GEN_16837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16839 = 8'h8b == r_count_82_io_out ? io_r_139_b : _GEN_16838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16840 = 8'h8c == r_count_82_io_out ? io_r_140_b : _GEN_16839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16841 = 8'h8d == r_count_82_io_out ? io_r_141_b : _GEN_16840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16842 = 8'h8e == r_count_82_io_out ? io_r_142_b : _GEN_16841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16843 = 8'h8f == r_count_82_io_out ? io_r_143_b : _GEN_16842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16844 = 8'h90 == r_count_82_io_out ? io_r_144_b : _GEN_16843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16845 = 8'h91 == r_count_82_io_out ? io_r_145_b : _GEN_16844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16846 = 8'h92 == r_count_82_io_out ? io_r_146_b : _GEN_16845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16847 = 8'h93 == r_count_82_io_out ? io_r_147_b : _GEN_16846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16848 = 8'h94 == r_count_82_io_out ? io_r_148_b : _GEN_16847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16849 = 8'h95 == r_count_82_io_out ? io_r_149_b : _GEN_16848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16850 = 8'h96 == r_count_82_io_out ? io_r_150_b : _GEN_16849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16851 = 8'h97 == r_count_82_io_out ? io_r_151_b : _GEN_16850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16852 = 8'h98 == r_count_82_io_out ? io_r_152_b : _GEN_16851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16853 = 8'h99 == r_count_82_io_out ? io_r_153_b : _GEN_16852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16854 = 8'h9a == r_count_82_io_out ? io_r_154_b : _GEN_16853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16855 = 8'h9b == r_count_82_io_out ? io_r_155_b : _GEN_16854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16856 = 8'h9c == r_count_82_io_out ? io_r_156_b : _GEN_16855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16857 = 8'h9d == r_count_82_io_out ? io_r_157_b : _GEN_16856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16858 = 8'h9e == r_count_82_io_out ? io_r_158_b : _GEN_16857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16859 = 8'h9f == r_count_82_io_out ? io_r_159_b : _GEN_16858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16860 = 8'ha0 == r_count_82_io_out ? io_r_160_b : _GEN_16859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16861 = 8'ha1 == r_count_82_io_out ? io_r_161_b : _GEN_16860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16862 = 8'ha2 == r_count_82_io_out ? io_r_162_b : _GEN_16861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16863 = 8'ha3 == r_count_82_io_out ? io_r_163_b : _GEN_16862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16864 = 8'ha4 == r_count_82_io_out ? io_r_164_b : _GEN_16863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16865 = 8'ha5 == r_count_82_io_out ? io_r_165_b : _GEN_16864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16866 = 8'ha6 == r_count_82_io_out ? io_r_166_b : _GEN_16865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16867 = 8'ha7 == r_count_82_io_out ? io_r_167_b : _GEN_16866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16868 = 8'ha8 == r_count_82_io_out ? io_r_168_b : _GEN_16867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16869 = 8'ha9 == r_count_82_io_out ? io_r_169_b : _GEN_16868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16870 = 8'haa == r_count_82_io_out ? io_r_170_b : _GEN_16869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16871 = 8'hab == r_count_82_io_out ? io_r_171_b : _GEN_16870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16872 = 8'hac == r_count_82_io_out ? io_r_172_b : _GEN_16871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16873 = 8'had == r_count_82_io_out ? io_r_173_b : _GEN_16872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16874 = 8'hae == r_count_82_io_out ? io_r_174_b : _GEN_16873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16875 = 8'haf == r_count_82_io_out ? io_r_175_b : _GEN_16874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16876 = 8'hb0 == r_count_82_io_out ? io_r_176_b : _GEN_16875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16877 = 8'hb1 == r_count_82_io_out ? io_r_177_b : _GEN_16876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16878 = 8'hb2 == r_count_82_io_out ? io_r_178_b : _GEN_16877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16879 = 8'hb3 == r_count_82_io_out ? io_r_179_b : _GEN_16878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16880 = 8'hb4 == r_count_82_io_out ? io_r_180_b : _GEN_16879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16881 = 8'hb5 == r_count_82_io_out ? io_r_181_b : _GEN_16880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16882 = 8'hb6 == r_count_82_io_out ? io_r_182_b : _GEN_16881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16883 = 8'hb7 == r_count_82_io_out ? io_r_183_b : _GEN_16882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16884 = 8'hb8 == r_count_82_io_out ? io_r_184_b : _GEN_16883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16885 = 8'hb9 == r_count_82_io_out ? io_r_185_b : _GEN_16884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16886 = 8'hba == r_count_82_io_out ? io_r_186_b : _GEN_16885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16887 = 8'hbb == r_count_82_io_out ? io_r_187_b : _GEN_16886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16888 = 8'hbc == r_count_82_io_out ? io_r_188_b : _GEN_16887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16889 = 8'hbd == r_count_82_io_out ? io_r_189_b : _GEN_16888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16890 = 8'hbe == r_count_82_io_out ? io_r_190_b : _GEN_16889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16891 = 8'hbf == r_count_82_io_out ? io_r_191_b : _GEN_16890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16892 = 8'hc0 == r_count_82_io_out ? io_r_192_b : _GEN_16891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16893 = 8'hc1 == r_count_82_io_out ? io_r_193_b : _GEN_16892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16894 = 8'hc2 == r_count_82_io_out ? io_r_194_b : _GEN_16893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16895 = 8'hc3 == r_count_82_io_out ? io_r_195_b : _GEN_16894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16896 = 8'hc4 == r_count_82_io_out ? io_r_196_b : _GEN_16895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16897 = 8'hc5 == r_count_82_io_out ? io_r_197_b : _GEN_16896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16898 = 8'hc6 == r_count_82_io_out ? io_r_198_b : _GEN_16897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16901 = 8'h1 == r_count_83_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16902 = 8'h2 == r_count_83_io_out ? io_r_2_b : _GEN_16901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16903 = 8'h3 == r_count_83_io_out ? io_r_3_b : _GEN_16902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16904 = 8'h4 == r_count_83_io_out ? io_r_4_b : _GEN_16903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16905 = 8'h5 == r_count_83_io_out ? io_r_5_b : _GEN_16904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16906 = 8'h6 == r_count_83_io_out ? io_r_6_b : _GEN_16905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16907 = 8'h7 == r_count_83_io_out ? io_r_7_b : _GEN_16906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16908 = 8'h8 == r_count_83_io_out ? io_r_8_b : _GEN_16907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16909 = 8'h9 == r_count_83_io_out ? io_r_9_b : _GEN_16908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16910 = 8'ha == r_count_83_io_out ? io_r_10_b : _GEN_16909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16911 = 8'hb == r_count_83_io_out ? io_r_11_b : _GEN_16910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16912 = 8'hc == r_count_83_io_out ? io_r_12_b : _GEN_16911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16913 = 8'hd == r_count_83_io_out ? io_r_13_b : _GEN_16912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16914 = 8'he == r_count_83_io_out ? io_r_14_b : _GEN_16913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16915 = 8'hf == r_count_83_io_out ? io_r_15_b : _GEN_16914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16916 = 8'h10 == r_count_83_io_out ? io_r_16_b : _GEN_16915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16917 = 8'h11 == r_count_83_io_out ? io_r_17_b : _GEN_16916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16918 = 8'h12 == r_count_83_io_out ? io_r_18_b : _GEN_16917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16919 = 8'h13 == r_count_83_io_out ? io_r_19_b : _GEN_16918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16920 = 8'h14 == r_count_83_io_out ? io_r_20_b : _GEN_16919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16921 = 8'h15 == r_count_83_io_out ? io_r_21_b : _GEN_16920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16922 = 8'h16 == r_count_83_io_out ? io_r_22_b : _GEN_16921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16923 = 8'h17 == r_count_83_io_out ? io_r_23_b : _GEN_16922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16924 = 8'h18 == r_count_83_io_out ? io_r_24_b : _GEN_16923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16925 = 8'h19 == r_count_83_io_out ? io_r_25_b : _GEN_16924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16926 = 8'h1a == r_count_83_io_out ? io_r_26_b : _GEN_16925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16927 = 8'h1b == r_count_83_io_out ? io_r_27_b : _GEN_16926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16928 = 8'h1c == r_count_83_io_out ? io_r_28_b : _GEN_16927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16929 = 8'h1d == r_count_83_io_out ? io_r_29_b : _GEN_16928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16930 = 8'h1e == r_count_83_io_out ? io_r_30_b : _GEN_16929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16931 = 8'h1f == r_count_83_io_out ? io_r_31_b : _GEN_16930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16932 = 8'h20 == r_count_83_io_out ? io_r_32_b : _GEN_16931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16933 = 8'h21 == r_count_83_io_out ? io_r_33_b : _GEN_16932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16934 = 8'h22 == r_count_83_io_out ? io_r_34_b : _GEN_16933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16935 = 8'h23 == r_count_83_io_out ? io_r_35_b : _GEN_16934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16936 = 8'h24 == r_count_83_io_out ? io_r_36_b : _GEN_16935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16937 = 8'h25 == r_count_83_io_out ? io_r_37_b : _GEN_16936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16938 = 8'h26 == r_count_83_io_out ? io_r_38_b : _GEN_16937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16939 = 8'h27 == r_count_83_io_out ? io_r_39_b : _GEN_16938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16940 = 8'h28 == r_count_83_io_out ? io_r_40_b : _GEN_16939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16941 = 8'h29 == r_count_83_io_out ? io_r_41_b : _GEN_16940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16942 = 8'h2a == r_count_83_io_out ? io_r_42_b : _GEN_16941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16943 = 8'h2b == r_count_83_io_out ? io_r_43_b : _GEN_16942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16944 = 8'h2c == r_count_83_io_out ? io_r_44_b : _GEN_16943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16945 = 8'h2d == r_count_83_io_out ? io_r_45_b : _GEN_16944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16946 = 8'h2e == r_count_83_io_out ? io_r_46_b : _GEN_16945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16947 = 8'h2f == r_count_83_io_out ? io_r_47_b : _GEN_16946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16948 = 8'h30 == r_count_83_io_out ? io_r_48_b : _GEN_16947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16949 = 8'h31 == r_count_83_io_out ? io_r_49_b : _GEN_16948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16950 = 8'h32 == r_count_83_io_out ? io_r_50_b : _GEN_16949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16951 = 8'h33 == r_count_83_io_out ? io_r_51_b : _GEN_16950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16952 = 8'h34 == r_count_83_io_out ? io_r_52_b : _GEN_16951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16953 = 8'h35 == r_count_83_io_out ? io_r_53_b : _GEN_16952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16954 = 8'h36 == r_count_83_io_out ? io_r_54_b : _GEN_16953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16955 = 8'h37 == r_count_83_io_out ? io_r_55_b : _GEN_16954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16956 = 8'h38 == r_count_83_io_out ? io_r_56_b : _GEN_16955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16957 = 8'h39 == r_count_83_io_out ? io_r_57_b : _GEN_16956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16958 = 8'h3a == r_count_83_io_out ? io_r_58_b : _GEN_16957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16959 = 8'h3b == r_count_83_io_out ? io_r_59_b : _GEN_16958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16960 = 8'h3c == r_count_83_io_out ? io_r_60_b : _GEN_16959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16961 = 8'h3d == r_count_83_io_out ? io_r_61_b : _GEN_16960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16962 = 8'h3e == r_count_83_io_out ? io_r_62_b : _GEN_16961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16963 = 8'h3f == r_count_83_io_out ? io_r_63_b : _GEN_16962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16964 = 8'h40 == r_count_83_io_out ? io_r_64_b : _GEN_16963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16965 = 8'h41 == r_count_83_io_out ? io_r_65_b : _GEN_16964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16966 = 8'h42 == r_count_83_io_out ? io_r_66_b : _GEN_16965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16967 = 8'h43 == r_count_83_io_out ? io_r_67_b : _GEN_16966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16968 = 8'h44 == r_count_83_io_out ? io_r_68_b : _GEN_16967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16969 = 8'h45 == r_count_83_io_out ? io_r_69_b : _GEN_16968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16970 = 8'h46 == r_count_83_io_out ? io_r_70_b : _GEN_16969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16971 = 8'h47 == r_count_83_io_out ? io_r_71_b : _GEN_16970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16972 = 8'h48 == r_count_83_io_out ? io_r_72_b : _GEN_16971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16973 = 8'h49 == r_count_83_io_out ? io_r_73_b : _GEN_16972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16974 = 8'h4a == r_count_83_io_out ? io_r_74_b : _GEN_16973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16975 = 8'h4b == r_count_83_io_out ? io_r_75_b : _GEN_16974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16976 = 8'h4c == r_count_83_io_out ? io_r_76_b : _GEN_16975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16977 = 8'h4d == r_count_83_io_out ? io_r_77_b : _GEN_16976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16978 = 8'h4e == r_count_83_io_out ? io_r_78_b : _GEN_16977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16979 = 8'h4f == r_count_83_io_out ? io_r_79_b : _GEN_16978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16980 = 8'h50 == r_count_83_io_out ? io_r_80_b : _GEN_16979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16981 = 8'h51 == r_count_83_io_out ? io_r_81_b : _GEN_16980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16982 = 8'h52 == r_count_83_io_out ? io_r_82_b : _GEN_16981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16983 = 8'h53 == r_count_83_io_out ? io_r_83_b : _GEN_16982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16984 = 8'h54 == r_count_83_io_out ? io_r_84_b : _GEN_16983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16985 = 8'h55 == r_count_83_io_out ? io_r_85_b : _GEN_16984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16986 = 8'h56 == r_count_83_io_out ? io_r_86_b : _GEN_16985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16987 = 8'h57 == r_count_83_io_out ? io_r_87_b : _GEN_16986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16988 = 8'h58 == r_count_83_io_out ? io_r_88_b : _GEN_16987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16989 = 8'h59 == r_count_83_io_out ? io_r_89_b : _GEN_16988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16990 = 8'h5a == r_count_83_io_out ? io_r_90_b : _GEN_16989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16991 = 8'h5b == r_count_83_io_out ? io_r_91_b : _GEN_16990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16992 = 8'h5c == r_count_83_io_out ? io_r_92_b : _GEN_16991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16993 = 8'h5d == r_count_83_io_out ? io_r_93_b : _GEN_16992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16994 = 8'h5e == r_count_83_io_out ? io_r_94_b : _GEN_16993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16995 = 8'h5f == r_count_83_io_out ? io_r_95_b : _GEN_16994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16996 = 8'h60 == r_count_83_io_out ? io_r_96_b : _GEN_16995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16997 = 8'h61 == r_count_83_io_out ? io_r_97_b : _GEN_16996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16998 = 8'h62 == r_count_83_io_out ? io_r_98_b : _GEN_16997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_16999 = 8'h63 == r_count_83_io_out ? io_r_99_b : _GEN_16998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17000 = 8'h64 == r_count_83_io_out ? io_r_100_b : _GEN_16999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17001 = 8'h65 == r_count_83_io_out ? io_r_101_b : _GEN_17000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17002 = 8'h66 == r_count_83_io_out ? io_r_102_b : _GEN_17001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17003 = 8'h67 == r_count_83_io_out ? io_r_103_b : _GEN_17002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17004 = 8'h68 == r_count_83_io_out ? io_r_104_b : _GEN_17003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17005 = 8'h69 == r_count_83_io_out ? io_r_105_b : _GEN_17004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17006 = 8'h6a == r_count_83_io_out ? io_r_106_b : _GEN_17005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17007 = 8'h6b == r_count_83_io_out ? io_r_107_b : _GEN_17006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17008 = 8'h6c == r_count_83_io_out ? io_r_108_b : _GEN_17007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17009 = 8'h6d == r_count_83_io_out ? io_r_109_b : _GEN_17008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17010 = 8'h6e == r_count_83_io_out ? io_r_110_b : _GEN_17009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17011 = 8'h6f == r_count_83_io_out ? io_r_111_b : _GEN_17010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17012 = 8'h70 == r_count_83_io_out ? io_r_112_b : _GEN_17011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17013 = 8'h71 == r_count_83_io_out ? io_r_113_b : _GEN_17012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17014 = 8'h72 == r_count_83_io_out ? io_r_114_b : _GEN_17013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17015 = 8'h73 == r_count_83_io_out ? io_r_115_b : _GEN_17014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17016 = 8'h74 == r_count_83_io_out ? io_r_116_b : _GEN_17015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17017 = 8'h75 == r_count_83_io_out ? io_r_117_b : _GEN_17016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17018 = 8'h76 == r_count_83_io_out ? io_r_118_b : _GEN_17017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17019 = 8'h77 == r_count_83_io_out ? io_r_119_b : _GEN_17018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17020 = 8'h78 == r_count_83_io_out ? io_r_120_b : _GEN_17019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17021 = 8'h79 == r_count_83_io_out ? io_r_121_b : _GEN_17020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17022 = 8'h7a == r_count_83_io_out ? io_r_122_b : _GEN_17021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17023 = 8'h7b == r_count_83_io_out ? io_r_123_b : _GEN_17022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17024 = 8'h7c == r_count_83_io_out ? io_r_124_b : _GEN_17023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17025 = 8'h7d == r_count_83_io_out ? io_r_125_b : _GEN_17024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17026 = 8'h7e == r_count_83_io_out ? io_r_126_b : _GEN_17025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17027 = 8'h7f == r_count_83_io_out ? io_r_127_b : _GEN_17026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17028 = 8'h80 == r_count_83_io_out ? io_r_128_b : _GEN_17027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17029 = 8'h81 == r_count_83_io_out ? io_r_129_b : _GEN_17028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17030 = 8'h82 == r_count_83_io_out ? io_r_130_b : _GEN_17029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17031 = 8'h83 == r_count_83_io_out ? io_r_131_b : _GEN_17030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17032 = 8'h84 == r_count_83_io_out ? io_r_132_b : _GEN_17031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17033 = 8'h85 == r_count_83_io_out ? io_r_133_b : _GEN_17032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17034 = 8'h86 == r_count_83_io_out ? io_r_134_b : _GEN_17033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17035 = 8'h87 == r_count_83_io_out ? io_r_135_b : _GEN_17034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17036 = 8'h88 == r_count_83_io_out ? io_r_136_b : _GEN_17035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17037 = 8'h89 == r_count_83_io_out ? io_r_137_b : _GEN_17036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17038 = 8'h8a == r_count_83_io_out ? io_r_138_b : _GEN_17037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17039 = 8'h8b == r_count_83_io_out ? io_r_139_b : _GEN_17038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17040 = 8'h8c == r_count_83_io_out ? io_r_140_b : _GEN_17039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17041 = 8'h8d == r_count_83_io_out ? io_r_141_b : _GEN_17040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17042 = 8'h8e == r_count_83_io_out ? io_r_142_b : _GEN_17041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17043 = 8'h8f == r_count_83_io_out ? io_r_143_b : _GEN_17042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17044 = 8'h90 == r_count_83_io_out ? io_r_144_b : _GEN_17043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17045 = 8'h91 == r_count_83_io_out ? io_r_145_b : _GEN_17044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17046 = 8'h92 == r_count_83_io_out ? io_r_146_b : _GEN_17045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17047 = 8'h93 == r_count_83_io_out ? io_r_147_b : _GEN_17046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17048 = 8'h94 == r_count_83_io_out ? io_r_148_b : _GEN_17047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17049 = 8'h95 == r_count_83_io_out ? io_r_149_b : _GEN_17048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17050 = 8'h96 == r_count_83_io_out ? io_r_150_b : _GEN_17049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17051 = 8'h97 == r_count_83_io_out ? io_r_151_b : _GEN_17050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17052 = 8'h98 == r_count_83_io_out ? io_r_152_b : _GEN_17051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17053 = 8'h99 == r_count_83_io_out ? io_r_153_b : _GEN_17052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17054 = 8'h9a == r_count_83_io_out ? io_r_154_b : _GEN_17053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17055 = 8'h9b == r_count_83_io_out ? io_r_155_b : _GEN_17054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17056 = 8'h9c == r_count_83_io_out ? io_r_156_b : _GEN_17055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17057 = 8'h9d == r_count_83_io_out ? io_r_157_b : _GEN_17056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17058 = 8'h9e == r_count_83_io_out ? io_r_158_b : _GEN_17057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17059 = 8'h9f == r_count_83_io_out ? io_r_159_b : _GEN_17058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17060 = 8'ha0 == r_count_83_io_out ? io_r_160_b : _GEN_17059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17061 = 8'ha1 == r_count_83_io_out ? io_r_161_b : _GEN_17060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17062 = 8'ha2 == r_count_83_io_out ? io_r_162_b : _GEN_17061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17063 = 8'ha3 == r_count_83_io_out ? io_r_163_b : _GEN_17062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17064 = 8'ha4 == r_count_83_io_out ? io_r_164_b : _GEN_17063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17065 = 8'ha5 == r_count_83_io_out ? io_r_165_b : _GEN_17064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17066 = 8'ha6 == r_count_83_io_out ? io_r_166_b : _GEN_17065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17067 = 8'ha7 == r_count_83_io_out ? io_r_167_b : _GEN_17066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17068 = 8'ha8 == r_count_83_io_out ? io_r_168_b : _GEN_17067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17069 = 8'ha9 == r_count_83_io_out ? io_r_169_b : _GEN_17068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17070 = 8'haa == r_count_83_io_out ? io_r_170_b : _GEN_17069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17071 = 8'hab == r_count_83_io_out ? io_r_171_b : _GEN_17070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17072 = 8'hac == r_count_83_io_out ? io_r_172_b : _GEN_17071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17073 = 8'had == r_count_83_io_out ? io_r_173_b : _GEN_17072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17074 = 8'hae == r_count_83_io_out ? io_r_174_b : _GEN_17073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17075 = 8'haf == r_count_83_io_out ? io_r_175_b : _GEN_17074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17076 = 8'hb0 == r_count_83_io_out ? io_r_176_b : _GEN_17075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17077 = 8'hb1 == r_count_83_io_out ? io_r_177_b : _GEN_17076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17078 = 8'hb2 == r_count_83_io_out ? io_r_178_b : _GEN_17077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17079 = 8'hb3 == r_count_83_io_out ? io_r_179_b : _GEN_17078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17080 = 8'hb4 == r_count_83_io_out ? io_r_180_b : _GEN_17079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17081 = 8'hb5 == r_count_83_io_out ? io_r_181_b : _GEN_17080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17082 = 8'hb6 == r_count_83_io_out ? io_r_182_b : _GEN_17081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17083 = 8'hb7 == r_count_83_io_out ? io_r_183_b : _GEN_17082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17084 = 8'hb8 == r_count_83_io_out ? io_r_184_b : _GEN_17083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17085 = 8'hb9 == r_count_83_io_out ? io_r_185_b : _GEN_17084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17086 = 8'hba == r_count_83_io_out ? io_r_186_b : _GEN_17085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17087 = 8'hbb == r_count_83_io_out ? io_r_187_b : _GEN_17086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17088 = 8'hbc == r_count_83_io_out ? io_r_188_b : _GEN_17087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17089 = 8'hbd == r_count_83_io_out ? io_r_189_b : _GEN_17088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17090 = 8'hbe == r_count_83_io_out ? io_r_190_b : _GEN_17089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17091 = 8'hbf == r_count_83_io_out ? io_r_191_b : _GEN_17090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17092 = 8'hc0 == r_count_83_io_out ? io_r_192_b : _GEN_17091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17093 = 8'hc1 == r_count_83_io_out ? io_r_193_b : _GEN_17092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17094 = 8'hc2 == r_count_83_io_out ? io_r_194_b : _GEN_17093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17095 = 8'hc3 == r_count_83_io_out ? io_r_195_b : _GEN_17094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17096 = 8'hc4 == r_count_83_io_out ? io_r_196_b : _GEN_17095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17097 = 8'hc5 == r_count_83_io_out ? io_r_197_b : _GEN_17096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17098 = 8'hc6 == r_count_83_io_out ? io_r_198_b : _GEN_17097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17101 = 8'h1 == r_count_84_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17102 = 8'h2 == r_count_84_io_out ? io_r_2_b : _GEN_17101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17103 = 8'h3 == r_count_84_io_out ? io_r_3_b : _GEN_17102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17104 = 8'h4 == r_count_84_io_out ? io_r_4_b : _GEN_17103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17105 = 8'h5 == r_count_84_io_out ? io_r_5_b : _GEN_17104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17106 = 8'h6 == r_count_84_io_out ? io_r_6_b : _GEN_17105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17107 = 8'h7 == r_count_84_io_out ? io_r_7_b : _GEN_17106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17108 = 8'h8 == r_count_84_io_out ? io_r_8_b : _GEN_17107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17109 = 8'h9 == r_count_84_io_out ? io_r_9_b : _GEN_17108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17110 = 8'ha == r_count_84_io_out ? io_r_10_b : _GEN_17109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17111 = 8'hb == r_count_84_io_out ? io_r_11_b : _GEN_17110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17112 = 8'hc == r_count_84_io_out ? io_r_12_b : _GEN_17111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17113 = 8'hd == r_count_84_io_out ? io_r_13_b : _GEN_17112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17114 = 8'he == r_count_84_io_out ? io_r_14_b : _GEN_17113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17115 = 8'hf == r_count_84_io_out ? io_r_15_b : _GEN_17114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17116 = 8'h10 == r_count_84_io_out ? io_r_16_b : _GEN_17115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17117 = 8'h11 == r_count_84_io_out ? io_r_17_b : _GEN_17116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17118 = 8'h12 == r_count_84_io_out ? io_r_18_b : _GEN_17117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17119 = 8'h13 == r_count_84_io_out ? io_r_19_b : _GEN_17118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17120 = 8'h14 == r_count_84_io_out ? io_r_20_b : _GEN_17119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17121 = 8'h15 == r_count_84_io_out ? io_r_21_b : _GEN_17120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17122 = 8'h16 == r_count_84_io_out ? io_r_22_b : _GEN_17121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17123 = 8'h17 == r_count_84_io_out ? io_r_23_b : _GEN_17122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17124 = 8'h18 == r_count_84_io_out ? io_r_24_b : _GEN_17123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17125 = 8'h19 == r_count_84_io_out ? io_r_25_b : _GEN_17124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17126 = 8'h1a == r_count_84_io_out ? io_r_26_b : _GEN_17125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17127 = 8'h1b == r_count_84_io_out ? io_r_27_b : _GEN_17126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17128 = 8'h1c == r_count_84_io_out ? io_r_28_b : _GEN_17127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17129 = 8'h1d == r_count_84_io_out ? io_r_29_b : _GEN_17128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17130 = 8'h1e == r_count_84_io_out ? io_r_30_b : _GEN_17129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17131 = 8'h1f == r_count_84_io_out ? io_r_31_b : _GEN_17130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17132 = 8'h20 == r_count_84_io_out ? io_r_32_b : _GEN_17131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17133 = 8'h21 == r_count_84_io_out ? io_r_33_b : _GEN_17132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17134 = 8'h22 == r_count_84_io_out ? io_r_34_b : _GEN_17133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17135 = 8'h23 == r_count_84_io_out ? io_r_35_b : _GEN_17134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17136 = 8'h24 == r_count_84_io_out ? io_r_36_b : _GEN_17135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17137 = 8'h25 == r_count_84_io_out ? io_r_37_b : _GEN_17136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17138 = 8'h26 == r_count_84_io_out ? io_r_38_b : _GEN_17137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17139 = 8'h27 == r_count_84_io_out ? io_r_39_b : _GEN_17138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17140 = 8'h28 == r_count_84_io_out ? io_r_40_b : _GEN_17139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17141 = 8'h29 == r_count_84_io_out ? io_r_41_b : _GEN_17140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17142 = 8'h2a == r_count_84_io_out ? io_r_42_b : _GEN_17141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17143 = 8'h2b == r_count_84_io_out ? io_r_43_b : _GEN_17142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17144 = 8'h2c == r_count_84_io_out ? io_r_44_b : _GEN_17143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17145 = 8'h2d == r_count_84_io_out ? io_r_45_b : _GEN_17144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17146 = 8'h2e == r_count_84_io_out ? io_r_46_b : _GEN_17145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17147 = 8'h2f == r_count_84_io_out ? io_r_47_b : _GEN_17146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17148 = 8'h30 == r_count_84_io_out ? io_r_48_b : _GEN_17147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17149 = 8'h31 == r_count_84_io_out ? io_r_49_b : _GEN_17148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17150 = 8'h32 == r_count_84_io_out ? io_r_50_b : _GEN_17149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17151 = 8'h33 == r_count_84_io_out ? io_r_51_b : _GEN_17150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17152 = 8'h34 == r_count_84_io_out ? io_r_52_b : _GEN_17151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17153 = 8'h35 == r_count_84_io_out ? io_r_53_b : _GEN_17152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17154 = 8'h36 == r_count_84_io_out ? io_r_54_b : _GEN_17153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17155 = 8'h37 == r_count_84_io_out ? io_r_55_b : _GEN_17154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17156 = 8'h38 == r_count_84_io_out ? io_r_56_b : _GEN_17155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17157 = 8'h39 == r_count_84_io_out ? io_r_57_b : _GEN_17156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17158 = 8'h3a == r_count_84_io_out ? io_r_58_b : _GEN_17157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17159 = 8'h3b == r_count_84_io_out ? io_r_59_b : _GEN_17158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17160 = 8'h3c == r_count_84_io_out ? io_r_60_b : _GEN_17159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17161 = 8'h3d == r_count_84_io_out ? io_r_61_b : _GEN_17160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17162 = 8'h3e == r_count_84_io_out ? io_r_62_b : _GEN_17161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17163 = 8'h3f == r_count_84_io_out ? io_r_63_b : _GEN_17162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17164 = 8'h40 == r_count_84_io_out ? io_r_64_b : _GEN_17163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17165 = 8'h41 == r_count_84_io_out ? io_r_65_b : _GEN_17164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17166 = 8'h42 == r_count_84_io_out ? io_r_66_b : _GEN_17165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17167 = 8'h43 == r_count_84_io_out ? io_r_67_b : _GEN_17166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17168 = 8'h44 == r_count_84_io_out ? io_r_68_b : _GEN_17167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17169 = 8'h45 == r_count_84_io_out ? io_r_69_b : _GEN_17168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17170 = 8'h46 == r_count_84_io_out ? io_r_70_b : _GEN_17169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17171 = 8'h47 == r_count_84_io_out ? io_r_71_b : _GEN_17170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17172 = 8'h48 == r_count_84_io_out ? io_r_72_b : _GEN_17171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17173 = 8'h49 == r_count_84_io_out ? io_r_73_b : _GEN_17172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17174 = 8'h4a == r_count_84_io_out ? io_r_74_b : _GEN_17173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17175 = 8'h4b == r_count_84_io_out ? io_r_75_b : _GEN_17174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17176 = 8'h4c == r_count_84_io_out ? io_r_76_b : _GEN_17175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17177 = 8'h4d == r_count_84_io_out ? io_r_77_b : _GEN_17176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17178 = 8'h4e == r_count_84_io_out ? io_r_78_b : _GEN_17177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17179 = 8'h4f == r_count_84_io_out ? io_r_79_b : _GEN_17178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17180 = 8'h50 == r_count_84_io_out ? io_r_80_b : _GEN_17179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17181 = 8'h51 == r_count_84_io_out ? io_r_81_b : _GEN_17180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17182 = 8'h52 == r_count_84_io_out ? io_r_82_b : _GEN_17181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17183 = 8'h53 == r_count_84_io_out ? io_r_83_b : _GEN_17182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17184 = 8'h54 == r_count_84_io_out ? io_r_84_b : _GEN_17183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17185 = 8'h55 == r_count_84_io_out ? io_r_85_b : _GEN_17184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17186 = 8'h56 == r_count_84_io_out ? io_r_86_b : _GEN_17185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17187 = 8'h57 == r_count_84_io_out ? io_r_87_b : _GEN_17186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17188 = 8'h58 == r_count_84_io_out ? io_r_88_b : _GEN_17187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17189 = 8'h59 == r_count_84_io_out ? io_r_89_b : _GEN_17188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17190 = 8'h5a == r_count_84_io_out ? io_r_90_b : _GEN_17189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17191 = 8'h5b == r_count_84_io_out ? io_r_91_b : _GEN_17190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17192 = 8'h5c == r_count_84_io_out ? io_r_92_b : _GEN_17191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17193 = 8'h5d == r_count_84_io_out ? io_r_93_b : _GEN_17192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17194 = 8'h5e == r_count_84_io_out ? io_r_94_b : _GEN_17193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17195 = 8'h5f == r_count_84_io_out ? io_r_95_b : _GEN_17194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17196 = 8'h60 == r_count_84_io_out ? io_r_96_b : _GEN_17195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17197 = 8'h61 == r_count_84_io_out ? io_r_97_b : _GEN_17196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17198 = 8'h62 == r_count_84_io_out ? io_r_98_b : _GEN_17197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17199 = 8'h63 == r_count_84_io_out ? io_r_99_b : _GEN_17198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17200 = 8'h64 == r_count_84_io_out ? io_r_100_b : _GEN_17199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17201 = 8'h65 == r_count_84_io_out ? io_r_101_b : _GEN_17200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17202 = 8'h66 == r_count_84_io_out ? io_r_102_b : _GEN_17201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17203 = 8'h67 == r_count_84_io_out ? io_r_103_b : _GEN_17202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17204 = 8'h68 == r_count_84_io_out ? io_r_104_b : _GEN_17203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17205 = 8'h69 == r_count_84_io_out ? io_r_105_b : _GEN_17204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17206 = 8'h6a == r_count_84_io_out ? io_r_106_b : _GEN_17205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17207 = 8'h6b == r_count_84_io_out ? io_r_107_b : _GEN_17206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17208 = 8'h6c == r_count_84_io_out ? io_r_108_b : _GEN_17207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17209 = 8'h6d == r_count_84_io_out ? io_r_109_b : _GEN_17208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17210 = 8'h6e == r_count_84_io_out ? io_r_110_b : _GEN_17209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17211 = 8'h6f == r_count_84_io_out ? io_r_111_b : _GEN_17210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17212 = 8'h70 == r_count_84_io_out ? io_r_112_b : _GEN_17211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17213 = 8'h71 == r_count_84_io_out ? io_r_113_b : _GEN_17212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17214 = 8'h72 == r_count_84_io_out ? io_r_114_b : _GEN_17213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17215 = 8'h73 == r_count_84_io_out ? io_r_115_b : _GEN_17214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17216 = 8'h74 == r_count_84_io_out ? io_r_116_b : _GEN_17215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17217 = 8'h75 == r_count_84_io_out ? io_r_117_b : _GEN_17216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17218 = 8'h76 == r_count_84_io_out ? io_r_118_b : _GEN_17217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17219 = 8'h77 == r_count_84_io_out ? io_r_119_b : _GEN_17218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17220 = 8'h78 == r_count_84_io_out ? io_r_120_b : _GEN_17219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17221 = 8'h79 == r_count_84_io_out ? io_r_121_b : _GEN_17220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17222 = 8'h7a == r_count_84_io_out ? io_r_122_b : _GEN_17221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17223 = 8'h7b == r_count_84_io_out ? io_r_123_b : _GEN_17222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17224 = 8'h7c == r_count_84_io_out ? io_r_124_b : _GEN_17223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17225 = 8'h7d == r_count_84_io_out ? io_r_125_b : _GEN_17224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17226 = 8'h7e == r_count_84_io_out ? io_r_126_b : _GEN_17225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17227 = 8'h7f == r_count_84_io_out ? io_r_127_b : _GEN_17226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17228 = 8'h80 == r_count_84_io_out ? io_r_128_b : _GEN_17227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17229 = 8'h81 == r_count_84_io_out ? io_r_129_b : _GEN_17228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17230 = 8'h82 == r_count_84_io_out ? io_r_130_b : _GEN_17229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17231 = 8'h83 == r_count_84_io_out ? io_r_131_b : _GEN_17230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17232 = 8'h84 == r_count_84_io_out ? io_r_132_b : _GEN_17231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17233 = 8'h85 == r_count_84_io_out ? io_r_133_b : _GEN_17232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17234 = 8'h86 == r_count_84_io_out ? io_r_134_b : _GEN_17233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17235 = 8'h87 == r_count_84_io_out ? io_r_135_b : _GEN_17234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17236 = 8'h88 == r_count_84_io_out ? io_r_136_b : _GEN_17235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17237 = 8'h89 == r_count_84_io_out ? io_r_137_b : _GEN_17236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17238 = 8'h8a == r_count_84_io_out ? io_r_138_b : _GEN_17237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17239 = 8'h8b == r_count_84_io_out ? io_r_139_b : _GEN_17238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17240 = 8'h8c == r_count_84_io_out ? io_r_140_b : _GEN_17239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17241 = 8'h8d == r_count_84_io_out ? io_r_141_b : _GEN_17240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17242 = 8'h8e == r_count_84_io_out ? io_r_142_b : _GEN_17241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17243 = 8'h8f == r_count_84_io_out ? io_r_143_b : _GEN_17242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17244 = 8'h90 == r_count_84_io_out ? io_r_144_b : _GEN_17243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17245 = 8'h91 == r_count_84_io_out ? io_r_145_b : _GEN_17244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17246 = 8'h92 == r_count_84_io_out ? io_r_146_b : _GEN_17245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17247 = 8'h93 == r_count_84_io_out ? io_r_147_b : _GEN_17246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17248 = 8'h94 == r_count_84_io_out ? io_r_148_b : _GEN_17247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17249 = 8'h95 == r_count_84_io_out ? io_r_149_b : _GEN_17248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17250 = 8'h96 == r_count_84_io_out ? io_r_150_b : _GEN_17249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17251 = 8'h97 == r_count_84_io_out ? io_r_151_b : _GEN_17250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17252 = 8'h98 == r_count_84_io_out ? io_r_152_b : _GEN_17251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17253 = 8'h99 == r_count_84_io_out ? io_r_153_b : _GEN_17252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17254 = 8'h9a == r_count_84_io_out ? io_r_154_b : _GEN_17253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17255 = 8'h9b == r_count_84_io_out ? io_r_155_b : _GEN_17254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17256 = 8'h9c == r_count_84_io_out ? io_r_156_b : _GEN_17255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17257 = 8'h9d == r_count_84_io_out ? io_r_157_b : _GEN_17256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17258 = 8'h9e == r_count_84_io_out ? io_r_158_b : _GEN_17257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17259 = 8'h9f == r_count_84_io_out ? io_r_159_b : _GEN_17258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17260 = 8'ha0 == r_count_84_io_out ? io_r_160_b : _GEN_17259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17261 = 8'ha1 == r_count_84_io_out ? io_r_161_b : _GEN_17260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17262 = 8'ha2 == r_count_84_io_out ? io_r_162_b : _GEN_17261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17263 = 8'ha3 == r_count_84_io_out ? io_r_163_b : _GEN_17262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17264 = 8'ha4 == r_count_84_io_out ? io_r_164_b : _GEN_17263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17265 = 8'ha5 == r_count_84_io_out ? io_r_165_b : _GEN_17264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17266 = 8'ha6 == r_count_84_io_out ? io_r_166_b : _GEN_17265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17267 = 8'ha7 == r_count_84_io_out ? io_r_167_b : _GEN_17266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17268 = 8'ha8 == r_count_84_io_out ? io_r_168_b : _GEN_17267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17269 = 8'ha9 == r_count_84_io_out ? io_r_169_b : _GEN_17268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17270 = 8'haa == r_count_84_io_out ? io_r_170_b : _GEN_17269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17271 = 8'hab == r_count_84_io_out ? io_r_171_b : _GEN_17270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17272 = 8'hac == r_count_84_io_out ? io_r_172_b : _GEN_17271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17273 = 8'had == r_count_84_io_out ? io_r_173_b : _GEN_17272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17274 = 8'hae == r_count_84_io_out ? io_r_174_b : _GEN_17273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17275 = 8'haf == r_count_84_io_out ? io_r_175_b : _GEN_17274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17276 = 8'hb0 == r_count_84_io_out ? io_r_176_b : _GEN_17275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17277 = 8'hb1 == r_count_84_io_out ? io_r_177_b : _GEN_17276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17278 = 8'hb2 == r_count_84_io_out ? io_r_178_b : _GEN_17277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17279 = 8'hb3 == r_count_84_io_out ? io_r_179_b : _GEN_17278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17280 = 8'hb4 == r_count_84_io_out ? io_r_180_b : _GEN_17279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17281 = 8'hb5 == r_count_84_io_out ? io_r_181_b : _GEN_17280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17282 = 8'hb6 == r_count_84_io_out ? io_r_182_b : _GEN_17281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17283 = 8'hb7 == r_count_84_io_out ? io_r_183_b : _GEN_17282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17284 = 8'hb8 == r_count_84_io_out ? io_r_184_b : _GEN_17283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17285 = 8'hb9 == r_count_84_io_out ? io_r_185_b : _GEN_17284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17286 = 8'hba == r_count_84_io_out ? io_r_186_b : _GEN_17285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17287 = 8'hbb == r_count_84_io_out ? io_r_187_b : _GEN_17286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17288 = 8'hbc == r_count_84_io_out ? io_r_188_b : _GEN_17287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17289 = 8'hbd == r_count_84_io_out ? io_r_189_b : _GEN_17288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17290 = 8'hbe == r_count_84_io_out ? io_r_190_b : _GEN_17289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17291 = 8'hbf == r_count_84_io_out ? io_r_191_b : _GEN_17290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17292 = 8'hc0 == r_count_84_io_out ? io_r_192_b : _GEN_17291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17293 = 8'hc1 == r_count_84_io_out ? io_r_193_b : _GEN_17292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17294 = 8'hc2 == r_count_84_io_out ? io_r_194_b : _GEN_17293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17295 = 8'hc3 == r_count_84_io_out ? io_r_195_b : _GEN_17294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17296 = 8'hc4 == r_count_84_io_out ? io_r_196_b : _GEN_17295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17297 = 8'hc5 == r_count_84_io_out ? io_r_197_b : _GEN_17296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17298 = 8'hc6 == r_count_84_io_out ? io_r_198_b : _GEN_17297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17301 = 8'h1 == r_count_85_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17302 = 8'h2 == r_count_85_io_out ? io_r_2_b : _GEN_17301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17303 = 8'h3 == r_count_85_io_out ? io_r_3_b : _GEN_17302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17304 = 8'h4 == r_count_85_io_out ? io_r_4_b : _GEN_17303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17305 = 8'h5 == r_count_85_io_out ? io_r_5_b : _GEN_17304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17306 = 8'h6 == r_count_85_io_out ? io_r_6_b : _GEN_17305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17307 = 8'h7 == r_count_85_io_out ? io_r_7_b : _GEN_17306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17308 = 8'h8 == r_count_85_io_out ? io_r_8_b : _GEN_17307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17309 = 8'h9 == r_count_85_io_out ? io_r_9_b : _GEN_17308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17310 = 8'ha == r_count_85_io_out ? io_r_10_b : _GEN_17309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17311 = 8'hb == r_count_85_io_out ? io_r_11_b : _GEN_17310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17312 = 8'hc == r_count_85_io_out ? io_r_12_b : _GEN_17311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17313 = 8'hd == r_count_85_io_out ? io_r_13_b : _GEN_17312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17314 = 8'he == r_count_85_io_out ? io_r_14_b : _GEN_17313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17315 = 8'hf == r_count_85_io_out ? io_r_15_b : _GEN_17314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17316 = 8'h10 == r_count_85_io_out ? io_r_16_b : _GEN_17315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17317 = 8'h11 == r_count_85_io_out ? io_r_17_b : _GEN_17316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17318 = 8'h12 == r_count_85_io_out ? io_r_18_b : _GEN_17317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17319 = 8'h13 == r_count_85_io_out ? io_r_19_b : _GEN_17318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17320 = 8'h14 == r_count_85_io_out ? io_r_20_b : _GEN_17319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17321 = 8'h15 == r_count_85_io_out ? io_r_21_b : _GEN_17320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17322 = 8'h16 == r_count_85_io_out ? io_r_22_b : _GEN_17321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17323 = 8'h17 == r_count_85_io_out ? io_r_23_b : _GEN_17322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17324 = 8'h18 == r_count_85_io_out ? io_r_24_b : _GEN_17323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17325 = 8'h19 == r_count_85_io_out ? io_r_25_b : _GEN_17324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17326 = 8'h1a == r_count_85_io_out ? io_r_26_b : _GEN_17325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17327 = 8'h1b == r_count_85_io_out ? io_r_27_b : _GEN_17326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17328 = 8'h1c == r_count_85_io_out ? io_r_28_b : _GEN_17327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17329 = 8'h1d == r_count_85_io_out ? io_r_29_b : _GEN_17328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17330 = 8'h1e == r_count_85_io_out ? io_r_30_b : _GEN_17329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17331 = 8'h1f == r_count_85_io_out ? io_r_31_b : _GEN_17330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17332 = 8'h20 == r_count_85_io_out ? io_r_32_b : _GEN_17331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17333 = 8'h21 == r_count_85_io_out ? io_r_33_b : _GEN_17332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17334 = 8'h22 == r_count_85_io_out ? io_r_34_b : _GEN_17333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17335 = 8'h23 == r_count_85_io_out ? io_r_35_b : _GEN_17334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17336 = 8'h24 == r_count_85_io_out ? io_r_36_b : _GEN_17335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17337 = 8'h25 == r_count_85_io_out ? io_r_37_b : _GEN_17336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17338 = 8'h26 == r_count_85_io_out ? io_r_38_b : _GEN_17337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17339 = 8'h27 == r_count_85_io_out ? io_r_39_b : _GEN_17338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17340 = 8'h28 == r_count_85_io_out ? io_r_40_b : _GEN_17339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17341 = 8'h29 == r_count_85_io_out ? io_r_41_b : _GEN_17340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17342 = 8'h2a == r_count_85_io_out ? io_r_42_b : _GEN_17341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17343 = 8'h2b == r_count_85_io_out ? io_r_43_b : _GEN_17342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17344 = 8'h2c == r_count_85_io_out ? io_r_44_b : _GEN_17343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17345 = 8'h2d == r_count_85_io_out ? io_r_45_b : _GEN_17344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17346 = 8'h2e == r_count_85_io_out ? io_r_46_b : _GEN_17345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17347 = 8'h2f == r_count_85_io_out ? io_r_47_b : _GEN_17346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17348 = 8'h30 == r_count_85_io_out ? io_r_48_b : _GEN_17347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17349 = 8'h31 == r_count_85_io_out ? io_r_49_b : _GEN_17348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17350 = 8'h32 == r_count_85_io_out ? io_r_50_b : _GEN_17349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17351 = 8'h33 == r_count_85_io_out ? io_r_51_b : _GEN_17350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17352 = 8'h34 == r_count_85_io_out ? io_r_52_b : _GEN_17351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17353 = 8'h35 == r_count_85_io_out ? io_r_53_b : _GEN_17352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17354 = 8'h36 == r_count_85_io_out ? io_r_54_b : _GEN_17353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17355 = 8'h37 == r_count_85_io_out ? io_r_55_b : _GEN_17354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17356 = 8'h38 == r_count_85_io_out ? io_r_56_b : _GEN_17355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17357 = 8'h39 == r_count_85_io_out ? io_r_57_b : _GEN_17356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17358 = 8'h3a == r_count_85_io_out ? io_r_58_b : _GEN_17357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17359 = 8'h3b == r_count_85_io_out ? io_r_59_b : _GEN_17358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17360 = 8'h3c == r_count_85_io_out ? io_r_60_b : _GEN_17359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17361 = 8'h3d == r_count_85_io_out ? io_r_61_b : _GEN_17360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17362 = 8'h3e == r_count_85_io_out ? io_r_62_b : _GEN_17361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17363 = 8'h3f == r_count_85_io_out ? io_r_63_b : _GEN_17362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17364 = 8'h40 == r_count_85_io_out ? io_r_64_b : _GEN_17363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17365 = 8'h41 == r_count_85_io_out ? io_r_65_b : _GEN_17364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17366 = 8'h42 == r_count_85_io_out ? io_r_66_b : _GEN_17365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17367 = 8'h43 == r_count_85_io_out ? io_r_67_b : _GEN_17366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17368 = 8'h44 == r_count_85_io_out ? io_r_68_b : _GEN_17367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17369 = 8'h45 == r_count_85_io_out ? io_r_69_b : _GEN_17368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17370 = 8'h46 == r_count_85_io_out ? io_r_70_b : _GEN_17369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17371 = 8'h47 == r_count_85_io_out ? io_r_71_b : _GEN_17370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17372 = 8'h48 == r_count_85_io_out ? io_r_72_b : _GEN_17371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17373 = 8'h49 == r_count_85_io_out ? io_r_73_b : _GEN_17372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17374 = 8'h4a == r_count_85_io_out ? io_r_74_b : _GEN_17373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17375 = 8'h4b == r_count_85_io_out ? io_r_75_b : _GEN_17374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17376 = 8'h4c == r_count_85_io_out ? io_r_76_b : _GEN_17375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17377 = 8'h4d == r_count_85_io_out ? io_r_77_b : _GEN_17376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17378 = 8'h4e == r_count_85_io_out ? io_r_78_b : _GEN_17377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17379 = 8'h4f == r_count_85_io_out ? io_r_79_b : _GEN_17378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17380 = 8'h50 == r_count_85_io_out ? io_r_80_b : _GEN_17379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17381 = 8'h51 == r_count_85_io_out ? io_r_81_b : _GEN_17380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17382 = 8'h52 == r_count_85_io_out ? io_r_82_b : _GEN_17381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17383 = 8'h53 == r_count_85_io_out ? io_r_83_b : _GEN_17382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17384 = 8'h54 == r_count_85_io_out ? io_r_84_b : _GEN_17383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17385 = 8'h55 == r_count_85_io_out ? io_r_85_b : _GEN_17384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17386 = 8'h56 == r_count_85_io_out ? io_r_86_b : _GEN_17385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17387 = 8'h57 == r_count_85_io_out ? io_r_87_b : _GEN_17386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17388 = 8'h58 == r_count_85_io_out ? io_r_88_b : _GEN_17387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17389 = 8'h59 == r_count_85_io_out ? io_r_89_b : _GEN_17388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17390 = 8'h5a == r_count_85_io_out ? io_r_90_b : _GEN_17389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17391 = 8'h5b == r_count_85_io_out ? io_r_91_b : _GEN_17390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17392 = 8'h5c == r_count_85_io_out ? io_r_92_b : _GEN_17391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17393 = 8'h5d == r_count_85_io_out ? io_r_93_b : _GEN_17392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17394 = 8'h5e == r_count_85_io_out ? io_r_94_b : _GEN_17393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17395 = 8'h5f == r_count_85_io_out ? io_r_95_b : _GEN_17394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17396 = 8'h60 == r_count_85_io_out ? io_r_96_b : _GEN_17395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17397 = 8'h61 == r_count_85_io_out ? io_r_97_b : _GEN_17396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17398 = 8'h62 == r_count_85_io_out ? io_r_98_b : _GEN_17397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17399 = 8'h63 == r_count_85_io_out ? io_r_99_b : _GEN_17398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17400 = 8'h64 == r_count_85_io_out ? io_r_100_b : _GEN_17399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17401 = 8'h65 == r_count_85_io_out ? io_r_101_b : _GEN_17400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17402 = 8'h66 == r_count_85_io_out ? io_r_102_b : _GEN_17401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17403 = 8'h67 == r_count_85_io_out ? io_r_103_b : _GEN_17402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17404 = 8'h68 == r_count_85_io_out ? io_r_104_b : _GEN_17403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17405 = 8'h69 == r_count_85_io_out ? io_r_105_b : _GEN_17404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17406 = 8'h6a == r_count_85_io_out ? io_r_106_b : _GEN_17405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17407 = 8'h6b == r_count_85_io_out ? io_r_107_b : _GEN_17406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17408 = 8'h6c == r_count_85_io_out ? io_r_108_b : _GEN_17407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17409 = 8'h6d == r_count_85_io_out ? io_r_109_b : _GEN_17408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17410 = 8'h6e == r_count_85_io_out ? io_r_110_b : _GEN_17409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17411 = 8'h6f == r_count_85_io_out ? io_r_111_b : _GEN_17410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17412 = 8'h70 == r_count_85_io_out ? io_r_112_b : _GEN_17411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17413 = 8'h71 == r_count_85_io_out ? io_r_113_b : _GEN_17412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17414 = 8'h72 == r_count_85_io_out ? io_r_114_b : _GEN_17413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17415 = 8'h73 == r_count_85_io_out ? io_r_115_b : _GEN_17414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17416 = 8'h74 == r_count_85_io_out ? io_r_116_b : _GEN_17415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17417 = 8'h75 == r_count_85_io_out ? io_r_117_b : _GEN_17416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17418 = 8'h76 == r_count_85_io_out ? io_r_118_b : _GEN_17417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17419 = 8'h77 == r_count_85_io_out ? io_r_119_b : _GEN_17418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17420 = 8'h78 == r_count_85_io_out ? io_r_120_b : _GEN_17419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17421 = 8'h79 == r_count_85_io_out ? io_r_121_b : _GEN_17420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17422 = 8'h7a == r_count_85_io_out ? io_r_122_b : _GEN_17421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17423 = 8'h7b == r_count_85_io_out ? io_r_123_b : _GEN_17422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17424 = 8'h7c == r_count_85_io_out ? io_r_124_b : _GEN_17423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17425 = 8'h7d == r_count_85_io_out ? io_r_125_b : _GEN_17424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17426 = 8'h7e == r_count_85_io_out ? io_r_126_b : _GEN_17425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17427 = 8'h7f == r_count_85_io_out ? io_r_127_b : _GEN_17426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17428 = 8'h80 == r_count_85_io_out ? io_r_128_b : _GEN_17427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17429 = 8'h81 == r_count_85_io_out ? io_r_129_b : _GEN_17428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17430 = 8'h82 == r_count_85_io_out ? io_r_130_b : _GEN_17429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17431 = 8'h83 == r_count_85_io_out ? io_r_131_b : _GEN_17430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17432 = 8'h84 == r_count_85_io_out ? io_r_132_b : _GEN_17431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17433 = 8'h85 == r_count_85_io_out ? io_r_133_b : _GEN_17432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17434 = 8'h86 == r_count_85_io_out ? io_r_134_b : _GEN_17433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17435 = 8'h87 == r_count_85_io_out ? io_r_135_b : _GEN_17434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17436 = 8'h88 == r_count_85_io_out ? io_r_136_b : _GEN_17435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17437 = 8'h89 == r_count_85_io_out ? io_r_137_b : _GEN_17436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17438 = 8'h8a == r_count_85_io_out ? io_r_138_b : _GEN_17437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17439 = 8'h8b == r_count_85_io_out ? io_r_139_b : _GEN_17438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17440 = 8'h8c == r_count_85_io_out ? io_r_140_b : _GEN_17439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17441 = 8'h8d == r_count_85_io_out ? io_r_141_b : _GEN_17440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17442 = 8'h8e == r_count_85_io_out ? io_r_142_b : _GEN_17441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17443 = 8'h8f == r_count_85_io_out ? io_r_143_b : _GEN_17442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17444 = 8'h90 == r_count_85_io_out ? io_r_144_b : _GEN_17443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17445 = 8'h91 == r_count_85_io_out ? io_r_145_b : _GEN_17444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17446 = 8'h92 == r_count_85_io_out ? io_r_146_b : _GEN_17445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17447 = 8'h93 == r_count_85_io_out ? io_r_147_b : _GEN_17446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17448 = 8'h94 == r_count_85_io_out ? io_r_148_b : _GEN_17447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17449 = 8'h95 == r_count_85_io_out ? io_r_149_b : _GEN_17448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17450 = 8'h96 == r_count_85_io_out ? io_r_150_b : _GEN_17449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17451 = 8'h97 == r_count_85_io_out ? io_r_151_b : _GEN_17450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17452 = 8'h98 == r_count_85_io_out ? io_r_152_b : _GEN_17451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17453 = 8'h99 == r_count_85_io_out ? io_r_153_b : _GEN_17452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17454 = 8'h9a == r_count_85_io_out ? io_r_154_b : _GEN_17453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17455 = 8'h9b == r_count_85_io_out ? io_r_155_b : _GEN_17454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17456 = 8'h9c == r_count_85_io_out ? io_r_156_b : _GEN_17455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17457 = 8'h9d == r_count_85_io_out ? io_r_157_b : _GEN_17456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17458 = 8'h9e == r_count_85_io_out ? io_r_158_b : _GEN_17457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17459 = 8'h9f == r_count_85_io_out ? io_r_159_b : _GEN_17458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17460 = 8'ha0 == r_count_85_io_out ? io_r_160_b : _GEN_17459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17461 = 8'ha1 == r_count_85_io_out ? io_r_161_b : _GEN_17460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17462 = 8'ha2 == r_count_85_io_out ? io_r_162_b : _GEN_17461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17463 = 8'ha3 == r_count_85_io_out ? io_r_163_b : _GEN_17462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17464 = 8'ha4 == r_count_85_io_out ? io_r_164_b : _GEN_17463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17465 = 8'ha5 == r_count_85_io_out ? io_r_165_b : _GEN_17464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17466 = 8'ha6 == r_count_85_io_out ? io_r_166_b : _GEN_17465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17467 = 8'ha7 == r_count_85_io_out ? io_r_167_b : _GEN_17466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17468 = 8'ha8 == r_count_85_io_out ? io_r_168_b : _GEN_17467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17469 = 8'ha9 == r_count_85_io_out ? io_r_169_b : _GEN_17468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17470 = 8'haa == r_count_85_io_out ? io_r_170_b : _GEN_17469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17471 = 8'hab == r_count_85_io_out ? io_r_171_b : _GEN_17470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17472 = 8'hac == r_count_85_io_out ? io_r_172_b : _GEN_17471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17473 = 8'had == r_count_85_io_out ? io_r_173_b : _GEN_17472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17474 = 8'hae == r_count_85_io_out ? io_r_174_b : _GEN_17473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17475 = 8'haf == r_count_85_io_out ? io_r_175_b : _GEN_17474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17476 = 8'hb0 == r_count_85_io_out ? io_r_176_b : _GEN_17475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17477 = 8'hb1 == r_count_85_io_out ? io_r_177_b : _GEN_17476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17478 = 8'hb2 == r_count_85_io_out ? io_r_178_b : _GEN_17477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17479 = 8'hb3 == r_count_85_io_out ? io_r_179_b : _GEN_17478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17480 = 8'hb4 == r_count_85_io_out ? io_r_180_b : _GEN_17479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17481 = 8'hb5 == r_count_85_io_out ? io_r_181_b : _GEN_17480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17482 = 8'hb6 == r_count_85_io_out ? io_r_182_b : _GEN_17481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17483 = 8'hb7 == r_count_85_io_out ? io_r_183_b : _GEN_17482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17484 = 8'hb8 == r_count_85_io_out ? io_r_184_b : _GEN_17483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17485 = 8'hb9 == r_count_85_io_out ? io_r_185_b : _GEN_17484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17486 = 8'hba == r_count_85_io_out ? io_r_186_b : _GEN_17485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17487 = 8'hbb == r_count_85_io_out ? io_r_187_b : _GEN_17486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17488 = 8'hbc == r_count_85_io_out ? io_r_188_b : _GEN_17487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17489 = 8'hbd == r_count_85_io_out ? io_r_189_b : _GEN_17488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17490 = 8'hbe == r_count_85_io_out ? io_r_190_b : _GEN_17489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17491 = 8'hbf == r_count_85_io_out ? io_r_191_b : _GEN_17490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17492 = 8'hc0 == r_count_85_io_out ? io_r_192_b : _GEN_17491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17493 = 8'hc1 == r_count_85_io_out ? io_r_193_b : _GEN_17492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17494 = 8'hc2 == r_count_85_io_out ? io_r_194_b : _GEN_17493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17495 = 8'hc3 == r_count_85_io_out ? io_r_195_b : _GEN_17494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17496 = 8'hc4 == r_count_85_io_out ? io_r_196_b : _GEN_17495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17497 = 8'hc5 == r_count_85_io_out ? io_r_197_b : _GEN_17496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17498 = 8'hc6 == r_count_85_io_out ? io_r_198_b : _GEN_17497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17501 = 8'h1 == r_count_86_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17502 = 8'h2 == r_count_86_io_out ? io_r_2_b : _GEN_17501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17503 = 8'h3 == r_count_86_io_out ? io_r_3_b : _GEN_17502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17504 = 8'h4 == r_count_86_io_out ? io_r_4_b : _GEN_17503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17505 = 8'h5 == r_count_86_io_out ? io_r_5_b : _GEN_17504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17506 = 8'h6 == r_count_86_io_out ? io_r_6_b : _GEN_17505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17507 = 8'h7 == r_count_86_io_out ? io_r_7_b : _GEN_17506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17508 = 8'h8 == r_count_86_io_out ? io_r_8_b : _GEN_17507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17509 = 8'h9 == r_count_86_io_out ? io_r_9_b : _GEN_17508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17510 = 8'ha == r_count_86_io_out ? io_r_10_b : _GEN_17509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17511 = 8'hb == r_count_86_io_out ? io_r_11_b : _GEN_17510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17512 = 8'hc == r_count_86_io_out ? io_r_12_b : _GEN_17511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17513 = 8'hd == r_count_86_io_out ? io_r_13_b : _GEN_17512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17514 = 8'he == r_count_86_io_out ? io_r_14_b : _GEN_17513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17515 = 8'hf == r_count_86_io_out ? io_r_15_b : _GEN_17514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17516 = 8'h10 == r_count_86_io_out ? io_r_16_b : _GEN_17515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17517 = 8'h11 == r_count_86_io_out ? io_r_17_b : _GEN_17516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17518 = 8'h12 == r_count_86_io_out ? io_r_18_b : _GEN_17517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17519 = 8'h13 == r_count_86_io_out ? io_r_19_b : _GEN_17518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17520 = 8'h14 == r_count_86_io_out ? io_r_20_b : _GEN_17519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17521 = 8'h15 == r_count_86_io_out ? io_r_21_b : _GEN_17520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17522 = 8'h16 == r_count_86_io_out ? io_r_22_b : _GEN_17521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17523 = 8'h17 == r_count_86_io_out ? io_r_23_b : _GEN_17522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17524 = 8'h18 == r_count_86_io_out ? io_r_24_b : _GEN_17523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17525 = 8'h19 == r_count_86_io_out ? io_r_25_b : _GEN_17524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17526 = 8'h1a == r_count_86_io_out ? io_r_26_b : _GEN_17525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17527 = 8'h1b == r_count_86_io_out ? io_r_27_b : _GEN_17526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17528 = 8'h1c == r_count_86_io_out ? io_r_28_b : _GEN_17527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17529 = 8'h1d == r_count_86_io_out ? io_r_29_b : _GEN_17528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17530 = 8'h1e == r_count_86_io_out ? io_r_30_b : _GEN_17529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17531 = 8'h1f == r_count_86_io_out ? io_r_31_b : _GEN_17530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17532 = 8'h20 == r_count_86_io_out ? io_r_32_b : _GEN_17531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17533 = 8'h21 == r_count_86_io_out ? io_r_33_b : _GEN_17532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17534 = 8'h22 == r_count_86_io_out ? io_r_34_b : _GEN_17533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17535 = 8'h23 == r_count_86_io_out ? io_r_35_b : _GEN_17534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17536 = 8'h24 == r_count_86_io_out ? io_r_36_b : _GEN_17535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17537 = 8'h25 == r_count_86_io_out ? io_r_37_b : _GEN_17536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17538 = 8'h26 == r_count_86_io_out ? io_r_38_b : _GEN_17537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17539 = 8'h27 == r_count_86_io_out ? io_r_39_b : _GEN_17538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17540 = 8'h28 == r_count_86_io_out ? io_r_40_b : _GEN_17539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17541 = 8'h29 == r_count_86_io_out ? io_r_41_b : _GEN_17540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17542 = 8'h2a == r_count_86_io_out ? io_r_42_b : _GEN_17541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17543 = 8'h2b == r_count_86_io_out ? io_r_43_b : _GEN_17542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17544 = 8'h2c == r_count_86_io_out ? io_r_44_b : _GEN_17543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17545 = 8'h2d == r_count_86_io_out ? io_r_45_b : _GEN_17544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17546 = 8'h2e == r_count_86_io_out ? io_r_46_b : _GEN_17545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17547 = 8'h2f == r_count_86_io_out ? io_r_47_b : _GEN_17546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17548 = 8'h30 == r_count_86_io_out ? io_r_48_b : _GEN_17547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17549 = 8'h31 == r_count_86_io_out ? io_r_49_b : _GEN_17548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17550 = 8'h32 == r_count_86_io_out ? io_r_50_b : _GEN_17549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17551 = 8'h33 == r_count_86_io_out ? io_r_51_b : _GEN_17550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17552 = 8'h34 == r_count_86_io_out ? io_r_52_b : _GEN_17551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17553 = 8'h35 == r_count_86_io_out ? io_r_53_b : _GEN_17552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17554 = 8'h36 == r_count_86_io_out ? io_r_54_b : _GEN_17553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17555 = 8'h37 == r_count_86_io_out ? io_r_55_b : _GEN_17554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17556 = 8'h38 == r_count_86_io_out ? io_r_56_b : _GEN_17555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17557 = 8'h39 == r_count_86_io_out ? io_r_57_b : _GEN_17556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17558 = 8'h3a == r_count_86_io_out ? io_r_58_b : _GEN_17557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17559 = 8'h3b == r_count_86_io_out ? io_r_59_b : _GEN_17558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17560 = 8'h3c == r_count_86_io_out ? io_r_60_b : _GEN_17559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17561 = 8'h3d == r_count_86_io_out ? io_r_61_b : _GEN_17560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17562 = 8'h3e == r_count_86_io_out ? io_r_62_b : _GEN_17561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17563 = 8'h3f == r_count_86_io_out ? io_r_63_b : _GEN_17562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17564 = 8'h40 == r_count_86_io_out ? io_r_64_b : _GEN_17563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17565 = 8'h41 == r_count_86_io_out ? io_r_65_b : _GEN_17564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17566 = 8'h42 == r_count_86_io_out ? io_r_66_b : _GEN_17565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17567 = 8'h43 == r_count_86_io_out ? io_r_67_b : _GEN_17566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17568 = 8'h44 == r_count_86_io_out ? io_r_68_b : _GEN_17567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17569 = 8'h45 == r_count_86_io_out ? io_r_69_b : _GEN_17568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17570 = 8'h46 == r_count_86_io_out ? io_r_70_b : _GEN_17569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17571 = 8'h47 == r_count_86_io_out ? io_r_71_b : _GEN_17570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17572 = 8'h48 == r_count_86_io_out ? io_r_72_b : _GEN_17571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17573 = 8'h49 == r_count_86_io_out ? io_r_73_b : _GEN_17572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17574 = 8'h4a == r_count_86_io_out ? io_r_74_b : _GEN_17573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17575 = 8'h4b == r_count_86_io_out ? io_r_75_b : _GEN_17574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17576 = 8'h4c == r_count_86_io_out ? io_r_76_b : _GEN_17575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17577 = 8'h4d == r_count_86_io_out ? io_r_77_b : _GEN_17576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17578 = 8'h4e == r_count_86_io_out ? io_r_78_b : _GEN_17577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17579 = 8'h4f == r_count_86_io_out ? io_r_79_b : _GEN_17578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17580 = 8'h50 == r_count_86_io_out ? io_r_80_b : _GEN_17579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17581 = 8'h51 == r_count_86_io_out ? io_r_81_b : _GEN_17580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17582 = 8'h52 == r_count_86_io_out ? io_r_82_b : _GEN_17581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17583 = 8'h53 == r_count_86_io_out ? io_r_83_b : _GEN_17582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17584 = 8'h54 == r_count_86_io_out ? io_r_84_b : _GEN_17583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17585 = 8'h55 == r_count_86_io_out ? io_r_85_b : _GEN_17584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17586 = 8'h56 == r_count_86_io_out ? io_r_86_b : _GEN_17585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17587 = 8'h57 == r_count_86_io_out ? io_r_87_b : _GEN_17586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17588 = 8'h58 == r_count_86_io_out ? io_r_88_b : _GEN_17587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17589 = 8'h59 == r_count_86_io_out ? io_r_89_b : _GEN_17588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17590 = 8'h5a == r_count_86_io_out ? io_r_90_b : _GEN_17589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17591 = 8'h5b == r_count_86_io_out ? io_r_91_b : _GEN_17590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17592 = 8'h5c == r_count_86_io_out ? io_r_92_b : _GEN_17591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17593 = 8'h5d == r_count_86_io_out ? io_r_93_b : _GEN_17592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17594 = 8'h5e == r_count_86_io_out ? io_r_94_b : _GEN_17593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17595 = 8'h5f == r_count_86_io_out ? io_r_95_b : _GEN_17594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17596 = 8'h60 == r_count_86_io_out ? io_r_96_b : _GEN_17595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17597 = 8'h61 == r_count_86_io_out ? io_r_97_b : _GEN_17596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17598 = 8'h62 == r_count_86_io_out ? io_r_98_b : _GEN_17597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17599 = 8'h63 == r_count_86_io_out ? io_r_99_b : _GEN_17598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17600 = 8'h64 == r_count_86_io_out ? io_r_100_b : _GEN_17599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17601 = 8'h65 == r_count_86_io_out ? io_r_101_b : _GEN_17600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17602 = 8'h66 == r_count_86_io_out ? io_r_102_b : _GEN_17601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17603 = 8'h67 == r_count_86_io_out ? io_r_103_b : _GEN_17602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17604 = 8'h68 == r_count_86_io_out ? io_r_104_b : _GEN_17603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17605 = 8'h69 == r_count_86_io_out ? io_r_105_b : _GEN_17604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17606 = 8'h6a == r_count_86_io_out ? io_r_106_b : _GEN_17605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17607 = 8'h6b == r_count_86_io_out ? io_r_107_b : _GEN_17606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17608 = 8'h6c == r_count_86_io_out ? io_r_108_b : _GEN_17607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17609 = 8'h6d == r_count_86_io_out ? io_r_109_b : _GEN_17608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17610 = 8'h6e == r_count_86_io_out ? io_r_110_b : _GEN_17609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17611 = 8'h6f == r_count_86_io_out ? io_r_111_b : _GEN_17610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17612 = 8'h70 == r_count_86_io_out ? io_r_112_b : _GEN_17611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17613 = 8'h71 == r_count_86_io_out ? io_r_113_b : _GEN_17612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17614 = 8'h72 == r_count_86_io_out ? io_r_114_b : _GEN_17613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17615 = 8'h73 == r_count_86_io_out ? io_r_115_b : _GEN_17614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17616 = 8'h74 == r_count_86_io_out ? io_r_116_b : _GEN_17615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17617 = 8'h75 == r_count_86_io_out ? io_r_117_b : _GEN_17616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17618 = 8'h76 == r_count_86_io_out ? io_r_118_b : _GEN_17617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17619 = 8'h77 == r_count_86_io_out ? io_r_119_b : _GEN_17618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17620 = 8'h78 == r_count_86_io_out ? io_r_120_b : _GEN_17619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17621 = 8'h79 == r_count_86_io_out ? io_r_121_b : _GEN_17620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17622 = 8'h7a == r_count_86_io_out ? io_r_122_b : _GEN_17621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17623 = 8'h7b == r_count_86_io_out ? io_r_123_b : _GEN_17622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17624 = 8'h7c == r_count_86_io_out ? io_r_124_b : _GEN_17623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17625 = 8'h7d == r_count_86_io_out ? io_r_125_b : _GEN_17624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17626 = 8'h7e == r_count_86_io_out ? io_r_126_b : _GEN_17625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17627 = 8'h7f == r_count_86_io_out ? io_r_127_b : _GEN_17626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17628 = 8'h80 == r_count_86_io_out ? io_r_128_b : _GEN_17627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17629 = 8'h81 == r_count_86_io_out ? io_r_129_b : _GEN_17628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17630 = 8'h82 == r_count_86_io_out ? io_r_130_b : _GEN_17629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17631 = 8'h83 == r_count_86_io_out ? io_r_131_b : _GEN_17630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17632 = 8'h84 == r_count_86_io_out ? io_r_132_b : _GEN_17631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17633 = 8'h85 == r_count_86_io_out ? io_r_133_b : _GEN_17632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17634 = 8'h86 == r_count_86_io_out ? io_r_134_b : _GEN_17633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17635 = 8'h87 == r_count_86_io_out ? io_r_135_b : _GEN_17634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17636 = 8'h88 == r_count_86_io_out ? io_r_136_b : _GEN_17635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17637 = 8'h89 == r_count_86_io_out ? io_r_137_b : _GEN_17636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17638 = 8'h8a == r_count_86_io_out ? io_r_138_b : _GEN_17637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17639 = 8'h8b == r_count_86_io_out ? io_r_139_b : _GEN_17638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17640 = 8'h8c == r_count_86_io_out ? io_r_140_b : _GEN_17639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17641 = 8'h8d == r_count_86_io_out ? io_r_141_b : _GEN_17640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17642 = 8'h8e == r_count_86_io_out ? io_r_142_b : _GEN_17641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17643 = 8'h8f == r_count_86_io_out ? io_r_143_b : _GEN_17642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17644 = 8'h90 == r_count_86_io_out ? io_r_144_b : _GEN_17643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17645 = 8'h91 == r_count_86_io_out ? io_r_145_b : _GEN_17644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17646 = 8'h92 == r_count_86_io_out ? io_r_146_b : _GEN_17645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17647 = 8'h93 == r_count_86_io_out ? io_r_147_b : _GEN_17646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17648 = 8'h94 == r_count_86_io_out ? io_r_148_b : _GEN_17647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17649 = 8'h95 == r_count_86_io_out ? io_r_149_b : _GEN_17648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17650 = 8'h96 == r_count_86_io_out ? io_r_150_b : _GEN_17649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17651 = 8'h97 == r_count_86_io_out ? io_r_151_b : _GEN_17650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17652 = 8'h98 == r_count_86_io_out ? io_r_152_b : _GEN_17651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17653 = 8'h99 == r_count_86_io_out ? io_r_153_b : _GEN_17652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17654 = 8'h9a == r_count_86_io_out ? io_r_154_b : _GEN_17653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17655 = 8'h9b == r_count_86_io_out ? io_r_155_b : _GEN_17654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17656 = 8'h9c == r_count_86_io_out ? io_r_156_b : _GEN_17655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17657 = 8'h9d == r_count_86_io_out ? io_r_157_b : _GEN_17656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17658 = 8'h9e == r_count_86_io_out ? io_r_158_b : _GEN_17657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17659 = 8'h9f == r_count_86_io_out ? io_r_159_b : _GEN_17658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17660 = 8'ha0 == r_count_86_io_out ? io_r_160_b : _GEN_17659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17661 = 8'ha1 == r_count_86_io_out ? io_r_161_b : _GEN_17660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17662 = 8'ha2 == r_count_86_io_out ? io_r_162_b : _GEN_17661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17663 = 8'ha3 == r_count_86_io_out ? io_r_163_b : _GEN_17662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17664 = 8'ha4 == r_count_86_io_out ? io_r_164_b : _GEN_17663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17665 = 8'ha5 == r_count_86_io_out ? io_r_165_b : _GEN_17664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17666 = 8'ha6 == r_count_86_io_out ? io_r_166_b : _GEN_17665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17667 = 8'ha7 == r_count_86_io_out ? io_r_167_b : _GEN_17666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17668 = 8'ha8 == r_count_86_io_out ? io_r_168_b : _GEN_17667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17669 = 8'ha9 == r_count_86_io_out ? io_r_169_b : _GEN_17668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17670 = 8'haa == r_count_86_io_out ? io_r_170_b : _GEN_17669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17671 = 8'hab == r_count_86_io_out ? io_r_171_b : _GEN_17670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17672 = 8'hac == r_count_86_io_out ? io_r_172_b : _GEN_17671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17673 = 8'had == r_count_86_io_out ? io_r_173_b : _GEN_17672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17674 = 8'hae == r_count_86_io_out ? io_r_174_b : _GEN_17673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17675 = 8'haf == r_count_86_io_out ? io_r_175_b : _GEN_17674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17676 = 8'hb0 == r_count_86_io_out ? io_r_176_b : _GEN_17675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17677 = 8'hb1 == r_count_86_io_out ? io_r_177_b : _GEN_17676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17678 = 8'hb2 == r_count_86_io_out ? io_r_178_b : _GEN_17677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17679 = 8'hb3 == r_count_86_io_out ? io_r_179_b : _GEN_17678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17680 = 8'hb4 == r_count_86_io_out ? io_r_180_b : _GEN_17679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17681 = 8'hb5 == r_count_86_io_out ? io_r_181_b : _GEN_17680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17682 = 8'hb6 == r_count_86_io_out ? io_r_182_b : _GEN_17681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17683 = 8'hb7 == r_count_86_io_out ? io_r_183_b : _GEN_17682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17684 = 8'hb8 == r_count_86_io_out ? io_r_184_b : _GEN_17683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17685 = 8'hb9 == r_count_86_io_out ? io_r_185_b : _GEN_17684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17686 = 8'hba == r_count_86_io_out ? io_r_186_b : _GEN_17685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17687 = 8'hbb == r_count_86_io_out ? io_r_187_b : _GEN_17686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17688 = 8'hbc == r_count_86_io_out ? io_r_188_b : _GEN_17687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17689 = 8'hbd == r_count_86_io_out ? io_r_189_b : _GEN_17688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17690 = 8'hbe == r_count_86_io_out ? io_r_190_b : _GEN_17689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17691 = 8'hbf == r_count_86_io_out ? io_r_191_b : _GEN_17690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17692 = 8'hc0 == r_count_86_io_out ? io_r_192_b : _GEN_17691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17693 = 8'hc1 == r_count_86_io_out ? io_r_193_b : _GEN_17692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17694 = 8'hc2 == r_count_86_io_out ? io_r_194_b : _GEN_17693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17695 = 8'hc3 == r_count_86_io_out ? io_r_195_b : _GEN_17694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17696 = 8'hc4 == r_count_86_io_out ? io_r_196_b : _GEN_17695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17697 = 8'hc5 == r_count_86_io_out ? io_r_197_b : _GEN_17696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17698 = 8'hc6 == r_count_86_io_out ? io_r_198_b : _GEN_17697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17701 = 8'h1 == r_count_87_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17702 = 8'h2 == r_count_87_io_out ? io_r_2_b : _GEN_17701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17703 = 8'h3 == r_count_87_io_out ? io_r_3_b : _GEN_17702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17704 = 8'h4 == r_count_87_io_out ? io_r_4_b : _GEN_17703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17705 = 8'h5 == r_count_87_io_out ? io_r_5_b : _GEN_17704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17706 = 8'h6 == r_count_87_io_out ? io_r_6_b : _GEN_17705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17707 = 8'h7 == r_count_87_io_out ? io_r_7_b : _GEN_17706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17708 = 8'h8 == r_count_87_io_out ? io_r_8_b : _GEN_17707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17709 = 8'h9 == r_count_87_io_out ? io_r_9_b : _GEN_17708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17710 = 8'ha == r_count_87_io_out ? io_r_10_b : _GEN_17709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17711 = 8'hb == r_count_87_io_out ? io_r_11_b : _GEN_17710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17712 = 8'hc == r_count_87_io_out ? io_r_12_b : _GEN_17711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17713 = 8'hd == r_count_87_io_out ? io_r_13_b : _GEN_17712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17714 = 8'he == r_count_87_io_out ? io_r_14_b : _GEN_17713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17715 = 8'hf == r_count_87_io_out ? io_r_15_b : _GEN_17714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17716 = 8'h10 == r_count_87_io_out ? io_r_16_b : _GEN_17715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17717 = 8'h11 == r_count_87_io_out ? io_r_17_b : _GEN_17716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17718 = 8'h12 == r_count_87_io_out ? io_r_18_b : _GEN_17717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17719 = 8'h13 == r_count_87_io_out ? io_r_19_b : _GEN_17718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17720 = 8'h14 == r_count_87_io_out ? io_r_20_b : _GEN_17719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17721 = 8'h15 == r_count_87_io_out ? io_r_21_b : _GEN_17720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17722 = 8'h16 == r_count_87_io_out ? io_r_22_b : _GEN_17721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17723 = 8'h17 == r_count_87_io_out ? io_r_23_b : _GEN_17722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17724 = 8'h18 == r_count_87_io_out ? io_r_24_b : _GEN_17723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17725 = 8'h19 == r_count_87_io_out ? io_r_25_b : _GEN_17724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17726 = 8'h1a == r_count_87_io_out ? io_r_26_b : _GEN_17725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17727 = 8'h1b == r_count_87_io_out ? io_r_27_b : _GEN_17726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17728 = 8'h1c == r_count_87_io_out ? io_r_28_b : _GEN_17727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17729 = 8'h1d == r_count_87_io_out ? io_r_29_b : _GEN_17728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17730 = 8'h1e == r_count_87_io_out ? io_r_30_b : _GEN_17729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17731 = 8'h1f == r_count_87_io_out ? io_r_31_b : _GEN_17730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17732 = 8'h20 == r_count_87_io_out ? io_r_32_b : _GEN_17731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17733 = 8'h21 == r_count_87_io_out ? io_r_33_b : _GEN_17732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17734 = 8'h22 == r_count_87_io_out ? io_r_34_b : _GEN_17733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17735 = 8'h23 == r_count_87_io_out ? io_r_35_b : _GEN_17734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17736 = 8'h24 == r_count_87_io_out ? io_r_36_b : _GEN_17735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17737 = 8'h25 == r_count_87_io_out ? io_r_37_b : _GEN_17736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17738 = 8'h26 == r_count_87_io_out ? io_r_38_b : _GEN_17737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17739 = 8'h27 == r_count_87_io_out ? io_r_39_b : _GEN_17738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17740 = 8'h28 == r_count_87_io_out ? io_r_40_b : _GEN_17739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17741 = 8'h29 == r_count_87_io_out ? io_r_41_b : _GEN_17740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17742 = 8'h2a == r_count_87_io_out ? io_r_42_b : _GEN_17741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17743 = 8'h2b == r_count_87_io_out ? io_r_43_b : _GEN_17742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17744 = 8'h2c == r_count_87_io_out ? io_r_44_b : _GEN_17743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17745 = 8'h2d == r_count_87_io_out ? io_r_45_b : _GEN_17744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17746 = 8'h2e == r_count_87_io_out ? io_r_46_b : _GEN_17745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17747 = 8'h2f == r_count_87_io_out ? io_r_47_b : _GEN_17746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17748 = 8'h30 == r_count_87_io_out ? io_r_48_b : _GEN_17747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17749 = 8'h31 == r_count_87_io_out ? io_r_49_b : _GEN_17748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17750 = 8'h32 == r_count_87_io_out ? io_r_50_b : _GEN_17749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17751 = 8'h33 == r_count_87_io_out ? io_r_51_b : _GEN_17750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17752 = 8'h34 == r_count_87_io_out ? io_r_52_b : _GEN_17751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17753 = 8'h35 == r_count_87_io_out ? io_r_53_b : _GEN_17752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17754 = 8'h36 == r_count_87_io_out ? io_r_54_b : _GEN_17753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17755 = 8'h37 == r_count_87_io_out ? io_r_55_b : _GEN_17754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17756 = 8'h38 == r_count_87_io_out ? io_r_56_b : _GEN_17755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17757 = 8'h39 == r_count_87_io_out ? io_r_57_b : _GEN_17756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17758 = 8'h3a == r_count_87_io_out ? io_r_58_b : _GEN_17757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17759 = 8'h3b == r_count_87_io_out ? io_r_59_b : _GEN_17758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17760 = 8'h3c == r_count_87_io_out ? io_r_60_b : _GEN_17759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17761 = 8'h3d == r_count_87_io_out ? io_r_61_b : _GEN_17760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17762 = 8'h3e == r_count_87_io_out ? io_r_62_b : _GEN_17761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17763 = 8'h3f == r_count_87_io_out ? io_r_63_b : _GEN_17762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17764 = 8'h40 == r_count_87_io_out ? io_r_64_b : _GEN_17763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17765 = 8'h41 == r_count_87_io_out ? io_r_65_b : _GEN_17764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17766 = 8'h42 == r_count_87_io_out ? io_r_66_b : _GEN_17765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17767 = 8'h43 == r_count_87_io_out ? io_r_67_b : _GEN_17766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17768 = 8'h44 == r_count_87_io_out ? io_r_68_b : _GEN_17767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17769 = 8'h45 == r_count_87_io_out ? io_r_69_b : _GEN_17768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17770 = 8'h46 == r_count_87_io_out ? io_r_70_b : _GEN_17769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17771 = 8'h47 == r_count_87_io_out ? io_r_71_b : _GEN_17770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17772 = 8'h48 == r_count_87_io_out ? io_r_72_b : _GEN_17771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17773 = 8'h49 == r_count_87_io_out ? io_r_73_b : _GEN_17772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17774 = 8'h4a == r_count_87_io_out ? io_r_74_b : _GEN_17773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17775 = 8'h4b == r_count_87_io_out ? io_r_75_b : _GEN_17774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17776 = 8'h4c == r_count_87_io_out ? io_r_76_b : _GEN_17775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17777 = 8'h4d == r_count_87_io_out ? io_r_77_b : _GEN_17776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17778 = 8'h4e == r_count_87_io_out ? io_r_78_b : _GEN_17777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17779 = 8'h4f == r_count_87_io_out ? io_r_79_b : _GEN_17778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17780 = 8'h50 == r_count_87_io_out ? io_r_80_b : _GEN_17779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17781 = 8'h51 == r_count_87_io_out ? io_r_81_b : _GEN_17780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17782 = 8'h52 == r_count_87_io_out ? io_r_82_b : _GEN_17781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17783 = 8'h53 == r_count_87_io_out ? io_r_83_b : _GEN_17782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17784 = 8'h54 == r_count_87_io_out ? io_r_84_b : _GEN_17783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17785 = 8'h55 == r_count_87_io_out ? io_r_85_b : _GEN_17784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17786 = 8'h56 == r_count_87_io_out ? io_r_86_b : _GEN_17785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17787 = 8'h57 == r_count_87_io_out ? io_r_87_b : _GEN_17786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17788 = 8'h58 == r_count_87_io_out ? io_r_88_b : _GEN_17787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17789 = 8'h59 == r_count_87_io_out ? io_r_89_b : _GEN_17788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17790 = 8'h5a == r_count_87_io_out ? io_r_90_b : _GEN_17789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17791 = 8'h5b == r_count_87_io_out ? io_r_91_b : _GEN_17790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17792 = 8'h5c == r_count_87_io_out ? io_r_92_b : _GEN_17791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17793 = 8'h5d == r_count_87_io_out ? io_r_93_b : _GEN_17792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17794 = 8'h5e == r_count_87_io_out ? io_r_94_b : _GEN_17793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17795 = 8'h5f == r_count_87_io_out ? io_r_95_b : _GEN_17794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17796 = 8'h60 == r_count_87_io_out ? io_r_96_b : _GEN_17795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17797 = 8'h61 == r_count_87_io_out ? io_r_97_b : _GEN_17796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17798 = 8'h62 == r_count_87_io_out ? io_r_98_b : _GEN_17797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17799 = 8'h63 == r_count_87_io_out ? io_r_99_b : _GEN_17798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17800 = 8'h64 == r_count_87_io_out ? io_r_100_b : _GEN_17799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17801 = 8'h65 == r_count_87_io_out ? io_r_101_b : _GEN_17800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17802 = 8'h66 == r_count_87_io_out ? io_r_102_b : _GEN_17801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17803 = 8'h67 == r_count_87_io_out ? io_r_103_b : _GEN_17802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17804 = 8'h68 == r_count_87_io_out ? io_r_104_b : _GEN_17803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17805 = 8'h69 == r_count_87_io_out ? io_r_105_b : _GEN_17804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17806 = 8'h6a == r_count_87_io_out ? io_r_106_b : _GEN_17805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17807 = 8'h6b == r_count_87_io_out ? io_r_107_b : _GEN_17806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17808 = 8'h6c == r_count_87_io_out ? io_r_108_b : _GEN_17807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17809 = 8'h6d == r_count_87_io_out ? io_r_109_b : _GEN_17808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17810 = 8'h6e == r_count_87_io_out ? io_r_110_b : _GEN_17809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17811 = 8'h6f == r_count_87_io_out ? io_r_111_b : _GEN_17810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17812 = 8'h70 == r_count_87_io_out ? io_r_112_b : _GEN_17811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17813 = 8'h71 == r_count_87_io_out ? io_r_113_b : _GEN_17812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17814 = 8'h72 == r_count_87_io_out ? io_r_114_b : _GEN_17813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17815 = 8'h73 == r_count_87_io_out ? io_r_115_b : _GEN_17814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17816 = 8'h74 == r_count_87_io_out ? io_r_116_b : _GEN_17815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17817 = 8'h75 == r_count_87_io_out ? io_r_117_b : _GEN_17816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17818 = 8'h76 == r_count_87_io_out ? io_r_118_b : _GEN_17817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17819 = 8'h77 == r_count_87_io_out ? io_r_119_b : _GEN_17818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17820 = 8'h78 == r_count_87_io_out ? io_r_120_b : _GEN_17819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17821 = 8'h79 == r_count_87_io_out ? io_r_121_b : _GEN_17820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17822 = 8'h7a == r_count_87_io_out ? io_r_122_b : _GEN_17821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17823 = 8'h7b == r_count_87_io_out ? io_r_123_b : _GEN_17822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17824 = 8'h7c == r_count_87_io_out ? io_r_124_b : _GEN_17823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17825 = 8'h7d == r_count_87_io_out ? io_r_125_b : _GEN_17824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17826 = 8'h7e == r_count_87_io_out ? io_r_126_b : _GEN_17825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17827 = 8'h7f == r_count_87_io_out ? io_r_127_b : _GEN_17826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17828 = 8'h80 == r_count_87_io_out ? io_r_128_b : _GEN_17827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17829 = 8'h81 == r_count_87_io_out ? io_r_129_b : _GEN_17828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17830 = 8'h82 == r_count_87_io_out ? io_r_130_b : _GEN_17829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17831 = 8'h83 == r_count_87_io_out ? io_r_131_b : _GEN_17830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17832 = 8'h84 == r_count_87_io_out ? io_r_132_b : _GEN_17831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17833 = 8'h85 == r_count_87_io_out ? io_r_133_b : _GEN_17832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17834 = 8'h86 == r_count_87_io_out ? io_r_134_b : _GEN_17833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17835 = 8'h87 == r_count_87_io_out ? io_r_135_b : _GEN_17834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17836 = 8'h88 == r_count_87_io_out ? io_r_136_b : _GEN_17835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17837 = 8'h89 == r_count_87_io_out ? io_r_137_b : _GEN_17836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17838 = 8'h8a == r_count_87_io_out ? io_r_138_b : _GEN_17837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17839 = 8'h8b == r_count_87_io_out ? io_r_139_b : _GEN_17838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17840 = 8'h8c == r_count_87_io_out ? io_r_140_b : _GEN_17839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17841 = 8'h8d == r_count_87_io_out ? io_r_141_b : _GEN_17840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17842 = 8'h8e == r_count_87_io_out ? io_r_142_b : _GEN_17841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17843 = 8'h8f == r_count_87_io_out ? io_r_143_b : _GEN_17842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17844 = 8'h90 == r_count_87_io_out ? io_r_144_b : _GEN_17843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17845 = 8'h91 == r_count_87_io_out ? io_r_145_b : _GEN_17844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17846 = 8'h92 == r_count_87_io_out ? io_r_146_b : _GEN_17845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17847 = 8'h93 == r_count_87_io_out ? io_r_147_b : _GEN_17846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17848 = 8'h94 == r_count_87_io_out ? io_r_148_b : _GEN_17847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17849 = 8'h95 == r_count_87_io_out ? io_r_149_b : _GEN_17848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17850 = 8'h96 == r_count_87_io_out ? io_r_150_b : _GEN_17849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17851 = 8'h97 == r_count_87_io_out ? io_r_151_b : _GEN_17850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17852 = 8'h98 == r_count_87_io_out ? io_r_152_b : _GEN_17851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17853 = 8'h99 == r_count_87_io_out ? io_r_153_b : _GEN_17852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17854 = 8'h9a == r_count_87_io_out ? io_r_154_b : _GEN_17853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17855 = 8'h9b == r_count_87_io_out ? io_r_155_b : _GEN_17854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17856 = 8'h9c == r_count_87_io_out ? io_r_156_b : _GEN_17855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17857 = 8'h9d == r_count_87_io_out ? io_r_157_b : _GEN_17856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17858 = 8'h9e == r_count_87_io_out ? io_r_158_b : _GEN_17857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17859 = 8'h9f == r_count_87_io_out ? io_r_159_b : _GEN_17858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17860 = 8'ha0 == r_count_87_io_out ? io_r_160_b : _GEN_17859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17861 = 8'ha1 == r_count_87_io_out ? io_r_161_b : _GEN_17860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17862 = 8'ha2 == r_count_87_io_out ? io_r_162_b : _GEN_17861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17863 = 8'ha3 == r_count_87_io_out ? io_r_163_b : _GEN_17862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17864 = 8'ha4 == r_count_87_io_out ? io_r_164_b : _GEN_17863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17865 = 8'ha5 == r_count_87_io_out ? io_r_165_b : _GEN_17864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17866 = 8'ha6 == r_count_87_io_out ? io_r_166_b : _GEN_17865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17867 = 8'ha7 == r_count_87_io_out ? io_r_167_b : _GEN_17866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17868 = 8'ha8 == r_count_87_io_out ? io_r_168_b : _GEN_17867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17869 = 8'ha9 == r_count_87_io_out ? io_r_169_b : _GEN_17868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17870 = 8'haa == r_count_87_io_out ? io_r_170_b : _GEN_17869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17871 = 8'hab == r_count_87_io_out ? io_r_171_b : _GEN_17870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17872 = 8'hac == r_count_87_io_out ? io_r_172_b : _GEN_17871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17873 = 8'had == r_count_87_io_out ? io_r_173_b : _GEN_17872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17874 = 8'hae == r_count_87_io_out ? io_r_174_b : _GEN_17873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17875 = 8'haf == r_count_87_io_out ? io_r_175_b : _GEN_17874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17876 = 8'hb0 == r_count_87_io_out ? io_r_176_b : _GEN_17875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17877 = 8'hb1 == r_count_87_io_out ? io_r_177_b : _GEN_17876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17878 = 8'hb2 == r_count_87_io_out ? io_r_178_b : _GEN_17877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17879 = 8'hb3 == r_count_87_io_out ? io_r_179_b : _GEN_17878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17880 = 8'hb4 == r_count_87_io_out ? io_r_180_b : _GEN_17879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17881 = 8'hb5 == r_count_87_io_out ? io_r_181_b : _GEN_17880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17882 = 8'hb6 == r_count_87_io_out ? io_r_182_b : _GEN_17881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17883 = 8'hb7 == r_count_87_io_out ? io_r_183_b : _GEN_17882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17884 = 8'hb8 == r_count_87_io_out ? io_r_184_b : _GEN_17883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17885 = 8'hb9 == r_count_87_io_out ? io_r_185_b : _GEN_17884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17886 = 8'hba == r_count_87_io_out ? io_r_186_b : _GEN_17885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17887 = 8'hbb == r_count_87_io_out ? io_r_187_b : _GEN_17886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17888 = 8'hbc == r_count_87_io_out ? io_r_188_b : _GEN_17887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17889 = 8'hbd == r_count_87_io_out ? io_r_189_b : _GEN_17888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17890 = 8'hbe == r_count_87_io_out ? io_r_190_b : _GEN_17889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17891 = 8'hbf == r_count_87_io_out ? io_r_191_b : _GEN_17890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17892 = 8'hc0 == r_count_87_io_out ? io_r_192_b : _GEN_17891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17893 = 8'hc1 == r_count_87_io_out ? io_r_193_b : _GEN_17892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17894 = 8'hc2 == r_count_87_io_out ? io_r_194_b : _GEN_17893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17895 = 8'hc3 == r_count_87_io_out ? io_r_195_b : _GEN_17894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17896 = 8'hc4 == r_count_87_io_out ? io_r_196_b : _GEN_17895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17897 = 8'hc5 == r_count_87_io_out ? io_r_197_b : _GEN_17896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17898 = 8'hc6 == r_count_87_io_out ? io_r_198_b : _GEN_17897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17901 = 8'h1 == r_count_88_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17902 = 8'h2 == r_count_88_io_out ? io_r_2_b : _GEN_17901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17903 = 8'h3 == r_count_88_io_out ? io_r_3_b : _GEN_17902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17904 = 8'h4 == r_count_88_io_out ? io_r_4_b : _GEN_17903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17905 = 8'h5 == r_count_88_io_out ? io_r_5_b : _GEN_17904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17906 = 8'h6 == r_count_88_io_out ? io_r_6_b : _GEN_17905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17907 = 8'h7 == r_count_88_io_out ? io_r_7_b : _GEN_17906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17908 = 8'h8 == r_count_88_io_out ? io_r_8_b : _GEN_17907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17909 = 8'h9 == r_count_88_io_out ? io_r_9_b : _GEN_17908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17910 = 8'ha == r_count_88_io_out ? io_r_10_b : _GEN_17909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17911 = 8'hb == r_count_88_io_out ? io_r_11_b : _GEN_17910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17912 = 8'hc == r_count_88_io_out ? io_r_12_b : _GEN_17911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17913 = 8'hd == r_count_88_io_out ? io_r_13_b : _GEN_17912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17914 = 8'he == r_count_88_io_out ? io_r_14_b : _GEN_17913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17915 = 8'hf == r_count_88_io_out ? io_r_15_b : _GEN_17914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17916 = 8'h10 == r_count_88_io_out ? io_r_16_b : _GEN_17915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17917 = 8'h11 == r_count_88_io_out ? io_r_17_b : _GEN_17916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17918 = 8'h12 == r_count_88_io_out ? io_r_18_b : _GEN_17917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17919 = 8'h13 == r_count_88_io_out ? io_r_19_b : _GEN_17918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17920 = 8'h14 == r_count_88_io_out ? io_r_20_b : _GEN_17919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17921 = 8'h15 == r_count_88_io_out ? io_r_21_b : _GEN_17920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17922 = 8'h16 == r_count_88_io_out ? io_r_22_b : _GEN_17921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17923 = 8'h17 == r_count_88_io_out ? io_r_23_b : _GEN_17922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17924 = 8'h18 == r_count_88_io_out ? io_r_24_b : _GEN_17923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17925 = 8'h19 == r_count_88_io_out ? io_r_25_b : _GEN_17924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17926 = 8'h1a == r_count_88_io_out ? io_r_26_b : _GEN_17925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17927 = 8'h1b == r_count_88_io_out ? io_r_27_b : _GEN_17926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17928 = 8'h1c == r_count_88_io_out ? io_r_28_b : _GEN_17927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17929 = 8'h1d == r_count_88_io_out ? io_r_29_b : _GEN_17928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17930 = 8'h1e == r_count_88_io_out ? io_r_30_b : _GEN_17929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17931 = 8'h1f == r_count_88_io_out ? io_r_31_b : _GEN_17930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17932 = 8'h20 == r_count_88_io_out ? io_r_32_b : _GEN_17931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17933 = 8'h21 == r_count_88_io_out ? io_r_33_b : _GEN_17932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17934 = 8'h22 == r_count_88_io_out ? io_r_34_b : _GEN_17933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17935 = 8'h23 == r_count_88_io_out ? io_r_35_b : _GEN_17934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17936 = 8'h24 == r_count_88_io_out ? io_r_36_b : _GEN_17935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17937 = 8'h25 == r_count_88_io_out ? io_r_37_b : _GEN_17936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17938 = 8'h26 == r_count_88_io_out ? io_r_38_b : _GEN_17937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17939 = 8'h27 == r_count_88_io_out ? io_r_39_b : _GEN_17938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17940 = 8'h28 == r_count_88_io_out ? io_r_40_b : _GEN_17939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17941 = 8'h29 == r_count_88_io_out ? io_r_41_b : _GEN_17940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17942 = 8'h2a == r_count_88_io_out ? io_r_42_b : _GEN_17941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17943 = 8'h2b == r_count_88_io_out ? io_r_43_b : _GEN_17942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17944 = 8'h2c == r_count_88_io_out ? io_r_44_b : _GEN_17943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17945 = 8'h2d == r_count_88_io_out ? io_r_45_b : _GEN_17944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17946 = 8'h2e == r_count_88_io_out ? io_r_46_b : _GEN_17945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17947 = 8'h2f == r_count_88_io_out ? io_r_47_b : _GEN_17946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17948 = 8'h30 == r_count_88_io_out ? io_r_48_b : _GEN_17947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17949 = 8'h31 == r_count_88_io_out ? io_r_49_b : _GEN_17948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17950 = 8'h32 == r_count_88_io_out ? io_r_50_b : _GEN_17949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17951 = 8'h33 == r_count_88_io_out ? io_r_51_b : _GEN_17950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17952 = 8'h34 == r_count_88_io_out ? io_r_52_b : _GEN_17951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17953 = 8'h35 == r_count_88_io_out ? io_r_53_b : _GEN_17952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17954 = 8'h36 == r_count_88_io_out ? io_r_54_b : _GEN_17953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17955 = 8'h37 == r_count_88_io_out ? io_r_55_b : _GEN_17954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17956 = 8'h38 == r_count_88_io_out ? io_r_56_b : _GEN_17955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17957 = 8'h39 == r_count_88_io_out ? io_r_57_b : _GEN_17956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17958 = 8'h3a == r_count_88_io_out ? io_r_58_b : _GEN_17957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17959 = 8'h3b == r_count_88_io_out ? io_r_59_b : _GEN_17958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17960 = 8'h3c == r_count_88_io_out ? io_r_60_b : _GEN_17959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17961 = 8'h3d == r_count_88_io_out ? io_r_61_b : _GEN_17960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17962 = 8'h3e == r_count_88_io_out ? io_r_62_b : _GEN_17961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17963 = 8'h3f == r_count_88_io_out ? io_r_63_b : _GEN_17962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17964 = 8'h40 == r_count_88_io_out ? io_r_64_b : _GEN_17963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17965 = 8'h41 == r_count_88_io_out ? io_r_65_b : _GEN_17964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17966 = 8'h42 == r_count_88_io_out ? io_r_66_b : _GEN_17965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17967 = 8'h43 == r_count_88_io_out ? io_r_67_b : _GEN_17966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17968 = 8'h44 == r_count_88_io_out ? io_r_68_b : _GEN_17967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17969 = 8'h45 == r_count_88_io_out ? io_r_69_b : _GEN_17968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17970 = 8'h46 == r_count_88_io_out ? io_r_70_b : _GEN_17969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17971 = 8'h47 == r_count_88_io_out ? io_r_71_b : _GEN_17970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17972 = 8'h48 == r_count_88_io_out ? io_r_72_b : _GEN_17971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17973 = 8'h49 == r_count_88_io_out ? io_r_73_b : _GEN_17972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17974 = 8'h4a == r_count_88_io_out ? io_r_74_b : _GEN_17973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17975 = 8'h4b == r_count_88_io_out ? io_r_75_b : _GEN_17974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17976 = 8'h4c == r_count_88_io_out ? io_r_76_b : _GEN_17975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17977 = 8'h4d == r_count_88_io_out ? io_r_77_b : _GEN_17976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17978 = 8'h4e == r_count_88_io_out ? io_r_78_b : _GEN_17977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17979 = 8'h4f == r_count_88_io_out ? io_r_79_b : _GEN_17978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17980 = 8'h50 == r_count_88_io_out ? io_r_80_b : _GEN_17979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17981 = 8'h51 == r_count_88_io_out ? io_r_81_b : _GEN_17980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17982 = 8'h52 == r_count_88_io_out ? io_r_82_b : _GEN_17981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17983 = 8'h53 == r_count_88_io_out ? io_r_83_b : _GEN_17982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17984 = 8'h54 == r_count_88_io_out ? io_r_84_b : _GEN_17983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17985 = 8'h55 == r_count_88_io_out ? io_r_85_b : _GEN_17984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17986 = 8'h56 == r_count_88_io_out ? io_r_86_b : _GEN_17985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17987 = 8'h57 == r_count_88_io_out ? io_r_87_b : _GEN_17986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17988 = 8'h58 == r_count_88_io_out ? io_r_88_b : _GEN_17987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17989 = 8'h59 == r_count_88_io_out ? io_r_89_b : _GEN_17988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17990 = 8'h5a == r_count_88_io_out ? io_r_90_b : _GEN_17989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17991 = 8'h5b == r_count_88_io_out ? io_r_91_b : _GEN_17990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17992 = 8'h5c == r_count_88_io_out ? io_r_92_b : _GEN_17991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17993 = 8'h5d == r_count_88_io_out ? io_r_93_b : _GEN_17992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17994 = 8'h5e == r_count_88_io_out ? io_r_94_b : _GEN_17993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17995 = 8'h5f == r_count_88_io_out ? io_r_95_b : _GEN_17994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17996 = 8'h60 == r_count_88_io_out ? io_r_96_b : _GEN_17995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17997 = 8'h61 == r_count_88_io_out ? io_r_97_b : _GEN_17996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17998 = 8'h62 == r_count_88_io_out ? io_r_98_b : _GEN_17997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_17999 = 8'h63 == r_count_88_io_out ? io_r_99_b : _GEN_17998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18000 = 8'h64 == r_count_88_io_out ? io_r_100_b : _GEN_17999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18001 = 8'h65 == r_count_88_io_out ? io_r_101_b : _GEN_18000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18002 = 8'h66 == r_count_88_io_out ? io_r_102_b : _GEN_18001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18003 = 8'h67 == r_count_88_io_out ? io_r_103_b : _GEN_18002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18004 = 8'h68 == r_count_88_io_out ? io_r_104_b : _GEN_18003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18005 = 8'h69 == r_count_88_io_out ? io_r_105_b : _GEN_18004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18006 = 8'h6a == r_count_88_io_out ? io_r_106_b : _GEN_18005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18007 = 8'h6b == r_count_88_io_out ? io_r_107_b : _GEN_18006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18008 = 8'h6c == r_count_88_io_out ? io_r_108_b : _GEN_18007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18009 = 8'h6d == r_count_88_io_out ? io_r_109_b : _GEN_18008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18010 = 8'h6e == r_count_88_io_out ? io_r_110_b : _GEN_18009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18011 = 8'h6f == r_count_88_io_out ? io_r_111_b : _GEN_18010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18012 = 8'h70 == r_count_88_io_out ? io_r_112_b : _GEN_18011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18013 = 8'h71 == r_count_88_io_out ? io_r_113_b : _GEN_18012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18014 = 8'h72 == r_count_88_io_out ? io_r_114_b : _GEN_18013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18015 = 8'h73 == r_count_88_io_out ? io_r_115_b : _GEN_18014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18016 = 8'h74 == r_count_88_io_out ? io_r_116_b : _GEN_18015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18017 = 8'h75 == r_count_88_io_out ? io_r_117_b : _GEN_18016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18018 = 8'h76 == r_count_88_io_out ? io_r_118_b : _GEN_18017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18019 = 8'h77 == r_count_88_io_out ? io_r_119_b : _GEN_18018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18020 = 8'h78 == r_count_88_io_out ? io_r_120_b : _GEN_18019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18021 = 8'h79 == r_count_88_io_out ? io_r_121_b : _GEN_18020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18022 = 8'h7a == r_count_88_io_out ? io_r_122_b : _GEN_18021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18023 = 8'h7b == r_count_88_io_out ? io_r_123_b : _GEN_18022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18024 = 8'h7c == r_count_88_io_out ? io_r_124_b : _GEN_18023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18025 = 8'h7d == r_count_88_io_out ? io_r_125_b : _GEN_18024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18026 = 8'h7e == r_count_88_io_out ? io_r_126_b : _GEN_18025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18027 = 8'h7f == r_count_88_io_out ? io_r_127_b : _GEN_18026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18028 = 8'h80 == r_count_88_io_out ? io_r_128_b : _GEN_18027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18029 = 8'h81 == r_count_88_io_out ? io_r_129_b : _GEN_18028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18030 = 8'h82 == r_count_88_io_out ? io_r_130_b : _GEN_18029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18031 = 8'h83 == r_count_88_io_out ? io_r_131_b : _GEN_18030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18032 = 8'h84 == r_count_88_io_out ? io_r_132_b : _GEN_18031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18033 = 8'h85 == r_count_88_io_out ? io_r_133_b : _GEN_18032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18034 = 8'h86 == r_count_88_io_out ? io_r_134_b : _GEN_18033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18035 = 8'h87 == r_count_88_io_out ? io_r_135_b : _GEN_18034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18036 = 8'h88 == r_count_88_io_out ? io_r_136_b : _GEN_18035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18037 = 8'h89 == r_count_88_io_out ? io_r_137_b : _GEN_18036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18038 = 8'h8a == r_count_88_io_out ? io_r_138_b : _GEN_18037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18039 = 8'h8b == r_count_88_io_out ? io_r_139_b : _GEN_18038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18040 = 8'h8c == r_count_88_io_out ? io_r_140_b : _GEN_18039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18041 = 8'h8d == r_count_88_io_out ? io_r_141_b : _GEN_18040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18042 = 8'h8e == r_count_88_io_out ? io_r_142_b : _GEN_18041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18043 = 8'h8f == r_count_88_io_out ? io_r_143_b : _GEN_18042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18044 = 8'h90 == r_count_88_io_out ? io_r_144_b : _GEN_18043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18045 = 8'h91 == r_count_88_io_out ? io_r_145_b : _GEN_18044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18046 = 8'h92 == r_count_88_io_out ? io_r_146_b : _GEN_18045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18047 = 8'h93 == r_count_88_io_out ? io_r_147_b : _GEN_18046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18048 = 8'h94 == r_count_88_io_out ? io_r_148_b : _GEN_18047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18049 = 8'h95 == r_count_88_io_out ? io_r_149_b : _GEN_18048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18050 = 8'h96 == r_count_88_io_out ? io_r_150_b : _GEN_18049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18051 = 8'h97 == r_count_88_io_out ? io_r_151_b : _GEN_18050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18052 = 8'h98 == r_count_88_io_out ? io_r_152_b : _GEN_18051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18053 = 8'h99 == r_count_88_io_out ? io_r_153_b : _GEN_18052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18054 = 8'h9a == r_count_88_io_out ? io_r_154_b : _GEN_18053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18055 = 8'h9b == r_count_88_io_out ? io_r_155_b : _GEN_18054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18056 = 8'h9c == r_count_88_io_out ? io_r_156_b : _GEN_18055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18057 = 8'h9d == r_count_88_io_out ? io_r_157_b : _GEN_18056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18058 = 8'h9e == r_count_88_io_out ? io_r_158_b : _GEN_18057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18059 = 8'h9f == r_count_88_io_out ? io_r_159_b : _GEN_18058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18060 = 8'ha0 == r_count_88_io_out ? io_r_160_b : _GEN_18059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18061 = 8'ha1 == r_count_88_io_out ? io_r_161_b : _GEN_18060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18062 = 8'ha2 == r_count_88_io_out ? io_r_162_b : _GEN_18061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18063 = 8'ha3 == r_count_88_io_out ? io_r_163_b : _GEN_18062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18064 = 8'ha4 == r_count_88_io_out ? io_r_164_b : _GEN_18063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18065 = 8'ha5 == r_count_88_io_out ? io_r_165_b : _GEN_18064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18066 = 8'ha6 == r_count_88_io_out ? io_r_166_b : _GEN_18065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18067 = 8'ha7 == r_count_88_io_out ? io_r_167_b : _GEN_18066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18068 = 8'ha8 == r_count_88_io_out ? io_r_168_b : _GEN_18067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18069 = 8'ha9 == r_count_88_io_out ? io_r_169_b : _GEN_18068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18070 = 8'haa == r_count_88_io_out ? io_r_170_b : _GEN_18069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18071 = 8'hab == r_count_88_io_out ? io_r_171_b : _GEN_18070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18072 = 8'hac == r_count_88_io_out ? io_r_172_b : _GEN_18071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18073 = 8'had == r_count_88_io_out ? io_r_173_b : _GEN_18072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18074 = 8'hae == r_count_88_io_out ? io_r_174_b : _GEN_18073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18075 = 8'haf == r_count_88_io_out ? io_r_175_b : _GEN_18074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18076 = 8'hb0 == r_count_88_io_out ? io_r_176_b : _GEN_18075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18077 = 8'hb1 == r_count_88_io_out ? io_r_177_b : _GEN_18076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18078 = 8'hb2 == r_count_88_io_out ? io_r_178_b : _GEN_18077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18079 = 8'hb3 == r_count_88_io_out ? io_r_179_b : _GEN_18078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18080 = 8'hb4 == r_count_88_io_out ? io_r_180_b : _GEN_18079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18081 = 8'hb5 == r_count_88_io_out ? io_r_181_b : _GEN_18080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18082 = 8'hb6 == r_count_88_io_out ? io_r_182_b : _GEN_18081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18083 = 8'hb7 == r_count_88_io_out ? io_r_183_b : _GEN_18082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18084 = 8'hb8 == r_count_88_io_out ? io_r_184_b : _GEN_18083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18085 = 8'hb9 == r_count_88_io_out ? io_r_185_b : _GEN_18084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18086 = 8'hba == r_count_88_io_out ? io_r_186_b : _GEN_18085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18087 = 8'hbb == r_count_88_io_out ? io_r_187_b : _GEN_18086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18088 = 8'hbc == r_count_88_io_out ? io_r_188_b : _GEN_18087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18089 = 8'hbd == r_count_88_io_out ? io_r_189_b : _GEN_18088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18090 = 8'hbe == r_count_88_io_out ? io_r_190_b : _GEN_18089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18091 = 8'hbf == r_count_88_io_out ? io_r_191_b : _GEN_18090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18092 = 8'hc0 == r_count_88_io_out ? io_r_192_b : _GEN_18091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18093 = 8'hc1 == r_count_88_io_out ? io_r_193_b : _GEN_18092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18094 = 8'hc2 == r_count_88_io_out ? io_r_194_b : _GEN_18093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18095 = 8'hc3 == r_count_88_io_out ? io_r_195_b : _GEN_18094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18096 = 8'hc4 == r_count_88_io_out ? io_r_196_b : _GEN_18095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18097 = 8'hc5 == r_count_88_io_out ? io_r_197_b : _GEN_18096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18098 = 8'hc6 == r_count_88_io_out ? io_r_198_b : _GEN_18097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18101 = 8'h1 == r_count_89_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18102 = 8'h2 == r_count_89_io_out ? io_r_2_b : _GEN_18101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18103 = 8'h3 == r_count_89_io_out ? io_r_3_b : _GEN_18102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18104 = 8'h4 == r_count_89_io_out ? io_r_4_b : _GEN_18103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18105 = 8'h5 == r_count_89_io_out ? io_r_5_b : _GEN_18104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18106 = 8'h6 == r_count_89_io_out ? io_r_6_b : _GEN_18105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18107 = 8'h7 == r_count_89_io_out ? io_r_7_b : _GEN_18106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18108 = 8'h8 == r_count_89_io_out ? io_r_8_b : _GEN_18107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18109 = 8'h9 == r_count_89_io_out ? io_r_9_b : _GEN_18108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18110 = 8'ha == r_count_89_io_out ? io_r_10_b : _GEN_18109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18111 = 8'hb == r_count_89_io_out ? io_r_11_b : _GEN_18110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18112 = 8'hc == r_count_89_io_out ? io_r_12_b : _GEN_18111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18113 = 8'hd == r_count_89_io_out ? io_r_13_b : _GEN_18112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18114 = 8'he == r_count_89_io_out ? io_r_14_b : _GEN_18113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18115 = 8'hf == r_count_89_io_out ? io_r_15_b : _GEN_18114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18116 = 8'h10 == r_count_89_io_out ? io_r_16_b : _GEN_18115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18117 = 8'h11 == r_count_89_io_out ? io_r_17_b : _GEN_18116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18118 = 8'h12 == r_count_89_io_out ? io_r_18_b : _GEN_18117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18119 = 8'h13 == r_count_89_io_out ? io_r_19_b : _GEN_18118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18120 = 8'h14 == r_count_89_io_out ? io_r_20_b : _GEN_18119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18121 = 8'h15 == r_count_89_io_out ? io_r_21_b : _GEN_18120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18122 = 8'h16 == r_count_89_io_out ? io_r_22_b : _GEN_18121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18123 = 8'h17 == r_count_89_io_out ? io_r_23_b : _GEN_18122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18124 = 8'h18 == r_count_89_io_out ? io_r_24_b : _GEN_18123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18125 = 8'h19 == r_count_89_io_out ? io_r_25_b : _GEN_18124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18126 = 8'h1a == r_count_89_io_out ? io_r_26_b : _GEN_18125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18127 = 8'h1b == r_count_89_io_out ? io_r_27_b : _GEN_18126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18128 = 8'h1c == r_count_89_io_out ? io_r_28_b : _GEN_18127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18129 = 8'h1d == r_count_89_io_out ? io_r_29_b : _GEN_18128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18130 = 8'h1e == r_count_89_io_out ? io_r_30_b : _GEN_18129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18131 = 8'h1f == r_count_89_io_out ? io_r_31_b : _GEN_18130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18132 = 8'h20 == r_count_89_io_out ? io_r_32_b : _GEN_18131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18133 = 8'h21 == r_count_89_io_out ? io_r_33_b : _GEN_18132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18134 = 8'h22 == r_count_89_io_out ? io_r_34_b : _GEN_18133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18135 = 8'h23 == r_count_89_io_out ? io_r_35_b : _GEN_18134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18136 = 8'h24 == r_count_89_io_out ? io_r_36_b : _GEN_18135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18137 = 8'h25 == r_count_89_io_out ? io_r_37_b : _GEN_18136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18138 = 8'h26 == r_count_89_io_out ? io_r_38_b : _GEN_18137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18139 = 8'h27 == r_count_89_io_out ? io_r_39_b : _GEN_18138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18140 = 8'h28 == r_count_89_io_out ? io_r_40_b : _GEN_18139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18141 = 8'h29 == r_count_89_io_out ? io_r_41_b : _GEN_18140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18142 = 8'h2a == r_count_89_io_out ? io_r_42_b : _GEN_18141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18143 = 8'h2b == r_count_89_io_out ? io_r_43_b : _GEN_18142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18144 = 8'h2c == r_count_89_io_out ? io_r_44_b : _GEN_18143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18145 = 8'h2d == r_count_89_io_out ? io_r_45_b : _GEN_18144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18146 = 8'h2e == r_count_89_io_out ? io_r_46_b : _GEN_18145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18147 = 8'h2f == r_count_89_io_out ? io_r_47_b : _GEN_18146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18148 = 8'h30 == r_count_89_io_out ? io_r_48_b : _GEN_18147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18149 = 8'h31 == r_count_89_io_out ? io_r_49_b : _GEN_18148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18150 = 8'h32 == r_count_89_io_out ? io_r_50_b : _GEN_18149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18151 = 8'h33 == r_count_89_io_out ? io_r_51_b : _GEN_18150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18152 = 8'h34 == r_count_89_io_out ? io_r_52_b : _GEN_18151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18153 = 8'h35 == r_count_89_io_out ? io_r_53_b : _GEN_18152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18154 = 8'h36 == r_count_89_io_out ? io_r_54_b : _GEN_18153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18155 = 8'h37 == r_count_89_io_out ? io_r_55_b : _GEN_18154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18156 = 8'h38 == r_count_89_io_out ? io_r_56_b : _GEN_18155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18157 = 8'h39 == r_count_89_io_out ? io_r_57_b : _GEN_18156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18158 = 8'h3a == r_count_89_io_out ? io_r_58_b : _GEN_18157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18159 = 8'h3b == r_count_89_io_out ? io_r_59_b : _GEN_18158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18160 = 8'h3c == r_count_89_io_out ? io_r_60_b : _GEN_18159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18161 = 8'h3d == r_count_89_io_out ? io_r_61_b : _GEN_18160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18162 = 8'h3e == r_count_89_io_out ? io_r_62_b : _GEN_18161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18163 = 8'h3f == r_count_89_io_out ? io_r_63_b : _GEN_18162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18164 = 8'h40 == r_count_89_io_out ? io_r_64_b : _GEN_18163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18165 = 8'h41 == r_count_89_io_out ? io_r_65_b : _GEN_18164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18166 = 8'h42 == r_count_89_io_out ? io_r_66_b : _GEN_18165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18167 = 8'h43 == r_count_89_io_out ? io_r_67_b : _GEN_18166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18168 = 8'h44 == r_count_89_io_out ? io_r_68_b : _GEN_18167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18169 = 8'h45 == r_count_89_io_out ? io_r_69_b : _GEN_18168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18170 = 8'h46 == r_count_89_io_out ? io_r_70_b : _GEN_18169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18171 = 8'h47 == r_count_89_io_out ? io_r_71_b : _GEN_18170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18172 = 8'h48 == r_count_89_io_out ? io_r_72_b : _GEN_18171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18173 = 8'h49 == r_count_89_io_out ? io_r_73_b : _GEN_18172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18174 = 8'h4a == r_count_89_io_out ? io_r_74_b : _GEN_18173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18175 = 8'h4b == r_count_89_io_out ? io_r_75_b : _GEN_18174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18176 = 8'h4c == r_count_89_io_out ? io_r_76_b : _GEN_18175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18177 = 8'h4d == r_count_89_io_out ? io_r_77_b : _GEN_18176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18178 = 8'h4e == r_count_89_io_out ? io_r_78_b : _GEN_18177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18179 = 8'h4f == r_count_89_io_out ? io_r_79_b : _GEN_18178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18180 = 8'h50 == r_count_89_io_out ? io_r_80_b : _GEN_18179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18181 = 8'h51 == r_count_89_io_out ? io_r_81_b : _GEN_18180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18182 = 8'h52 == r_count_89_io_out ? io_r_82_b : _GEN_18181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18183 = 8'h53 == r_count_89_io_out ? io_r_83_b : _GEN_18182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18184 = 8'h54 == r_count_89_io_out ? io_r_84_b : _GEN_18183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18185 = 8'h55 == r_count_89_io_out ? io_r_85_b : _GEN_18184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18186 = 8'h56 == r_count_89_io_out ? io_r_86_b : _GEN_18185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18187 = 8'h57 == r_count_89_io_out ? io_r_87_b : _GEN_18186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18188 = 8'h58 == r_count_89_io_out ? io_r_88_b : _GEN_18187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18189 = 8'h59 == r_count_89_io_out ? io_r_89_b : _GEN_18188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18190 = 8'h5a == r_count_89_io_out ? io_r_90_b : _GEN_18189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18191 = 8'h5b == r_count_89_io_out ? io_r_91_b : _GEN_18190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18192 = 8'h5c == r_count_89_io_out ? io_r_92_b : _GEN_18191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18193 = 8'h5d == r_count_89_io_out ? io_r_93_b : _GEN_18192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18194 = 8'h5e == r_count_89_io_out ? io_r_94_b : _GEN_18193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18195 = 8'h5f == r_count_89_io_out ? io_r_95_b : _GEN_18194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18196 = 8'h60 == r_count_89_io_out ? io_r_96_b : _GEN_18195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18197 = 8'h61 == r_count_89_io_out ? io_r_97_b : _GEN_18196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18198 = 8'h62 == r_count_89_io_out ? io_r_98_b : _GEN_18197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18199 = 8'h63 == r_count_89_io_out ? io_r_99_b : _GEN_18198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18200 = 8'h64 == r_count_89_io_out ? io_r_100_b : _GEN_18199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18201 = 8'h65 == r_count_89_io_out ? io_r_101_b : _GEN_18200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18202 = 8'h66 == r_count_89_io_out ? io_r_102_b : _GEN_18201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18203 = 8'h67 == r_count_89_io_out ? io_r_103_b : _GEN_18202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18204 = 8'h68 == r_count_89_io_out ? io_r_104_b : _GEN_18203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18205 = 8'h69 == r_count_89_io_out ? io_r_105_b : _GEN_18204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18206 = 8'h6a == r_count_89_io_out ? io_r_106_b : _GEN_18205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18207 = 8'h6b == r_count_89_io_out ? io_r_107_b : _GEN_18206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18208 = 8'h6c == r_count_89_io_out ? io_r_108_b : _GEN_18207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18209 = 8'h6d == r_count_89_io_out ? io_r_109_b : _GEN_18208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18210 = 8'h6e == r_count_89_io_out ? io_r_110_b : _GEN_18209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18211 = 8'h6f == r_count_89_io_out ? io_r_111_b : _GEN_18210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18212 = 8'h70 == r_count_89_io_out ? io_r_112_b : _GEN_18211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18213 = 8'h71 == r_count_89_io_out ? io_r_113_b : _GEN_18212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18214 = 8'h72 == r_count_89_io_out ? io_r_114_b : _GEN_18213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18215 = 8'h73 == r_count_89_io_out ? io_r_115_b : _GEN_18214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18216 = 8'h74 == r_count_89_io_out ? io_r_116_b : _GEN_18215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18217 = 8'h75 == r_count_89_io_out ? io_r_117_b : _GEN_18216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18218 = 8'h76 == r_count_89_io_out ? io_r_118_b : _GEN_18217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18219 = 8'h77 == r_count_89_io_out ? io_r_119_b : _GEN_18218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18220 = 8'h78 == r_count_89_io_out ? io_r_120_b : _GEN_18219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18221 = 8'h79 == r_count_89_io_out ? io_r_121_b : _GEN_18220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18222 = 8'h7a == r_count_89_io_out ? io_r_122_b : _GEN_18221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18223 = 8'h7b == r_count_89_io_out ? io_r_123_b : _GEN_18222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18224 = 8'h7c == r_count_89_io_out ? io_r_124_b : _GEN_18223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18225 = 8'h7d == r_count_89_io_out ? io_r_125_b : _GEN_18224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18226 = 8'h7e == r_count_89_io_out ? io_r_126_b : _GEN_18225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18227 = 8'h7f == r_count_89_io_out ? io_r_127_b : _GEN_18226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18228 = 8'h80 == r_count_89_io_out ? io_r_128_b : _GEN_18227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18229 = 8'h81 == r_count_89_io_out ? io_r_129_b : _GEN_18228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18230 = 8'h82 == r_count_89_io_out ? io_r_130_b : _GEN_18229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18231 = 8'h83 == r_count_89_io_out ? io_r_131_b : _GEN_18230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18232 = 8'h84 == r_count_89_io_out ? io_r_132_b : _GEN_18231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18233 = 8'h85 == r_count_89_io_out ? io_r_133_b : _GEN_18232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18234 = 8'h86 == r_count_89_io_out ? io_r_134_b : _GEN_18233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18235 = 8'h87 == r_count_89_io_out ? io_r_135_b : _GEN_18234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18236 = 8'h88 == r_count_89_io_out ? io_r_136_b : _GEN_18235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18237 = 8'h89 == r_count_89_io_out ? io_r_137_b : _GEN_18236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18238 = 8'h8a == r_count_89_io_out ? io_r_138_b : _GEN_18237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18239 = 8'h8b == r_count_89_io_out ? io_r_139_b : _GEN_18238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18240 = 8'h8c == r_count_89_io_out ? io_r_140_b : _GEN_18239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18241 = 8'h8d == r_count_89_io_out ? io_r_141_b : _GEN_18240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18242 = 8'h8e == r_count_89_io_out ? io_r_142_b : _GEN_18241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18243 = 8'h8f == r_count_89_io_out ? io_r_143_b : _GEN_18242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18244 = 8'h90 == r_count_89_io_out ? io_r_144_b : _GEN_18243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18245 = 8'h91 == r_count_89_io_out ? io_r_145_b : _GEN_18244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18246 = 8'h92 == r_count_89_io_out ? io_r_146_b : _GEN_18245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18247 = 8'h93 == r_count_89_io_out ? io_r_147_b : _GEN_18246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18248 = 8'h94 == r_count_89_io_out ? io_r_148_b : _GEN_18247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18249 = 8'h95 == r_count_89_io_out ? io_r_149_b : _GEN_18248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18250 = 8'h96 == r_count_89_io_out ? io_r_150_b : _GEN_18249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18251 = 8'h97 == r_count_89_io_out ? io_r_151_b : _GEN_18250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18252 = 8'h98 == r_count_89_io_out ? io_r_152_b : _GEN_18251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18253 = 8'h99 == r_count_89_io_out ? io_r_153_b : _GEN_18252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18254 = 8'h9a == r_count_89_io_out ? io_r_154_b : _GEN_18253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18255 = 8'h9b == r_count_89_io_out ? io_r_155_b : _GEN_18254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18256 = 8'h9c == r_count_89_io_out ? io_r_156_b : _GEN_18255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18257 = 8'h9d == r_count_89_io_out ? io_r_157_b : _GEN_18256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18258 = 8'h9e == r_count_89_io_out ? io_r_158_b : _GEN_18257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18259 = 8'h9f == r_count_89_io_out ? io_r_159_b : _GEN_18258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18260 = 8'ha0 == r_count_89_io_out ? io_r_160_b : _GEN_18259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18261 = 8'ha1 == r_count_89_io_out ? io_r_161_b : _GEN_18260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18262 = 8'ha2 == r_count_89_io_out ? io_r_162_b : _GEN_18261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18263 = 8'ha3 == r_count_89_io_out ? io_r_163_b : _GEN_18262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18264 = 8'ha4 == r_count_89_io_out ? io_r_164_b : _GEN_18263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18265 = 8'ha5 == r_count_89_io_out ? io_r_165_b : _GEN_18264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18266 = 8'ha6 == r_count_89_io_out ? io_r_166_b : _GEN_18265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18267 = 8'ha7 == r_count_89_io_out ? io_r_167_b : _GEN_18266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18268 = 8'ha8 == r_count_89_io_out ? io_r_168_b : _GEN_18267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18269 = 8'ha9 == r_count_89_io_out ? io_r_169_b : _GEN_18268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18270 = 8'haa == r_count_89_io_out ? io_r_170_b : _GEN_18269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18271 = 8'hab == r_count_89_io_out ? io_r_171_b : _GEN_18270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18272 = 8'hac == r_count_89_io_out ? io_r_172_b : _GEN_18271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18273 = 8'had == r_count_89_io_out ? io_r_173_b : _GEN_18272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18274 = 8'hae == r_count_89_io_out ? io_r_174_b : _GEN_18273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18275 = 8'haf == r_count_89_io_out ? io_r_175_b : _GEN_18274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18276 = 8'hb0 == r_count_89_io_out ? io_r_176_b : _GEN_18275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18277 = 8'hb1 == r_count_89_io_out ? io_r_177_b : _GEN_18276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18278 = 8'hb2 == r_count_89_io_out ? io_r_178_b : _GEN_18277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18279 = 8'hb3 == r_count_89_io_out ? io_r_179_b : _GEN_18278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18280 = 8'hb4 == r_count_89_io_out ? io_r_180_b : _GEN_18279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18281 = 8'hb5 == r_count_89_io_out ? io_r_181_b : _GEN_18280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18282 = 8'hb6 == r_count_89_io_out ? io_r_182_b : _GEN_18281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18283 = 8'hb7 == r_count_89_io_out ? io_r_183_b : _GEN_18282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18284 = 8'hb8 == r_count_89_io_out ? io_r_184_b : _GEN_18283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18285 = 8'hb9 == r_count_89_io_out ? io_r_185_b : _GEN_18284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18286 = 8'hba == r_count_89_io_out ? io_r_186_b : _GEN_18285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18287 = 8'hbb == r_count_89_io_out ? io_r_187_b : _GEN_18286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18288 = 8'hbc == r_count_89_io_out ? io_r_188_b : _GEN_18287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18289 = 8'hbd == r_count_89_io_out ? io_r_189_b : _GEN_18288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18290 = 8'hbe == r_count_89_io_out ? io_r_190_b : _GEN_18289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18291 = 8'hbf == r_count_89_io_out ? io_r_191_b : _GEN_18290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18292 = 8'hc0 == r_count_89_io_out ? io_r_192_b : _GEN_18291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18293 = 8'hc1 == r_count_89_io_out ? io_r_193_b : _GEN_18292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18294 = 8'hc2 == r_count_89_io_out ? io_r_194_b : _GEN_18293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18295 = 8'hc3 == r_count_89_io_out ? io_r_195_b : _GEN_18294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18296 = 8'hc4 == r_count_89_io_out ? io_r_196_b : _GEN_18295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18297 = 8'hc5 == r_count_89_io_out ? io_r_197_b : _GEN_18296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18298 = 8'hc6 == r_count_89_io_out ? io_r_198_b : _GEN_18297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18301 = 8'h1 == r_count_90_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18302 = 8'h2 == r_count_90_io_out ? io_r_2_b : _GEN_18301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18303 = 8'h3 == r_count_90_io_out ? io_r_3_b : _GEN_18302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18304 = 8'h4 == r_count_90_io_out ? io_r_4_b : _GEN_18303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18305 = 8'h5 == r_count_90_io_out ? io_r_5_b : _GEN_18304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18306 = 8'h6 == r_count_90_io_out ? io_r_6_b : _GEN_18305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18307 = 8'h7 == r_count_90_io_out ? io_r_7_b : _GEN_18306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18308 = 8'h8 == r_count_90_io_out ? io_r_8_b : _GEN_18307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18309 = 8'h9 == r_count_90_io_out ? io_r_9_b : _GEN_18308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18310 = 8'ha == r_count_90_io_out ? io_r_10_b : _GEN_18309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18311 = 8'hb == r_count_90_io_out ? io_r_11_b : _GEN_18310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18312 = 8'hc == r_count_90_io_out ? io_r_12_b : _GEN_18311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18313 = 8'hd == r_count_90_io_out ? io_r_13_b : _GEN_18312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18314 = 8'he == r_count_90_io_out ? io_r_14_b : _GEN_18313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18315 = 8'hf == r_count_90_io_out ? io_r_15_b : _GEN_18314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18316 = 8'h10 == r_count_90_io_out ? io_r_16_b : _GEN_18315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18317 = 8'h11 == r_count_90_io_out ? io_r_17_b : _GEN_18316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18318 = 8'h12 == r_count_90_io_out ? io_r_18_b : _GEN_18317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18319 = 8'h13 == r_count_90_io_out ? io_r_19_b : _GEN_18318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18320 = 8'h14 == r_count_90_io_out ? io_r_20_b : _GEN_18319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18321 = 8'h15 == r_count_90_io_out ? io_r_21_b : _GEN_18320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18322 = 8'h16 == r_count_90_io_out ? io_r_22_b : _GEN_18321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18323 = 8'h17 == r_count_90_io_out ? io_r_23_b : _GEN_18322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18324 = 8'h18 == r_count_90_io_out ? io_r_24_b : _GEN_18323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18325 = 8'h19 == r_count_90_io_out ? io_r_25_b : _GEN_18324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18326 = 8'h1a == r_count_90_io_out ? io_r_26_b : _GEN_18325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18327 = 8'h1b == r_count_90_io_out ? io_r_27_b : _GEN_18326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18328 = 8'h1c == r_count_90_io_out ? io_r_28_b : _GEN_18327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18329 = 8'h1d == r_count_90_io_out ? io_r_29_b : _GEN_18328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18330 = 8'h1e == r_count_90_io_out ? io_r_30_b : _GEN_18329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18331 = 8'h1f == r_count_90_io_out ? io_r_31_b : _GEN_18330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18332 = 8'h20 == r_count_90_io_out ? io_r_32_b : _GEN_18331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18333 = 8'h21 == r_count_90_io_out ? io_r_33_b : _GEN_18332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18334 = 8'h22 == r_count_90_io_out ? io_r_34_b : _GEN_18333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18335 = 8'h23 == r_count_90_io_out ? io_r_35_b : _GEN_18334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18336 = 8'h24 == r_count_90_io_out ? io_r_36_b : _GEN_18335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18337 = 8'h25 == r_count_90_io_out ? io_r_37_b : _GEN_18336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18338 = 8'h26 == r_count_90_io_out ? io_r_38_b : _GEN_18337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18339 = 8'h27 == r_count_90_io_out ? io_r_39_b : _GEN_18338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18340 = 8'h28 == r_count_90_io_out ? io_r_40_b : _GEN_18339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18341 = 8'h29 == r_count_90_io_out ? io_r_41_b : _GEN_18340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18342 = 8'h2a == r_count_90_io_out ? io_r_42_b : _GEN_18341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18343 = 8'h2b == r_count_90_io_out ? io_r_43_b : _GEN_18342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18344 = 8'h2c == r_count_90_io_out ? io_r_44_b : _GEN_18343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18345 = 8'h2d == r_count_90_io_out ? io_r_45_b : _GEN_18344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18346 = 8'h2e == r_count_90_io_out ? io_r_46_b : _GEN_18345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18347 = 8'h2f == r_count_90_io_out ? io_r_47_b : _GEN_18346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18348 = 8'h30 == r_count_90_io_out ? io_r_48_b : _GEN_18347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18349 = 8'h31 == r_count_90_io_out ? io_r_49_b : _GEN_18348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18350 = 8'h32 == r_count_90_io_out ? io_r_50_b : _GEN_18349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18351 = 8'h33 == r_count_90_io_out ? io_r_51_b : _GEN_18350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18352 = 8'h34 == r_count_90_io_out ? io_r_52_b : _GEN_18351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18353 = 8'h35 == r_count_90_io_out ? io_r_53_b : _GEN_18352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18354 = 8'h36 == r_count_90_io_out ? io_r_54_b : _GEN_18353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18355 = 8'h37 == r_count_90_io_out ? io_r_55_b : _GEN_18354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18356 = 8'h38 == r_count_90_io_out ? io_r_56_b : _GEN_18355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18357 = 8'h39 == r_count_90_io_out ? io_r_57_b : _GEN_18356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18358 = 8'h3a == r_count_90_io_out ? io_r_58_b : _GEN_18357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18359 = 8'h3b == r_count_90_io_out ? io_r_59_b : _GEN_18358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18360 = 8'h3c == r_count_90_io_out ? io_r_60_b : _GEN_18359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18361 = 8'h3d == r_count_90_io_out ? io_r_61_b : _GEN_18360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18362 = 8'h3e == r_count_90_io_out ? io_r_62_b : _GEN_18361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18363 = 8'h3f == r_count_90_io_out ? io_r_63_b : _GEN_18362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18364 = 8'h40 == r_count_90_io_out ? io_r_64_b : _GEN_18363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18365 = 8'h41 == r_count_90_io_out ? io_r_65_b : _GEN_18364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18366 = 8'h42 == r_count_90_io_out ? io_r_66_b : _GEN_18365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18367 = 8'h43 == r_count_90_io_out ? io_r_67_b : _GEN_18366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18368 = 8'h44 == r_count_90_io_out ? io_r_68_b : _GEN_18367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18369 = 8'h45 == r_count_90_io_out ? io_r_69_b : _GEN_18368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18370 = 8'h46 == r_count_90_io_out ? io_r_70_b : _GEN_18369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18371 = 8'h47 == r_count_90_io_out ? io_r_71_b : _GEN_18370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18372 = 8'h48 == r_count_90_io_out ? io_r_72_b : _GEN_18371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18373 = 8'h49 == r_count_90_io_out ? io_r_73_b : _GEN_18372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18374 = 8'h4a == r_count_90_io_out ? io_r_74_b : _GEN_18373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18375 = 8'h4b == r_count_90_io_out ? io_r_75_b : _GEN_18374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18376 = 8'h4c == r_count_90_io_out ? io_r_76_b : _GEN_18375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18377 = 8'h4d == r_count_90_io_out ? io_r_77_b : _GEN_18376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18378 = 8'h4e == r_count_90_io_out ? io_r_78_b : _GEN_18377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18379 = 8'h4f == r_count_90_io_out ? io_r_79_b : _GEN_18378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18380 = 8'h50 == r_count_90_io_out ? io_r_80_b : _GEN_18379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18381 = 8'h51 == r_count_90_io_out ? io_r_81_b : _GEN_18380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18382 = 8'h52 == r_count_90_io_out ? io_r_82_b : _GEN_18381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18383 = 8'h53 == r_count_90_io_out ? io_r_83_b : _GEN_18382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18384 = 8'h54 == r_count_90_io_out ? io_r_84_b : _GEN_18383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18385 = 8'h55 == r_count_90_io_out ? io_r_85_b : _GEN_18384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18386 = 8'h56 == r_count_90_io_out ? io_r_86_b : _GEN_18385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18387 = 8'h57 == r_count_90_io_out ? io_r_87_b : _GEN_18386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18388 = 8'h58 == r_count_90_io_out ? io_r_88_b : _GEN_18387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18389 = 8'h59 == r_count_90_io_out ? io_r_89_b : _GEN_18388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18390 = 8'h5a == r_count_90_io_out ? io_r_90_b : _GEN_18389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18391 = 8'h5b == r_count_90_io_out ? io_r_91_b : _GEN_18390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18392 = 8'h5c == r_count_90_io_out ? io_r_92_b : _GEN_18391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18393 = 8'h5d == r_count_90_io_out ? io_r_93_b : _GEN_18392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18394 = 8'h5e == r_count_90_io_out ? io_r_94_b : _GEN_18393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18395 = 8'h5f == r_count_90_io_out ? io_r_95_b : _GEN_18394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18396 = 8'h60 == r_count_90_io_out ? io_r_96_b : _GEN_18395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18397 = 8'h61 == r_count_90_io_out ? io_r_97_b : _GEN_18396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18398 = 8'h62 == r_count_90_io_out ? io_r_98_b : _GEN_18397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18399 = 8'h63 == r_count_90_io_out ? io_r_99_b : _GEN_18398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18400 = 8'h64 == r_count_90_io_out ? io_r_100_b : _GEN_18399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18401 = 8'h65 == r_count_90_io_out ? io_r_101_b : _GEN_18400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18402 = 8'h66 == r_count_90_io_out ? io_r_102_b : _GEN_18401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18403 = 8'h67 == r_count_90_io_out ? io_r_103_b : _GEN_18402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18404 = 8'h68 == r_count_90_io_out ? io_r_104_b : _GEN_18403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18405 = 8'h69 == r_count_90_io_out ? io_r_105_b : _GEN_18404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18406 = 8'h6a == r_count_90_io_out ? io_r_106_b : _GEN_18405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18407 = 8'h6b == r_count_90_io_out ? io_r_107_b : _GEN_18406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18408 = 8'h6c == r_count_90_io_out ? io_r_108_b : _GEN_18407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18409 = 8'h6d == r_count_90_io_out ? io_r_109_b : _GEN_18408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18410 = 8'h6e == r_count_90_io_out ? io_r_110_b : _GEN_18409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18411 = 8'h6f == r_count_90_io_out ? io_r_111_b : _GEN_18410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18412 = 8'h70 == r_count_90_io_out ? io_r_112_b : _GEN_18411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18413 = 8'h71 == r_count_90_io_out ? io_r_113_b : _GEN_18412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18414 = 8'h72 == r_count_90_io_out ? io_r_114_b : _GEN_18413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18415 = 8'h73 == r_count_90_io_out ? io_r_115_b : _GEN_18414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18416 = 8'h74 == r_count_90_io_out ? io_r_116_b : _GEN_18415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18417 = 8'h75 == r_count_90_io_out ? io_r_117_b : _GEN_18416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18418 = 8'h76 == r_count_90_io_out ? io_r_118_b : _GEN_18417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18419 = 8'h77 == r_count_90_io_out ? io_r_119_b : _GEN_18418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18420 = 8'h78 == r_count_90_io_out ? io_r_120_b : _GEN_18419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18421 = 8'h79 == r_count_90_io_out ? io_r_121_b : _GEN_18420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18422 = 8'h7a == r_count_90_io_out ? io_r_122_b : _GEN_18421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18423 = 8'h7b == r_count_90_io_out ? io_r_123_b : _GEN_18422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18424 = 8'h7c == r_count_90_io_out ? io_r_124_b : _GEN_18423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18425 = 8'h7d == r_count_90_io_out ? io_r_125_b : _GEN_18424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18426 = 8'h7e == r_count_90_io_out ? io_r_126_b : _GEN_18425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18427 = 8'h7f == r_count_90_io_out ? io_r_127_b : _GEN_18426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18428 = 8'h80 == r_count_90_io_out ? io_r_128_b : _GEN_18427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18429 = 8'h81 == r_count_90_io_out ? io_r_129_b : _GEN_18428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18430 = 8'h82 == r_count_90_io_out ? io_r_130_b : _GEN_18429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18431 = 8'h83 == r_count_90_io_out ? io_r_131_b : _GEN_18430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18432 = 8'h84 == r_count_90_io_out ? io_r_132_b : _GEN_18431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18433 = 8'h85 == r_count_90_io_out ? io_r_133_b : _GEN_18432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18434 = 8'h86 == r_count_90_io_out ? io_r_134_b : _GEN_18433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18435 = 8'h87 == r_count_90_io_out ? io_r_135_b : _GEN_18434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18436 = 8'h88 == r_count_90_io_out ? io_r_136_b : _GEN_18435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18437 = 8'h89 == r_count_90_io_out ? io_r_137_b : _GEN_18436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18438 = 8'h8a == r_count_90_io_out ? io_r_138_b : _GEN_18437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18439 = 8'h8b == r_count_90_io_out ? io_r_139_b : _GEN_18438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18440 = 8'h8c == r_count_90_io_out ? io_r_140_b : _GEN_18439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18441 = 8'h8d == r_count_90_io_out ? io_r_141_b : _GEN_18440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18442 = 8'h8e == r_count_90_io_out ? io_r_142_b : _GEN_18441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18443 = 8'h8f == r_count_90_io_out ? io_r_143_b : _GEN_18442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18444 = 8'h90 == r_count_90_io_out ? io_r_144_b : _GEN_18443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18445 = 8'h91 == r_count_90_io_out ? io_r_145_b : _GEN_18444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18446 = 8'h92 == r_count_90_io_out ? io_r_146_b : _GEN_18445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18447 = 8'h93 == r_count_90_io_out ? io_r_147_b : _GEN_18446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18448 = 8'h94 == r_count_90_io_out ? io_r_148_b : _GEN_18447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18449 = 8'h95 == r_count_90_io_out ? io_r_149_b : _GEN_18448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18450 = 8'h96 == r_count_90_io_out ? io_r_150_b : _GEN_18449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18451 = 8'h97 == r_count_90_io_out ? io_r_151_b : _GEN_18450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18452 = 8'h98 == r_count_90_io_out ? io_r_152_b : _GEN_18451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18453 = 8'h99 == r_count_90_io_out ? io_r_153_b : _GEN_18452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18454 = 8'h9a == r_count_90_io_out ? io_r_154_b : _GEN_18453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18455 = 8'h9b == r_count_90_io_out ? io_r_155_b : _GEN_18454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18456 = 8'h9c == r_count_90_io_out ? io_r_156_b : _GEN_18455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18457 = 8'h9d == r_count_90_io_out ? io_r_157_b : _GEN_18456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18458 = 8'h9e == r_count_90_io_out ? io_r_158_b : _GEN_18457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18459 = 8'h9f == r_count_90_io_out ? io_r_159_b : _GEN_18458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18460 = 8'ha0 == r_count_90_io_out ? io_r_160_b : _GEN_18459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18461 = 8'ha1 == r_count_90_io_out ? io_r_161_b : _GEN_18460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18462 = 8'ha2 == r_count_90_io_out ? io_r_162_b : _GEN_18461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18463 = 8'ha3 == r_count_90_io_out ? io_r_163_b : _GEN_18462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18464 = 8'ha4 == r_count_90_io_out ? io_r_164_b : _GEN_18463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18465 = 8'ha5 == r_count_90_io_out ? io_r_165_b : _GEN_18464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18466 = 8'ha6 == r_count_90_io_out ? io_r_166_b : _GEN_18465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18467 = 8'ha7 == r_count_90_io_out ? io_r_167_b : _GEN_18466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18468 = 8'ha8 == r_count_90_io_out ? io_r_168_b : _GEN_18467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18469 = 8'ha9 == r_count_90_io_out ? io_r_169_b : _GEN_18468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18470 = 8'haa == r_count_90_io_out ? io_r_170_b : _GEN_18469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18471 = 8'hab == r_count_90_io_out ? io_r_171_b : _GEN_18470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18472 = 8'hac == r_count_90_io_out ? io_r_172_b : _GEN_18471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18473 = 8'had == r_count_90_io_out ? io_r_173_b : _GEN_18472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18474 = 8'hae == r_count_90_io_out ? io_r_174_b : _GEN_18473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18475 = 8'haf == r_count_90_io_out ? io_r_175_b : _GEN_18474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18476 = 8'hb0 == r_count_90_io_out ? io_r_176_b : _GEN_18475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18477 = 8'hb1 == r_count_90_io_out ? io_r_177_b : _GEN_18476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18478 = 8'hb2 == r_count_90_io_out ? io_r_178_b : _GEN_18477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18479 = 8'hb3 == r_count_90_io_out ? io_r_179_b : _GEN_18478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18480 = 8'hb4 == r_count_90_io_out ? io_r_180_b : _GEN_18479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18481 = 8'hb5 == r_count_90_io_out ? io_r_181_b : _GEN_18480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18482 = 8'hb6 == r_count_90_io_out ? io_r_182_b : _GEN_18481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18483 = 8'hb7 == r_count_90_io_out ? io_r_183_b : _GEN_18482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18484 = 8'hb8 == r_count_90_io_out ? io_r_184_b : _GEN_18483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18485 = 8'hb9 == r_count_90_io_out ? io_r_185_b : _GEN_18484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18486 = 8'hba == r_count_90_io_out ? io_r_186_b : _GEN_18485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18487 = 8'hbb == r_count_90_io_out ? io_r_187_b : _GEN_18486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18488 = 8'hbc == r_count_90_io_out ? io_r_188_b : _GEN_18487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18489 = 8'hbd == r_count_90_io_out ? io_r_189_b : _GEN_18488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18490 = 8'hbe == r_count_90_io_out ? io_r_190_b : _GEN_18489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18491 = 8'hbf == r_count_90_io_out ? io_r_191_b : _GEN_18490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18492 = 8'hc0 == r_count_90_io_out ? io_r_192_b : _GEN_18491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18493 = 8'hc1 == r_count_90_io_out ? io_r_193_b : _GEN_18492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18494 = 8'hc2 == r_count_90_io_out ? io_r_194_b : _GEN_18493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18495 = 8'hc3 == r_count_90_io_out ? io_r_195_b : _GEN_18494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18496 = 8'hc4 == r_count_90_io_out ? io_r_196_b : _GEN_18495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18497 = 8'hc5 == r_count_90_io_out ? io_r_197_b : _GEN_18496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18498 = 8'hc6 == r_count_90_io_out ? io_r_198_b : _GEN_18497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18501 = 8'h1 == r_count_91_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18502 = 8'h2 == r_count_91_io_out ? io_r_2_b : _GEN_18501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18503 = 8'h3 == r_count_91_io_out ? io_r_3_b : _GEN_18502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18504 = 8'h4 == r_count_91_io_out ? io_r_4_b : _GEN_18503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18505 = 8'h5 == r_count_91_io_out ? io_r_5_b : _GEN_18504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18506 = 8'h6 == r_count_91_io_out ? io_r_6_b : _GEN_18505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18507 = 8'h7 == r_count_91_io_out ? io_r_7_b : _GEN_18506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18508 = 8'h8 == r_count_91_io_out ? io_r_8_b : _GEN_18507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18509 = 8'h9 == r_count_91_io_out ? io_r_9_b : _GEN_18508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18510 = 8'ha == r_count_91_io_out ? io_r_10_b : _GEN_18509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18511 = 8'hb == r_count_91_io_out ? io_r_11_b : _GEN_18510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18512 = 8'hc == r_count_91_io_out ? io_r_12_b : _GEN_18511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18513 = 8'hd == r_count_91_io_out ? io_r_13_b : _GEN_18512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18514 = 8'he == r_count_91_io_out ? io_r_14_b : _GEN_18513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18515 = 8'hf == r_count_91_io_out ? io_r_15_b : _GEN_18514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18516 = 8'h10 == r_count_91_io_out ? io_r_16_b : _GEN_18515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18517 = 8'h11 == r_count_91_io_out ? io_r_17_b : _GEN_18516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18518 = 8'h12 == r_count_91_io_out ? io_r_18_b : _GEN_18517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18519 = 8'h13 == r_count_91_io_out ? io_r_19_b : _GEN_18518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18520 = 8'h14 == r_count_91_io_out ? io_r_20_b : _GEN_18519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18521 = 8'h15 == r_count_91_io_out ? io_r_21_b : _GEN_18520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18522 = 8'h16 == r_count_91_io_out ? io_r_22_b : _GEN_18521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18523 = 8'h17 == r_count_91_io_out ? io_r_23_b : _GEN_18522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18524 = 8'h18 == r_count_91_io_out ? io_r_24_b : _GEN_18523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18525 = 8'h19 == r_count_91_io_out ? io_r_25_b : _GEN_18524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18526 = 8'h1a == r_count_91_io_out ? io_r_26_b : _GEN_18525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18527 = 8'h1b == r_count_91_io_out ? io_r_27_b : _GEN_18526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18528 = 8'h1c == r_count_91_io_out ? io_r_28_b : _GEN_18527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18529 = 8'h1d == r_count_91_io_out ? io_r_29_b : _GEN_18528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18530 = 8'h1e == r_count_91_io_out ? io_r_30_b : _GEN_18529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18531 = 8'h1f == r_count_91_io_out ? io_r_31_b : _GEN_18530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18532 = 8'h20 == r_count_91_io_out ? io_r_32_b : _GEN_18531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18533 = 8'h21 == r_count_91_io_out ? io_r_33_b : _GEN_18532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18534 = 8'h22 == r_count_91_io_out ? io_r_34_b : _GEN_18533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18535 = 8'h23 == r_count_91_io_out ? io_r_35_b : _GEN_18534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18536 = 8'h24 == r_count_91_io_out ? io_r_36_b : _GEN_18535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18537 = 8'h25 == r_count_91_io_out ? io_r_37_b : _GEN_18536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18538 = 8'h26 == r_count_91_io_out ? io_r_38_b : _GEN_18537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18539 = 8'h27 == r_count_91_io_out ? io_r_39_b : _GEN_18538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18540 = 8'h28 == r_count_91_io_out ? io_r_40_b : _GEN_18539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18541 = 8'h29 == r_count_91_io_out ? io_r_41_b : _GEN_18540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18542 = 8'h2a == r_count_91_io_out ? io_r_42_b : _GEN_18541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18543 = 8'h2b == r_count_91_io_out ? io_r_43_b : _GEN_18542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18544 = 8'h2c == r_count_91_io_out ? io_r_44_b : _GEN_18543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18545 = 8'h2d == r_count_91_io_out ? io_r_45_b : _GEN_18544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18546 = 8'h2e == r_count_91_io_out ? io_r_46_b : _GEN_18545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18547 = 8'h2f == r_count_91_io_out ? io_r_47_b : _GEN_18546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18548 = 8'h30 == r_count_91_io_out ? io_r_48_b : _GEN_18547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18549 = 8'h31 == r_count_91_io_out ? io_r_49_b : _GEN_18548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18550 = 8'h32 == r_count_91_io_out ? io_r_50_b : _GEN_18549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18551 = 8'h33 == r_count_91_io_out ? io_r_51_b : _GEN_18550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18552 = 8'h34 == r_count_91_io_out ? io_r_52_b : _GEN_18551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18553 = 8'h35 == r_count_91_io_out ? io_r_53_b : _GEN_18552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18554 = 8'h36 == r_count_91_io_out ? io_r_54_b : _GEN_18553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18555 = 8'h37 == r_count_91_io_out ? io_r_55_b : _GEN_18554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18556 = 8'h38 == r_count_91_io_out ? io_r_56_b : _GEN_18555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18557 = 8'h39 == r_count_91_io_out ? io_r_57_b : _GEN_18556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18558 = 8'h3a == r_count_91_io_out ? io_r_58_b : _GEN_18557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18559 = 8'h3b == r_count_91_io_out ? io_r_59_b : _GEN_18558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18560 = 8'h3c == r_count_91_io_out ? io_r_60_b : _GEN_18559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18561 = 8'h3d == r_count_91_io_out ? io_r_61_b : _GEN_18560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18562 = 8'h3e == r_count_91_io_out ? io_r_62_b : _GEN_18561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18563 = 8'h3f == r_count_91_io_out ? io_r_63_b : _GEN_18562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18564 = 8'h40 == r_count_91_io_out ? io_r_64_b : _GEN_18563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18565 = 8'h41 == r_count_91_io_out ? io_r_65_b : _GEN_18564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18566 = 8'h42 == r_count_91_io_out ? io_r_66_b : _GEN_18565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18567 = 8'h43 == r_count_91_io_out ? io_r_67_b : _GEN_18566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18568 = 8'h44 == r_count_91_io_out ? io_r_68_b : _GEN_18567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18569 = 8'h45 == r_count_91_io_out ? io_r_69_b : _GEN_18568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18570 = 8'h46 == r_count_91_io_out ? io_r_70_b : _GEN_18569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18571 = 8'h47 == r_count_91_io_out ? io_r_71_b : _GEN_18570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18572 = 8'h48 == r_count_91_io_out ? io_r_72_b : _GEN_18571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18573 = 8'h49 == r_count_91_io_out ? io_r_73_b : _GEN_18572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18574 = 8'h4a == r_count_91_io_out ? io_r_74_b : _GEN_18573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18575 = 8'h4b == r_count_91_io_out ? io_r_75_b : _GEN_18574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18576 = 8'h4c == r_count_91_io_out ? io_r_76_b : _GEN_18575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18577 = 8'h4d == r_count_91_io_out ? io_r_77_b : _GEN_18576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18578 = 8'h4e == r_count_91_io_out ? io_r_78_b : _GEN_18577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18579 = 8'h4f == r_count_91_io_out ? io_r_79_b : _GEN_18578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18580 = 8'h50 == r_count_91_io_out ? io_r_80_b : _GEN_18579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18581 = 8'h51 == r_count_91_io_out ? io_r_81_b : _GEN_18580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18582 = 8'h52 == r_count_91_io_out ? io_r_82_b : _GEN_18581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18583 = 8'h53 == r_count_91_io_out ? io_r_83_b : _GEN_18582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18584 = 8'h54 == r_count_91_io_out ? io_r_84_b : _GEN_18583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18585 = 8'h55 == r_count_91_io_out ? io_r_85_b : _GEN_18584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18586 = 8'h56 == r_count_91_io_out ? io_r_86_b : _GEN_18585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18587 = 8'h57 == r_count_91_io_out ? io_r_87_b : _GEN_18586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18588 = 8'h58 == r_count_91_io_out ? io_r_88_b : _GEN_18587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18589 = 8'h59 == r_count_91_io_out ? io_r_89_b : _GEN_18588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18590 = 8'h5a == r_count_91_io_out ? io_r_90_b : _GEN_18589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18591 = 8'h5b == r_count_91_io_out ? io_r_91_b : _GEN_18590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18592 = 8'h5c == r_count_91_io_out ? io_r_92_b : _GEN_18591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18593 = 8'h5d == r_count_91_io_out ? io_r_93_b : _GEN_18592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18594 = 8'h5e == r_count_91_io_out ? io_r_94_b : _GEN_18593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18595 = 8'h5f == r_count_91_io_out ? io_r_95_b : _GEN_18594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18596 = 8'h60 == r_count_91_io_out ? io_r_96_b : _GEN_18595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18597 = 8'h61 == r_count_91_io_out ? io_r_97_b : _GEN_18596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18598 = 8'h62 == r_count_91_io_out ? io_r_98_b : _GEN_18597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18599 = 8'h63 == r_count_91_io_out ? io_r_99_b : _GEN_18598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18600 = 8'h64 == r_count_91_io_out ? io_r_100_b : _GEN_18599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18601 = 8'h65 == r_count_91_io_out ? io_r_101_b : _GEN_18600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18602 = 8'h66 == r_count_91_io_out ? io_r_102_b : _GEN_18601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18603 = 8'h67 == r_count_91_io_out ? io_r_103_b : _GEN_18602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18604 = 8'h68 == r_count_91_io_out ? io_r_104_b : _GEN_18603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18605 = 8'h69 == r_count_91_io_out ? io_r_105_b : _GEN_18604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18606 = 8'h6a == r_count_91_io_out ? io_r_106_b : _GEN_18605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18607 = 8'h6b == r_count_91_io_out ? io_r_107_b : _GEN_18606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18608 = 8'h6c == r_count_91_io_out ? io_r_108_b : _GEN_18607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18609 = 8'h6d == r_count_91_io_out ? io_r_109_b : _GEN_18608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18610 = 8'h6e == r_count_91_io_out ? io_r_110_b : _GEN_18609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18611 = 8'h6f == r_count_91_io_out ? io_r_111_b : _GEN_18610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18612 = 8'h70 == r_count_91_io_out ? io_r_112_b : _GEN_18611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18613 = 8'h71 == r_count_91_io_out ? io_r_113_b : _GEN_18612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18614 = 8'h72 == r_count_91_io_out ? io_r_114_b : _GEN_18613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18615 = 8'h73 == r_count_91_io_out ? io_r_115_b : _GEN_18614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18616 = 8'h74 == r_count_91_io_out ? io_r_116_b : _GEN_18615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18617 = 8'h75 == r_count_91_io_out ? io_r_117_b : _GEN_18616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18618 = 8'h76 == r_count_91_io_out ? io_r_118_b : _GEN_18617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18619 = 8'h77 == r_count_91_io_out ? io_r_119_b : _GEN_18618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18620 = 8'h78 == r_count_91_io_out ? io_r_120_b : _GEN_18619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18621 = 8'h79 == r_count_91_io_out ? io_r_121_b : _GEN_18620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18622 = 8'h7a == r_count_91_io_out ? io_r_122_b : _GEN_18621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18623 = 8'h7b == r_count_91_io_out ? io_r_123_b : _GEN_18622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18624 = 8'h7c == r_count_91_io_out ? io_r_124_b : _GEN_18623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18625 = 8'h7d == r_count_91_io_out ? io_r_125_b : _GEN_18624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18626 = 8'h7e == r_count_91_io_out ? io_r_126_b : _GEN_18625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18627 = 8'h7f == r_count_91_io_out ? io_r_127_b : _GEN_18626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18628 = 8'h80 == r_count_91_io_out ? io_r_128_b : _GEN_18627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18629 = 8'h81 == r_count_91_io_out ? io_r_129_b : _GEN_18628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18630 = 8'h82 == r_count_91_io_out ? io_r_130_b : _GEN_18629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18631 = 8'h83 == r_count_91_io_out ? io_r_131_b : _GEN_18630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18632 = 8'h84 == r_count_91_io_out ? io_r_132_b : _GEN_18631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18633 = 8'h85 == r_count_91_io_out ? io_r_133_b : _GEN_18632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18634 = 8'h86 == r_count_91_io_out ? io_r_134_b : _GEN_18633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18635 = 8'h87 == r_count_91_io_out ? io_r_135_b : _GEN_18634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18636 = 8'h88 == r_count_91_io_out ? io_r_136_b : _GEN_18635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18637 = 8'h89 == r_count_91_io_out ? io_r_137_b : _GEN_18636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18638 = 8'h8a == r_count_91_io_out ? io_r_138_b : _GEN_18637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18639 = 8'h8b == r_count_91_io_out ? io_r_139_b : _GEN_18638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18640 = 8'h8c == r_count_91_io_out ? io_r_140_b : _GEN_18639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18641 = 8'h8d == r_count_91_io_out ? io_r_141_b : _GEN_18640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18642 = 8'h8e == r_count_91_io_out ? io_r_142_b : _GEN_18641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18643 = 8'h8f == r_count_91_io_out ? io_r_143_b : _GEN_18642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18644 = 8'h90 == r_count_91_io_out ? io_r_144_b : _GEN_18643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18645 = 8'h91 == r_count_91_io_out ? io_r_145_b : _GEN_18644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18646 = 8'h92 == r_count_91_io_out ? io_r_146_b : _GEN_18645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18647 = 8'h93 == r_count_91_io_out ? io_r_147_b : _GEN_18646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18648 = 8'h94 == r_count_91_io_out ? io_r_148_b : _GEN_18647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18649 = 8'h95 == r_count_91_io_out ? io_r_149_b : _GEN_18648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18650 = 8'h96 == r_count_91_io_out ? io_r_150_b : _GEN_18649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18651 = 8'h97 == r_count_91_io_out ? io_r_151_b : _GEN_18650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18652 = 8'h98 == r_count_91_io_out ? io_r_152_b : _GEN_18651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18653 = 8'h99 == r_count_91_io_out ? io_r_153_b : _GEN_18652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18654 = 8'h9a == r_count_91_io_out ? io_r_154_b : _GEN_18653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18655 = 8'h9b == r_count_91_io_out ? io_r_155_b : _GEN_18654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18656 = 8'h9c == r_count_91_io_out ? io_r_156_b : _GEN_18655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18657 = 8'h9d == r_count_91_io_out ? io_r_157_b : _GEN_18656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18658 = 8'h9e == r_count_91_io_out ? io_r_158_b : _GEN_18657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18659 = 8'h9f == r_count_91_io_out ? io_r_159_b : _GEN_18658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18660 = 8'ha0 == r_count_91_io_out ? io_r_160_b : _GEN_18659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18661 = 8'ha1 == r_count_91_io_out ? io_r_161_b : _GEN_18660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18662 = 8'ha2 == r_count_91_io_out ? io_r_162_b : _GEN_18661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18663 = 8'ha3 == r_count_91_io_out ? io_r_163_b : _GEN_18662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18664 = 8'ha4 == r_count_91_io_out ? io_r_164_b : _GEN_18663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18665 = 8'ha5 == r_count_91_io_out ? io_r_165_b : _GEN_18664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18666 = 8'ha6 == r_count_91_io_out ? io_r_166_b : _GEN_18665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18667 = 8'ha7 == r_count_91_io_out ? io_r_167_b : _GEN_18666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18668 = 8'ha8 == r_count_91_io_out ? io_r_168_b : _GEN_18667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18669 = 8'ha9 == r_count_91_io_out ? io_r_169_b : _GEN_18668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18670 = 8'haa == r_count_91_io_out ? io_r_170_b : _GEN_18669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18671 = 8'hab == r_count_91_io_out ? io_r_171_b : _GEN_18670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18672 = 8'hac == r_count_91_io_out ? io_r_172_b : _GEN_18671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18673 = 8'had == r_count_91_io_out ? io_r_173_b : _GEN_18672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18674 = 8'hae == r_count_91_io_out ? io_r_174_b : _GEN_18673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18675 = 8'haf == r_count_91_io_out ? io_r_175_b : _GEN_18674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18676 = 8'hb0 == r_count_91_io_out ? io_r_176_b : _GEN_18675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18677 = 8'hb1 == r_count_91_io_out ? io_r_177_b : _GEN_18676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18678 = 8'hb2 == r_count_91_io_out ? io_r_178_b : _GEN_18677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18679 = 8'hb3 == r_count_91_io_out ? io_r_179_b : _GEN_18678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18680 = 8'hb4 == r_count_91_io_out ? io_r_180_b : _GEN_18679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18681 = 8'hb5 == r_count_91_io_out ? io_r_181_b : _GEN_18680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18682 = 8'hb6 == r_count_91_io_out ? io_r_182_b : _GEN_18681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18683 = 8'hb7 == r_count_91_io_out ? io_r_183_b : _GEN_18682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18684 = 8'hb8 == r_count_91_io_out ? io_r_184_b : _GEN_18683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18685 = 8'hb9 == r_count_91_io_out ? io_r_185_b : _GEN_18684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18686 = 8'hba == r_count_91_io_out ? io_r_186_b : _GEN_18685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18687 = 8'hbb == r_count_91_io_out ? io_r_187_b : _GEN_18686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18688 = 8'hbc == r_count_91_io_out ? io_r_188_b : _GEN_18687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18689 = 8'hbd == r_count_91_io_out ? io_r_189_b : _GEN_18688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18690 = 8'hbe == r_count_91_io_out ? io_r_190_b : _GEN_18689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18691 = 8'hbf == r_count_91_io_out ? io_r_191_b : _GEN_18690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18692 = 8'hc0 == r_count_91_io_out ? io_r_192_b : _GEN_18691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18693 = 8'hc1 == r_count_91_io_out ? io_r_193_b : _GEN_18692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18694 = 8'hc2 == r_count_91_io_out ? io_r_194_b : _GEN_18693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18695 = 8'hc3 == r_count_91_io_out ? io_r_195_b : _GEN_18694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18696 = 8'hc4 == r_count_91_io_out ? io_r_196_b : _GEN_18695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18697 = 8'hc5 == r_count_91_io_out ? io_r_197_b : _GEN_18696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18698 = 8'hc6 == r_count_91_io_out ? io_r_198_b : _GEN_18697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18701 = 8'h1 == r_count_92_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18702 = 8'h2 == r_count_92_io_out ? io_r_2_b : _GEN_18701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18703 = 8'h3 == r_count_92_io_out ? io_r_3_b : _GEN_18702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18704 = 8'h4 == r_count_92_io_out ? io_r_4_b : _GEN_18703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18705 = 8'h5 == r_count_92_io_out ? io_r_5_b : _GEN_18704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18706 = 8'h6 == r_count_92_io_out ? io_r_6_b : _GEN_18705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18707 = 8'h7 == r_count_92_io_out ? io_r_7_b : _GEN_18706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18708 = 8'h8 == r_count_92_io_out ? io_r_8_b : _GEN_18707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18709 = 8'h9 == r_count_92_io_out ? io_r_9_b : _GEN_18708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18710 = 8'ha == r_count_92_io_out ? io_r_10_b : _GEN_18709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18711 = 8'hb == r_count_92_io_out ? io_r_11_b : _GEN_18710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18712 = 8'hc == r_count_92_io_out ? io_r_12_b : _GEN_18711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18713 = 8'hd == r_count_92_io_out ? io_r_13_b : _GEN_18712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18714 = 8'he == r_count_92_io_out ? io_r_14_b : _GEN_18713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18715 = 8'hf == r_count_92_io_out ? io_r_15_b : _GEN_18714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18716 = 8'h10 == r_count_92_io_out ? io_r_16_b : _GEN_18715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18717 = 8'h11 == r_count_92_io_out ? io_r_17_b : _GEN_18716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18718 = 8'h12 == r_count_92_io_out ? io_r_18_b : _GEN_18717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18719 = 8'h13 == r_count_92_io_out ? io_r_19_b : _GEN_18718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18720 = 8'h14 == r_count_92_io_out ? io_r_20_b : _GEN_18719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18721 = 8'h15 == r_count_92_io_out ? io_r_21_b : _GEN_18720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18722 = 8'h16 == r_count_92_io_out ? io_r_22_b : _GEN_18721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18723 = 8'h17 == r_count_92_io_out ? io_r_23_b : _GEN_18722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18724 = 8'h18 == r_count_92_io_out ? io_r_24_b : _GEN_18723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18725 = 8'h19 == r_count_92_io_out ? io_r_25_b : _GEN_18724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18726 = 8'h1a == r_count_92_io_out ? io_r_26_b : _GEN_18725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18727 = 8'h1b == r_count_92_io_out ? io_r_27_b : _GEN_18726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18728 = 8'h1c == r_count_92_io_out ? io_r_28_b : _GEN_18727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18729 = 8'h1d == r_count_92_io_out ? io_r_29_b : _GEN_18728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18730 = 8'h1e == r_count_92_io_out ? io_r_30_b : _GEN_18729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18731 = 8'h1f == r_count_92_io_out ? io_r_31_b : _GEN_18730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18732 = 8'h20 == r_count_92_io_out ? io_r_32_b : _GEN_18731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18733 = 8'h21 == r_count_92_io_out ? io_r_33_b : _GEN_18732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18734 = 8'h22 == r_count_92_io_out ? io_r_34_b : _GEN_18733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18735 = 8'h23 == r_count_92_io_out ? io_r_35_b : _GEN_18734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18736 = 8'h24 == r_count_92_io_out ? io_r_36_b : _GEN_18735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18737 = 8'h25 == r_count_92_io_out ? io_r_37_b : _GEN_18736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18738 = 8'h26 == r_count_92_io_out ? io_r_38_b : _GEN_18737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18739 = 8'h27 == r_count_92_io_out ? io_r_39_b : _GEN_18738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18740 = 8'h28 == r_count_92_io_out ? io_r_40_b : _GEN_18739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18741 = 8'h29 == r_count_92_io_out ? io_r_41_b : _GEN_18740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18742 = 8'h2a == r_count_92_io_out ? io_r_42_b : _GEN_18741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18743 = 8'h2b == r_count_92_io_out ? io_r_43_b : _GEN_18742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18744 = 8'h2c == r_count_92_io_out ? io_r_44_b : _GEN_18743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18745 = 8'h2d == r_count_92_io_out ? io_r_45_b : _GEN_18744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18746 = 8'h2e == r_count_92_io_out ? io_r_46_b : _GEN_18745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18747 = 8'h2f == r_count_92_io_out ? io_r_47_b : _GEN_18746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18748 = 8'h30 == r_count_92_io_out ? io_r_48_b : _GEN_18747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18749 = 8'h31 == r_count_92_io_out ? io_r_49_b : _GEN_18748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18750 = 8'h32 == r_count_92_io_out ? io_r_50_b : _GEN_18749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18751 = 8'h33 == r_count_92_io_out ? io_r_51_b : _GEN_18750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18752 = 8'h34 == r_count_92_io_out ? io_r_52_b : _GEN_18751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18753 = 8'h35 == r_count_92_io_out ? io_r_53_b : _GEN_18752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18754 = 8'h36 == r_count_92_io_out ? io_r_54_b : _GEN_18753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18755 = 8'h37 == r_count_92_io_out ? io_r_55_b : _GEN_18754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18756 = 8'h38 == r_count_92_io_out ? io_r_56_b : _GEN_18755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18757 = 8'h39 == r_count_92_io_out ? io_r_57_b : _GEN_18756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18758 = 8'h3a == r_count_92_io_out ? io_r_58_b : _GEN_18757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18759 = 8'h3b == r_count_92_io_out ? io_r_59_b : _GEN_18758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18760 = 8'h3c == r_count_92_io_out ? io_r_60_b : _GEN_18759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18761 = 8'h3d == r_count_92_io_out ? io_r_61_b : _GEN_18760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18762 = 8'h3e == r_count_92_io_out ? io_r_62_b : _GEN_18761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18763 = 8'h3f == r_count_92_io_out ? io_r_63_b : _GEN_18762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18764 = 8'h40 == r_count_92_io_out ? io_r_64_b : _GEN_18763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18765 = 8'h41 == r_count_92_io_out ? io_r_65_b : _GEN_18764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18766 = 8'h42 == r_count_92_io_out ? io_r_66_b : _GEN_18765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18767 = 8'h43 == r_count_92_io_out ? io_r_67_b : _GEN_18766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18768 = 8'h44 == r_count_92_io_out ? io_r_68_b : _GEN_18767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18769 = 8'h45 == r_count_92_io_out ? io_r_69_b : _GEN_18768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18770 = 8'h46 == r_count_92_io_out ? io_r_70_b : _GEN_18769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18771 = 8'h47 == r_count_92_io_out ? io_r_71_b : _GEN_18770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18772 = 8'h48 == r_count_92_io_out ? io_r_72_b : _GEN_18771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18773 = 8'h49 == r_count_92_io_out ? io_r_73_b : _GEN_18772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18774 = 8'h4a == r_count_92_io_out ? io_r_74_b : _GEN_18773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18775 = 8'h4b == r_count_92_io_out ? io_r_75_b : _GEN_18774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18776 = 8'h4c == r_count_92_io_out ? io_r_76_b : _GEN_18775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18777 = 8'h4d == r_count_92_io_out ? io_r_77_b : _GEN_18776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18778 = 8'h4e == r_count_92_io_out ? io_r_78_b : _GEN_18777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18779 = 8'h4f == r_count_92_io_out ? io_r_79_b : _GEN_18778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18780 = 8'h50 == r_count_92_io_out ? io_r_80_b : _GEN_18779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18781 = 8'h51 == r_count_92_io_out ? io_r_81_b : _GEN_18780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18782 = 8'h52 == r_count_92_io_out ? io_r_82_b : _GEN_18781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18783 = 8'h53 == r_count_92_io_out ? io_r_83_b : _GEN_18782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18784 = 8'h54 == r_count_92_io_out ? io_r_84_b : _GEN_18783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18785 = 8'h55 == r_count_92_io_out ? io_r_85_b : _GEN_18784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18786 = 8'h56 == r_count_92_io_out ? io_r_86_b : _GEN_18785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18787 = 8'h57 == r_count_92_io_out ? io_r_87_b : _GEN_18786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18788 = 8'h58 == r_count_92_io_out ? io_r_88_b : _GEN_18787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18789 = 8'h59 == r_count_92_io_out ? io_r_89_b : _GEN_18788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18790 = 8'h5a == r_count_92_io_out ? io_r_90_b : _GEN_18789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18791 = 8'h5b == r_count_92_io_out ? io_r_91_b : _GEN_18790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18792 = 8'h5c == r_count_92_io_out ? io_r_92_b : _GEN_18791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18793 = 8'h5d == r_count_92_io_out ? io_r_93_b : _GEN_18792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18794 = 8'h5e == r_count_92_io_out ? io_r_94_b : _GEN_18793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18795 = 8'h5f == r_count_92_io_out ? io_r_95_b : _GEN_18794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18796 = 8'h60 == r_count_92_io_out ? io_r_96_b : _GEN_18795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18797 = 8'h61 == r_count_92_io_out ? io_r_97_b : _GEN_18796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18798 = 8'h62 == r_count_92_io_out ? io_r_98_b : _GEN_18797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18799 = 8'h63 == r_count_92_io_out ? io_r_99_b : _GEN_18798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18800 = 8'h64 == r_count_92_io_out ? io_r_100_b : _GEN_18799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18801 = 8'h65 == r_count_92_io_out ? io_r_101_b : _GEN_18800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18802 = 8'h66 == r_count_92_io_out ? io_r_102_b : _GEN_18801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18803 = 8'h67 == r_count_92_io_out ? io_r_103_b : _GEN_18802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18804 = 8'h68 == r_count_92_io_out ? io_r_104_b : _GEN_18803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18805 = 8'h69 == r_count_92_io_out ? io_r_105_b : _GEN_18804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18806 = 8'h6a == r_count_92_io_out ? io_r_106_b : _GEN_18805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18807 = 8'h6b == r_count_92_io_out ? io_r_107_b : _GEN_18806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18808 = 8'h6c == r_count_92_io_out ? io_r_108_b : _GEN_18807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18809 = 8'h6d == r_count_92_io_out ? io_r_109_b : _GEN_18808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18810 = 8'h6e == r_count_92_io_out ? io_r_110_b : _GEN_18809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18811 = 8'h6f == r_count_92_io_out ? io_r_111_b : _GEN_18810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18812 = 8'h70 == r_count_92_io_out ? io_r_112_b : _GEN_18811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18813 = 8'h71 == r_count_92_io_out ? io_r_113_b : _GEN_18812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18814 = 8'h72 == r_count_92_io_out ? io_r_114_b : _GEN_18813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18815 = 8'h73 == r_count_92_io_out ? io_r_115_b : _GEN_18814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18816 = 8'h74 == r_count_92_io_out ? io_r_116_b : _GEN_18815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18817 = 8'h75 == r_count_92_io_out ? io_r_117_b : _GEN_18816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18818 = 8'h76 == r_count_92_io_out ? io_r_118_b : _GEN_18817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18819 = 8'h77 == r_count_92_io_out ? io_r_119_b : _GEN_18818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18820 = 8'h78 == r_count_92_io_out ? io_r_120_b : _GEN_18819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18821 = 8'h79 == r_count_92_io_out ? io_r_121_b : _GEN_18820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18822 = 8'h7a == r_count_92_io_out ? io_r_122_b : _GEN_18821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18823 = 8'h7b == r_count_92_io_out ? io_r_123_b : _GEN_18822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18824 = 8'h7c == r_count_92_io_out ? io_r_124_b : _GEN_18823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18825 = 8'h7d == r_count_92_io_out ? io_r_125_b : _GEN_18824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18826 = 8'h7e == r_count_92_io_out ? io_r_126_b : _GEN_18825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18827 = 8'h7f == r_count_92_io_out ? io_r_127_b : _GEN_18826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18828 = 8'h80 == r_count_92_io_out ? io_r_128_b : _GEN_18827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18829 = 8'h81 == r_count_92_io_out ? io_r_129_b : _GEN_18828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18830 = 8'h82 == r_count_92_io_out ? io_r_130_b : _GEN_18829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18831 = 8'h83 == r_count_92_io_out ? io_r_131_b : _GEN_18830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18832 = 8'h84 == r_count_92_io_out ? io_r_132_b : _GEN_18831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18833 = 8'h85 == r_count_92_io_out ? io_r_133_b : _GEN_18832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18834 = 8'h86 == r_count_92_io_out ? io_r_134_b : _GEN_18833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18835 = 8'h87 == r_count_92_io_out ? io_r_135_b : _GEN_18834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18836 = 8'h88 == r_count_92_io_out ? io_r_136_b : _GEN_18835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18837 = 8'h89 == r_count_92_io_out ? io_r_137_b : _GEN_18836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18838 = 8'h8a == r_count_92_io_out ? io_r_138_b : _GEN_18837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18839 = 8'h8b == r_count_92_io_out ? io_r_139_b : _GEN_18838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18840 = 8'h8c == r_count_92_io_out ? io_r_140_b : _GEN_18839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18841 = 8'h8d == r_count_92_io_out ? io_r_141_b : _GEN_18840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18842 = 8'h8e == r_count_92_io_out ? io_r_142_b : _GEN_18841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18843 = 8'h8f == r_count_92_io_out ? io_r_143_b : _GEN_18842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18844 = 8'h90 == r_count_92_io_out ? io_r_144_b : _GEN_18843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18845 = 8'h91 == r_count_92_io_out ? io_r_145_b : _GEN_18844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18846 = 8'h92 == r_count_92_io_out ? io_r_146_b : _GEN_18845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18847 = 8'h93 == r_count_92_io_out ? io_r_147_b : _GEN_18846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18848 = 8'h94 == r_count_92_io_out ? io_r_148_b : _GEN_18847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18849 = 8'h95 == r_count_92_io_out ? io_r_149_b : _GEN_18848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18850 = 8'h96 == r_count_92_io_out ? io_r_150_b : _GEN_18849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18851 = 8'h97 == r_count_92_io_out ? io_r_151_b : _GEN_18850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18852 = 8'h98 == r_count_92_io_out ? io_r_152_b : _GEN_18851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18853 = 8'h99 == r_count_92_io_out ? io_r_153_b : _GEN_18852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18854 = 8'h9a == r_count_92_io_out ? io_r_154_b : _GEN_18853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18855 = 8'h9b == r_count_92_io_out ? io_r_155_b : _GEN_18854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18856 = 8'h9c == r_count_92_io_out ? io_r_156_b : _GEN_18855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18857 = 8'h9d == r_count_92_io_out ? io_r_157_b : _GEN_18856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18858 = 8'h9e == r_count_92_io_out ? io_r_158_b : _GEN_18857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18859 = 8'h9f == r_count_92_io_out ? io_r_159_b : _GEN_18858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18860 = 8'ha0 == r_count_92_io_out ? io_r_160_b : _GEN_18859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18861 = 8'ha1 == r_count_92_io_out ? io_r_161_b : _GEN_18860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18862 = 8'ha2 == r_count_92_io_out ? io_r_162_b : _GEN_18861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18863 = 8'ha3 == r_count_92_io_out ? io_r_163_b : _GEN_18862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18864 = 8'ha4 == r_count_92_io_out ? io_r_164_b : _GEN_18863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18865 = 8'ha5 == r_count_92_io_out ? io_r_165_b : _GEN_18864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18866 = 8'ha6 == r_count_92_io_out ? io_r_166_b : _GEN_18865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18867 = 8'ha7 == r_count_92_io_out ? io_r_167_b : _GEN_18866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18868 = 8'ha8 == r_count_92_io_out ? io_r_168_b : _GEN_18867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18869 = 8'ha9 == r_count_92_io_out ? io_r_169_b : _GEN_18868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18870 = 8'haa == r_count_92_io_out ? io_r_170_b : _GEN_18869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18871 = 8'hab == r_count_92_io_out ? io_r_171_b : _GEN_18870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18872 = 8'hac == r_count_92_io_out ? io_r_172_b : _GEN_18871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18873 = 8'had == r_count_92_io_out ? io_r_173_b : _GEN_18872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18874 = 8'hae == r_count_92_io_out ? io_r_174_b : _GEN_18873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18875 = 8'haf == r_count_92_io_out ? io_r_175_b : _GEN_18874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18876 = 8'hb0 == r_count_92_io_out ? io_r_176_b : _GEN_18875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18877 = 8'hb1 == r_count_92_io_out ? io_r_177_b : _GEN_18876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18878 = 8'hb2 == r_count_92_io_out ? io_r_178_b : _GEN_18877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18879 = 8'hb3 == r_count_92_io_out ? io_r_179_b : _GEN_18878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18880 = 8'hb4 == r_count_92_io_out ? io_r_180_b : _GEN_18879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18881 = 8'hb5 == r_count_92_io_out ? io_r_181_b : _GEN_18880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18882 = 8'hb6 == r_count_92_io_out ? io_r_182_b : _GEN_18881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18883 = 8'hb7 == r_count_92_io_out ? io_r_183_b : _GEN_18882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18884 = 8'hb8 == r_count_92_io_out ? io_r_184_b : _GEN_18883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18885 = 8'hb9 == r_count_92_io_out ? io_r_185_b : _GEN_18884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18886 = 8'hba == r_count_92_io_out ? io_r_186_b : _GEN_18885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18887 = 8'hbb == r_count_92_io_out ? io_r_187_b : _GEN_18886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18888 = 8'hbc == r_count_92_io_out ? io_r_188_b : _GEN_18887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18889 = 8'hbd == r_count_92_io_out ? io_r_189_b : _GEN_18888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18890 = 8'hbe == r_count_92_io_out ? io_r_190_b : _GEN_18889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18891 = 8'hbf == r_count_92_io_out ? io_r_191_b : _GEN_18890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18892 = 8'hc0 == r_count_92_io_out ? io_r_192_b : _GEN_18891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18893 = 8'hc1 == r_count_92_io_out ? io_r_193_b : _GEN_18892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18894 = 8'hc2 == r_count_92_io_out ? io_r_194_b : _GEN_18893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18895 = 8'hc3 == r_count_92_io_out ? io_r_195_b : _GEN_18894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18896 = 8'hc4 == r_count_92_io_out ? io_r_196_b : _GEN_18895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18897 = 8'hc5 == r_count_92_io_out ? io_r_197_b : _GEN_18896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18898 = 8'hc6 == r_count_92_io_out ? io_r_198_b : _GEN_18897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18901 = 8'h1 == r_count_93_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18902 = 8'h2 == r_count_93_io_out ? io_r_2_b : _GEN_18901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18903 = 8'h3 == r_count_93_io_out ? io_r_3_b : _GEN_18902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18904 = 8'h4 == r_count_93_io_out ? io_r_4_b : _GEN_18903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18905 = 8'h5 == r_count_93_io_out ? io_r_5_b : _GEN_18904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18906 = 8'h6 == r_count_93_io_out ? io_r_6_b : _GEN_18905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18907 = 8'h7 == r_count_93_io_out ? io_r_7_b : _GEN_18906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18908 = 8'h8 == r_count_93_io_out ? io_r_8_b : _GEN_18907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18909 = 8'h9 == r_count_93_io_out ? io_r_9_b : _GEN_18908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18910 = 8'ha == r_count_93_io_out ? io_r_10_b : _GEN_18909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18911 = 8'hb == r_count_93_io_out ? io_r_11_b : _GEN_18910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18912 = 8'hc == r_count_93_io_out ? io_r_12_b : _GEN_18911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18913 = 8'hd == r_count_93_io_out ? io_r_13_b : _GEN_18912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18914 = 8'he == r_count_93_io_out ? io_r_14_b : _GEN_18913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18915 = 8'hf == r_count_93_io_out ? io_r_15_b : _GEN_18914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18916 = 8'h10 == r_count_93_io_out ? io_r_16_b : _GEN_18915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18917 = 8'h11 == r_count_93_io_out ? io_r_17_b : _GEN_18916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18918 = 8'h12 == r_count_93_io_out ? io_r_18_b : _GEN_18917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18919 = 8'h13 == r_count_93_io_out ? io_r_19_b : _GEN_18918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18920 = 8'h14 == r_count_93_io_out ? io_r_20_b : _GEN_18919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18921 = 8'h15 == r_count_93_io_out ? io_r_21_b : _GEN_18920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18922 = 8'h16 == r_count_93_io_out ? io_r_22_b : _GEN_18921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18923 = 8'h17 == r_count_93_io_out ? io_r_23_b : _GEN_18922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18924 = 8'h18 == r_count_93_io_out ? io_r_24_b : _GEN_18923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18925 = 8'h19 == r_count_93_io_out ? io_r_25_b : _GEN_18924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18926 = 8'h1a == r_count_93_io_out ? io_r_26_b : _GEN_18925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18927 = 8'h1b == r_count_93_io_out ? io_r_27_b : _GEN_18926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18928 = 8'h1c == r_count_93_io_out ? io_r_28_b : _GEN_18927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18929 = 8'h1d == r_count_93_io_out ? io_r_29_b : _GEN_18928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18930 = 8'h1e == r_count_93_io_out ? io_r_30_b : _GEN_18929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18931 = 8'h1f == r_count_93_io_out ? io_r_31_b : _GEN_18930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18932 = 8'h20 == r_count_93_io_out ? io_r_32_b : _GEN_18931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18933 = 8'h21 == r_count_93_io_out ? io_r_33_b : _GEN_18932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18934 = 8'h22 == r_count_93_io_out ? io_r_34_b : _GEN_18933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18935 = 8'h23 == r_count_93_io_out ? io_r_35_b : _GEN_18934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18936 = 8'h24 == r_count_93_io_out ? io_r_36_b : _GEN_18935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18937 = 8'h25 == r_count_93_io_out ? io_r_37_b : _GEN_18936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18938 = 8'h26 == r_count_93_io_out ? io_r_38_b : _GEN_18937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18939 = 8'h27 == r_count_93_io_out ? io_r_39_b : _GEN_18938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18940 = 8'h28 == r_count_93_io_out ? io_r_40_b : _GEN_18939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18941 = 8'h29 == r_count_93_io_out ? io_r_41_b : _GEN_18940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18942 = 8'h2a == r_count_93_io_out ? io_r_42_b : _GEN_18941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18943 = 8'h2b == r_count_93_io_out ? io_r_43_b : _GEN_18942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18944 = 8'h2c == r_count_93_io_out ? io_r_44_b : _GEN_18943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18945 = 8'h2d == r_count_93_io_out ? io_r_45_b : _GEN_18944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18946 = 8'h2e == r_count_93_io_out ? io_r_46_b : _GEN_18945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18947 = 8'h2f == r_count_93_io_out ? io_r_47_b : _GEN_18946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18948 = 8'h30 == r_count_93_io_out ? io_r_48_b : _GEN_18947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18949 = 8'h31 == r_count_93_io_out ? io_r_49_b : _GEN_18948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18950 = 8'h32 == r_count_93_io_out ? io_r_50_b : _GEN_18949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18951 = 8'h33 == r_count_93_io_out ? io_r_51_b : _GEN_18950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18952 = 8'h34 == r_count_93_io_out ? io_r_52_b : _GEN_18951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18953 = 8'h35 == r_count_93_io_out ? io_r_53_b : _GEN_18952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18954 = 8'h36 == r_count_93_io_out ? io_r_54_b : _GEN_18953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18955 = 8'h37 == r_count_93_io_out ? io_r_55_b : _GEN_18954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18956 = 8'h38 == r_count_93_io_out ? io_r_56_b : _GEN_18955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18957 = 8'h39 == r_count_93_io_out ? io_r_57_b : _GEN_18956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18958 = 8'h3a == r_count_93_io_out ? io_r_58_b : _GEN_18957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18959 = 8'h3b == r_count_93_io_out ? io_r_59_b : _GEN_18958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18960 = 8'h3c == r_count_93_io_out ? io_r_60_b : _GEN_18959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18961 = 8'h3d == r_count_93_io_out ? io_r_61_b : _GEN_18960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18962 = 8'h3e == r_count_93_io_out ? io_r_62_b : _GEN_18961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18963 = 8'h3f == r_count_93_io_out ? io_r_63_b : _GEN_18962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18964 = 8'h40 == r_count_93_io_out ? io_r_64_b : _GEN_18963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18965 = 8'h41 == r_count_93_io_out ? io_r_65_b : _GEN_18964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18966 = 8'h42 == r_count_93_io_out ? io_r_66_b : _GEN_18965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18967 = 8'h43 == r_count_93_io_out ? io_r_67_b : _GEN_18966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18968 = 8'h44 == r_count_93_io_out ? io_r_68_b : _GEN_18967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18969 = 8'h45 == r_count_93_io_out ? io_r_69_b : _GEN_18968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18970 = 8'h46 == r_count_93_io_out ? io_r_70_b : _GEN_18969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18971 = 8'h47 == r_count_93_io_out ? io_r_71_b : _GEN_18970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18972 = 8'h48 == r_count_93_io_out ? io_r_72_b : _GEN_18971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18973 = 8'h49 == r_count_93_io_out ? io_r_73_b : _GEN_18972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18974 = 8'h4a == r_count_93_io_out ? io_r_74_b : _GEN_18973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18975 = 8'h4b == r_count_93_io_out ? io_r_75_b : _GEN_18974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18976 = 8'h4c == r_count_93_io_out ? io_r_76_b : _GEN_18975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18977 = 8'h4d == r_count_93_io_out ? io_r_77_b : _GEN_18976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18978 = 8'h4e == r_count_93_io_out ? io_r_78_b : _GEN_18977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18979 = 8'h4f == r_count_93_io_out ? io_r_79_b : _GEN_18978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18980 = 8'h50 == r_count_93_io_out ? io_r_80_b : _GEN_18979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18981 = 8'h51 == r_count_93_io_out ? io_r_81_b : _GEN_18980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18982 = 8'h52 == r_count_93_io_out ? io_r_82_b : _GEN_18981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18983 = 8'h53 == r_count_93_io_out ? io_r_83_b : _GEN_18982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18984 = 8'h54 == r_count_93_io_out ? io_r_84_b : _GEN_18983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18985 = 8'h55 == r_count_93_io_out ? io_r_85_b : _GEN_18984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18986 = 8'h56 == r_count_93_io_out ? io_r_86_b : _GEN_18985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18987 = 8'h57 == r_count_93_io_out ? io_r_87_b : _GEN_18986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18988 = 8'h58 == r_count_93_io_out ? io_r_88_b : _GEN_18987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18989 = 8'h59 == r_count_93_io_out ? io_r_89_b : _GEN_18988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18990 = 8'h5a == r_count_93_io_out ? io_r_90_b : _GEN_18989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18991 = 8'h5b == r_count_93_io_out ? io_r_91_b : _GEN_18990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18992 = 8'h5c == r_count_93_io_out ? io_r_92_b : _GEN_18991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18993 = 8'h5d == r_count_93_io_out ? io_r_93_b : _GEN_18992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18994 = 8'h5e == r_count_93_io_out ? io_r_94_b : _GEN_18993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18995 = 8'h5f == r_count_93_io_out ? io_r_95_b : _GEN_18994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18996 = 8'h60 == r_count_93_io_out ? io_r_96_b : _GEN_18995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18997 = 8'h61 == r_count_93_io_out ? io_r_97_b : _GEN_18996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18998 = 8'h62 == r_count_93_io_out ? io_r_98_b : _GEN_18997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_18999 = 8'h63 == r_count_93_io_out ? io_r_99_b : _GEN_18998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19000 = 8'h64 == r_count_93_io_out ? io_r_100_b : _GEN_18999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19001 = 8'h65 == r_count_93_io_out ? io_r_101_b : _GEN_19000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19002 = 8'h66 == r_count_93_io_out ? io_r_102_b : _GEN_19001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19003 = 8'h67 == r_count_93_io_out ? io_r_103_b : _GEN_19002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19004 = 8'h68 == r_count_93_io_out ? io_r_104_b : _GEN_19003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19005 = 8'h69 == r_count_93_io_out ? io_r_105_b : _GEN_19004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19006 = 8'h6a == r_count_93_io_out ? io_r_106_b : _GEN_19005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19007 = 8'h6b == r_count_93_io_out ? io_r_107_b : _GEN_19006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19008 = 8'h6c == r_count_93_io_out ? io_r_108_b : _GEN_19007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19009 = 8'h6d == r_count_93_io_out ? io_r_109_b : _GEN_19008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19010 = 8'h6e == r_count_93_io_out ? io_r_110_b : _GEN_19009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19011 = 8'h6f == r_count_93_io_out ? io_r_111_b : _GEN_19010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19012 = 8'h70 == r_count_93_io_out ? io_r_112_b : _GEN_19011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19013 = 8'h71 == r_count_93_io_out ? io_r_113_b : _GEN_19012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19014 = 8'h72 == r_count_93_io_out ? io_r_114_b : _GEN_19013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19015 = 8'h73 == r_count_93_io_out ? io_r_115_b : _GEN_19014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19016 = 8'h74 == r_count_93_io_out ? io_r_116_b : _GEN_19015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19017 = 8'h75 == r_count_93_io_out ? io_r_117_b : _GEN_19016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19018 = 8'h76 == r_count_93_io_out ? io_r_118_b : _GEN_19017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19019 = 8'h77 == r_count_93_io_out ? io_r_119_b : _GEN_19018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19020 = 8'h78 == r_count_93_io_out ? io_r_120_b : _GEN_19019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19021 = 8'h79 == r_count_93_io_out ? io_r_121_b : _GEN_19020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19022 = 8'h7a == r_count_93_io_out ? io_r_122_b : _GEN_19021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19023 = 8'h7b == r_count_93_io_out ? io_r_123_b : _GEN_19022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19024 = 8'h7c == r_count_93_io_out ? io_r_124_b : _GEN_19023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19025 = 8'h7d == r_count_93_io_out ? io_r_125_b : _GEN_19024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19026 = 8'h7e == r_count_93_io_out ? io_r_126_b : _GEN_19025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19027 = 8'h7f == r_count_93_io_out ? io_r_127_b : _GEN_19026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19028 = 8'h80 == r_count_93_io_out ? io_r_128_b : _GEN_19027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19029 = 8'h81 == r_count_93_io_out ? io_r_129_b : _GEN_19028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19030 = 8'h82 == r_count_93_io_out ? io_r_130_b : _GEN_19029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19031 = 8'h83 == r_count_93_io_out ? io_r_131_b : _GEN_19030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19032 = 8'h84 == r_count_93_io_out ? io_r_132_b : _GEN_19031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19033 = 8'h85 == r_count_93_io_out ? io_r_133_b : _GEN_19032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19034 = 8'h86 == r_count_93_io_out ? io_r_134_b : _GEN_19033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19035 = 8'h87 == r_count_93_io_out ? io_r_135_b : _GEN_19034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19036 = 8'h88 == r_count_93_io_out ? io_r_136_b : _GEN_19035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19037 = 8'h89 == r_count_93_io_out ? io_r_137_b : _GEN_19036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19038 = 8'h8a == r_count_93_io_out ? io_r_138_b : _GEN_19037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19039 = 8'h8b == r_count_93_io_out ? io_r_139_b : _GEN_19038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19040 = 8'h8c == r_count_93_io_out ? io_r_140_b : _GEN_19039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19041 = 8'h8d == r_count_93_io_out ? io_r_141_b : _GEN_19040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19042 = 8'h8e == r_count_93_io_out ? io_r_142_b : _GEN_19041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19043 = 8'h8f == r_count_93_io_out ? io_r_143_b : _GEN_19042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19044 = 8'h90 == r_count_93_io_out ? io_r_144_b : _GEN_19043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19045 = 8'h91 == r_count_93_io_out ? io_r_145_b : _GEN_19044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19046 = 8'h92 == r_count_93_io_out ? io_r_146_b : _GEN_19045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19047 = 8'h93 == r_count_93_io_out ? io_r_147_b : _GEN_19046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19048 = 8'h94 == r_count_93_io_out ? io_r_148_b : _GEN_19047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19049 = 8'h95 == r_count_93_io_out ? io_r_149_b : _GEN_19048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19050 = 8'h96 == r_count_93_io_out ? io_r_150_b : _GEN_19049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19051 = 8'h97 == r_count_93_io_out ? io_r_151_b : _GEN_19050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19052 = 8'h98 == r_count_93_io_out ? io_r_152_b : _GEN_19051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19053 = 8'h99 == r_count_93_io_out ? io_r_153_b : _GEN_19052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19054 = 8'h9a == r_count_93_io_out ? io_r_154_b : _GEN_19053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19055 = 8'h9b == r_count_93_io_out ? io_r_155_b : _GEN_19054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19056 = 8'h9c == r_count_93_io_out ? io_r_156_b : _GEN_19055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19057 = 8'h9d == r_count_93_io_out ? io_r_157_b : _GEN_19056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19058 = 8'h9e == r_count_93_io_out ? io_r_158_b : _GEN_19057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19059 = 8'h9f == r_count_93_io_out ? io_r_159_b : _GEN_19058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19060 = 8'ha0 == r_count_93_io_out ? io_r_160_b : _GEN_19059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19061 = 8'ha1 == r_count_93_io_out ? io_r_161_b : _GEN_19060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19062 = 8'ha2 == r_count_93_io_out ? io_r_162_b : _GEN_19061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19063 = 8'ha3 == r_count_93_io_out ? io_r_163_b : _GEN_19062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19064 = 8'ha4 == r_count_93_io_out ? io_r_164_b : _GEN_19063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19065 = 8'ha5 == r_count_93_io_out ? io_r_165_b : _GEN_19064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19066 = 8'ha6 == r_count_93_io_out ? io_r_166_b : _GEN_19065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19067 = 8'ha7 == r_count_93_io_out ? io_r_167_b : _GEN_19066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19068 = 8'ha8 == r_count_93_io_out ? io_r_168_b : _GEN_19067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19069 = 8'ha9 == r_count_93_io_out ? io_r_169_b : _GEN_19068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19070 = 8'haa == r_count_93_io_out ? io_r_170_b : _GEN_19069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19071 = 8'hab == r_count_93_io_out ? io_r_171_b : _GEN_19070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19072 = 8'hac == r_count_93_io_out ? io_r_172_b : _GEN_19071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19073 = 8'had == r_count_93_io_out ? io_r_173_b : _GEN_19072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19074 = 8'hae == r_count_93_io_out ? io_r_174_b : _GEN_19073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19075 = 8'haf == r_count_93_io_out ? io_r_175_b : _GEN_19074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19076 = 8'hb0 == r_count_93_io_out ? io_r_176_b : _GEN_19075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19077 = 8'hb1 == r_count_93_io_out ? io_r_177_b : _GEN_19076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19078 = 8'hb2 == r_count_93_io_out ? io_r_178_b : _GEN_19077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19079 = 8'hb3 == r_count_93_io_out ? io_r_179_b : _GEN_19078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19080 = 8'hb4 == r_count_93_io_out ? io_r_180_b : _GEN_19079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19081 = 8'hb5 == r_count_93_io_out ? io_r_181_b : _GEN_19080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19082 = 8'hb6 == r_count_93_io_out ? io_r_182_b : _GEN_19081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19083 = 8'hb7 == r_count_93_io_out ? io_r_183_b : _GEN_19082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19084 = 8'hb8 == r_count_93_io_out ? io_r_184_b : _GEN_19083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19085 = 8'hb9 == r_count_93_io_out ? io_r_185_b : _GEN_19084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19086 = 8'hba == r_count_93_io_out ? io_r_186_b : _GEN_19085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19087 = 8'hbb == r_count_93_io_out ? io_r_187_b : _GEN_19086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19088 = 8'hbc == r_count_93_io_out ? io_r_188_b : _GEN_19087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19089 = 8'hbd == r_count_93_io_out ? io_r_189_b : _GEN_19088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19090 = 8'hbe == r_count_93_io_out ? io_r_190_b : _GEN_19089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19091 = 8'hbf == r_count_93_io_out ? io_r_191_b : _GEN_19090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19092 = 8'hc0 == r_count_93_io_out ? io_r_192_b : _GEN_19091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19093 = 8'hc1 == r_count_93_io_out ? io_r_193_b : _GEN_19092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19094 = 8'hc2 == r_count_93_io_out ? io_r_194_b : _GEN_19093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19095 = 8'hc3 == r_count_93_io_out ? io_r_195_b : _GEN_19094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19096 = 8'hc4 == r_count_93_io_out ? io_r_196_b : _GEN_19095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19097 = 8'hc5 == r_count_93_io_out ? io_r_197_b : _GEN_19096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19098 = 8'hc6 == r_count_93_io_out ? io_r_198_b : _GEN_19097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19101 = 8'h1 == r_count_94_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19102 = 8'h2 == r_count_94_io_out ? io_r_2_b : _GEN_19101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19103 = 8'h3 == r_count_94_io_out ? io_r_3_b : _GEN_19102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19104 = 8'h4 == r_count_94_io_out ? io_r_4_b : _GEN_19103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19105 = 8'h5 == r_count_94_io_out ? io_r_5_b : _GEN_19104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19106 = 8'h6 == r_count_94_io_out ? io_r_6_b : _GEN_19105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19107 = 8'h7 == r_count_94_io_out ? io_r_7_b : _GEN_19106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19108 = 8'h8 == r_count_94_io_out ? io_r_8_b : _GEN_19107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19109 = 8'h9 == r_count_94_io_out ? io_r_9_b : _GEN_19108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19110 = 8'ha == r_count_94_io_out ? io_r_10_b : _GEN_19109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19111 = 8'hb == r_count_94_io_out ? io_r_11_b : _GEN_19110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19112 = 8'hc == r_count_94_io_out ? io_r_12_b : _GEN_19111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19113 = 8'hd == r_count_94_io_out ? io_r_13_b : _GEN_19112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19114 = 8'he == r_count_94_io_out ? io_r_14_b : _GEN_19113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19115 = 8'hf == r_count_94_io_out ? io_r_15_b : _GEN_19114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19116 = 8'h10 == r_count_94_io_out ? io_r_16_b : _GEN_19115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19117 = 8'h11 == r_count_94_io_out ? io_r_17_b : _GEN_19116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19118 = 8'h12 == r_count_94_io_out ? io_r_18_b : _GEN_19117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19119 = 8'h13 == r_count_94_io_out ? io_r_19_b : _GEN_19118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19120 = 8'h14 == r_count_94_io_out ? io_r_20_b : _GEN_19119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19121 = 8'h15 == r_count_94_io_out ? io_r_21_b : _GEN_19120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19122 = 8'h16 == r_count_94_io_out ? io_r_22_b : _GEN_19121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19123 = 8'h17 == r_count_94_io_out ? io_r_23_b : _GEN_19122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19124 = 8'h18 == r_count_94_io_out ? io_r_24_b : _GEN_19123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19125 = 8'h19 == r_count_94_io_out ? io_r_25_b : _GEN_19124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19126 = 8'h1a == r_count_94_io_out ? io_r_26_b : _GEN_19125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19127 = 8'h1b == r_count_94_io_out ? io_r_27_b : _GEN_19126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19128 = 8'h1c == r_count_94_io_out ? io_r_28_b : _GEN_19127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19129 = 8'h1d == r_count_94_io_out ? io_r_29_b : _GEN_19128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19130 = 8'h1e == r_count_94_io_out ? io_r_30_b : _GEN_19129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19131 = 8'h1f == r_count_94_io_out ? io_r_31_b : _GEN_19130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19132 = 8'h20 == r_count_94_io_out ? io_r_32_b : _GEN_19131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19133 = 8'h21 == r_count_94_io_out ? io_r_33_b : _GEN_19132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19134 = 8'h22 == r_count_94_io_out ? io_r_34_b : _GEN_19133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19135 = 8'h23 == r_count_94_io_out ? io_r_35_b : _GEN_19134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19136 = 8'h24 == r_count_94_io_out ? io_r_36_b : _GEN_19135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19137 = 8'h25 == r_count_94_io_out ? io_r_37_b : _GEN_19136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19138 = 8'h26 == r_count_94_io_out ? io_r_38_b : _GEN_19137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19139 = 8'h27 == r_count_94_io_out ? io_r_39_b : _GEN_19138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19140 = 8'h28 == r_count_94_io_out ? io_r_40_b : _GEN_19139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19141 = 8'h29 == r_count_94_io_out ? io_r_41_b : _GEN_19140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19142 = 8'h2a == r_count_94_io_out ? io_r_42_b : _GEN_19141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19143 = 8'h2b == r_count_94_io_out ? io_r_43_b : _GEN_19142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19144 = 8'h2c == r_count_94_io_out ? io_r_44_b : _GEN_19143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19145 = 8'h2d == r_count_94_io_out ? io_r_45_b : _GEN_19144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19146 = 8'h2e == r_count_94_io_out ? io_r_46_b : _GEN_19145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19147 = 8'h2f == r_count_94_io_out ? io_r_47_b : _GEN_19146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19148 = 8'h30 == r_count_94_io_out ? io_r_48_b : _GEN_19147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19149 = 8'h31 == r_count_94_io_out ? io_r_49_b : _GEN_19148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19150 = 8'h32 == r_count_94_io_out ? io_r_50_b : _GEN_19149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19151 = 8'h33 == r_count_94_io_out ? io_r_51_b : _GEN_19150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19152 = 8'h34 == r_count_94_io_out ? io_r_52_b : _GEN_19151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19153 = 8'h35 == r_count_94_io_out ? io_r_53_b : _GEN_19152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19154 = 8'h36 == r_count_94_io_out ? io_r_54_b : _GEN_19153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19155 = 8'h37 == r_count_94_io_out ? io_r_55_b : _GEN_19154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19156 = 8'h38 == r_count_94_io_out ? io_r_56_b : _GEN_19155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19157 = 8'h39 == r_count_94_io_out ? io_r_57_b : _GEN_19156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19158 = 8'h3a == r_count_94_io_out ? io_r_58_b : _GEN_19157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19159 = 8'h3b == r_count_94_io_out ? io_r_59_b : _GEN_19158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19160 = 8'h3c == r_count_94_io_out ? io_r_60_b : _GEN_19159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19161 = 8'h3d == r_count_94_io_out ? io_r_61_b : _GEN_19160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19162 = 8'h3e == r_count_94_io_out ? io_r_62_b : _GEN_19161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19163 = 8'h3f == r_count_94_io_out ? io_r_63_b : _GEN_19162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19164 = 8'h40 == r_count_94_io_out ? io_r_64_b : _GEN_19163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19165 = 8'h41 == r_count_94_io_out ? io_r_65_b : _GEN_19164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19166 = 8'h42 == r_count_94_io_out ? io_r_66_b : _GEN_19165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19167 = 8'h43 == r_count_94_io_out ? io_r_67_b : _GEN_19166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19168 = 8'h44 == r_count_94_io_out ? io_r_68_b : _GEN_19167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19169 = 8'h45 == r_count_94_io_out ? io_r_69_b : _GEN_19168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19170 = 8'h46 == r_count_94_io_out ? io_r_70_b : _GEN_19169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19171 = 8'h47 == r_count_94_io_out ? io_r_71_b : _GEN_19170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19172 = 8'h48 == r_count_94_io_out ? io_r_72_b : _GEN_19171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19173 = 8'h49 == r_count_94_io_out ? io_r_73_b : _GEN_19172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19174 = 8'h4a == r_count_94_io_out ? io_r_74_b : _GEN_19173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19175 = 8'h4b == r_count_94_io_out ? io_r_75_b : _GEN_19174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19176 = 8'h4c == r_count_94_io_out ? io_r_76_b : _GEN_19175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19177 = 8'h4d == r_count_94_io_out ? io_r_77_b : _GEN_19176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19178 = 8'h4e == r_count_94_io_out ? io_r_78_b : _GEN_19177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19179 = 8'h4f == r_count_94_io_out ? io_r_79_b : _GEN_19178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19180 = 8'h50 == r_count_94_io_out ? io_r_80_b : _GEN_19179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19181 = 8'h51 == r_count_94_io_out ? io_r_81_b : _GEN_19180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19182 = 8'h52 == r_count_94_io_out ? io_r_82_b : _GEN_19181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19183 = 8'h53 == r_count_94_io_out ? io_r_83_b : _GEN_19182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19184 = 8'h54 == r_count_94_io_out ? io_r_84_b : _GEN_19183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19185 = 8'h55 == r_count_94_io_out ? io_r_85_b : _GEN_19184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19186 = 8'h56 == r_count_94_io_out ? io_r_86_b : _GEN_19185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19187 = 8'h57 == r_count_94_io_out ? io_r_87_b : _GEN_19186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19188 = 8'h58 == r_count_94_io_out ? io_r_88_b : _GEN_19187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19189 = 8'h59 == r_count_94_io_out ? io_r_89_b : _GEN_19188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19190 = 8'h5a == r_count_94_io_out ? io_r_90_b : _GEN_19189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19191 = 8'h5b == r_count_94_io_out ? io_r_91_b : _GEN_19190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19192 = 8'h5c == r_count_94_io_out ? io_r_92_b : _GEN_19191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19193 = 8'h5d == r_count_94_io_out ? io_r_93_b : _GEN_19192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19194 = 8'h5e == r_count_94_io_out ? io_r_94_b : _GEN_19193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19195 = 8'h5f == r_count_94_io_out ? io_r_95_b : _GEN_19194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19196 = 8'h60 == r_count_94_io_out ? io_r_96_b : _GEN_19195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19197 = 8'h61 == r_count_94_io_out ? io_r_97_b : _GEN_19196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19198 = 8'h62 == r_count_94_io_out ? io_r_98_b : _GEN_19197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19199 = 8'h63 == r_count_94_io_out ? io_r_99_b : _GEN_19198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19200 = 8'h64 == r_count_94_io_out ? io_r_100_b : _GEN_19199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19201 = 8'h65 == r_count_94_io_out ? io_r_101_b : _GEN_19200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19202 = 8'h66 == r_count_94_io_out ? io_r_102_b : _GEN_19201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19203 = 8'h67 == r_count_94_io_out ? io_r_103_b : _GEN_19202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19204 = 8'h68 == r_count_94_io_out ? io_r_104_b : _GEN_19203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19205 = 8'h69 == r_count_94_io_out ? io_r_105_b : _GEN_19204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19206 = 8'h6a == r_count_94_io_out ? io_r_106_b : _GEN_19205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19207 = 8'h6b == r_count_94_io_out ? io_r_107_b : _GEN_19206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19208 = 8'h6c == r_count_94_io_out ? io_r_108_b : _GEN_19207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19209 = 8'h6d == r_count_94_io_out ? io_r_109_b : _GEN_19208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19210 = 8'h6e == r_count_94_io_out ? io_r_110_b : _GEN_19209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19211 = 8'h6f == r_count_94_io_out ? io_r_111_b : _GEN_19210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19212 = 8'h70 == r_count_94_io_out ? io_r_112_b : _GEN_19211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19213 = 8'h71 == r_count_94_io_out ? io_r_113_b : _GEN_19212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19214 = 8'h72 == r_count_94_io_out ? io_r_114_b : _GEN_19213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19215 = 8'h73 == r_count_94_io_out ? io_r_115_b : _GEN_19214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19216 = 8'h74 == r_count_94_io_out ? io_r_116_b : _GEN_19215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19217 = 8'h75 == r_count_94_io_out ? io_r_117_b : _GEN_19216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19218 = 8'h76 == r_count_94_io_out ? io_r_118_b : _GEN_19217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19219 = 8'h77 == r_count_94_io_out ? io_r_119_b : _GEN_19218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19220 = 8'h78 == r_count_94_io_out ? io_r_120_b : _GEN_19219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19221 = 8'h79 == r_count_94_io_out ? io_r_121_b : _GEN_19220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19222 = 8'h7a == r_count_94_io_out ? io_r_122_b : _GEN_19221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19223 = 8'h7b == r_count_94_io_out ? io_r_123_b : _GEN_19222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19224 = 8'h7c == r_count_94_io_out ? io_r_124_b : _GEN_19223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19225 = 8'h7d == r_count_94_io_out ? io_r_125_b : _GEN_19224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19226 = 8'h7e == r_count_94_io_out ? io_r_126_b : _GEN_19225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19227 = 8'h7f == r_count_94_io_out ? io_r_127_b : _GEN_19226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19228 = 8'h80 == r_count_94_io_out ? io_r_128_b : _GEN_19227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19229 = 8'h81 == r_count_94_io_out ? io_r_129_b : _GEN_19228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19230 = 8'h82 == r_count_94_io_out ? io_r_130_b : _GEN_19229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19231 = 8'h83 == r_count_94_io_out ? io_r_131_b : _GEN_19230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19232 = 8'h84 == r_count_94_io_out ? io_r_132_b : _GEN_19231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19233 = 8'h85 == r_count_94_io_out ? io_r_133_b : _GEN_19232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19234 = 8'h86 == r_count_94_io_out ? io_r_134_b : _GEN_19233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19235 = 8'h87 == r_count_94_io_out ? io_r_135_b : _GEN_19234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19236 = 8'h88 == r_count_94_io_out ? io_r_136_b : _GEN_19235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19237 = 8'h89 == r_count_94_io_out ? io_r_137_b : _GEN_19236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19238 = 8'h8a == r_count_94_io_out ? io_r_138_b : _GEN_19237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19239 = 8'h8b == r_count_94_io_out ? io_r_139_b : _GEN_19238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19240 = 8'h8c == r_count_94_io_out ? io_r_140_b : _GEN_19239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19241 = 8'h8d == r_count_94_io_out ? io_r_141_b : _GEN_19240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19242 = 8'h8e == r_count_94_io_out ? io_r_142_b : _GEN_19241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19243 = 8'h8f == r_count_94_io_out ? io_r_143_b : _GEN_19242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19244 = 8'h90 == r_count_94_io_out ? io_r_144_b : _GEN_19243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19245 = 8'h91 == r_count_94_io_out ? io_r_145_b : _GEN_19244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19246 = 8'h92 == r_count_94_io_out ? io_r_146_b : _GEN_19245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19247 = 8'h93 == r_count_94_io_out ? io_r_147_b : _GEN_19246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19248 = 8'h94 == r_count_94_io_out ? io_r_148_b : _GEN_19247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19249 = 8'h95 == r_count_94_io_out ? io_r_149_b : _GEN_19248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19250 = 8'h96 == r_count_94_io_out ? io_r_150_b : _GEN_19249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19251 = 8'h97 == r_count_94_io_out ? io_r_151_b : _GEN_19250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19252 = 8'h98 == r_count_94_io_out ? io_r_152_b : _GEN_19251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19253 = 8'h99 == r_count_94_io_out ? io_r_153_b : _GEN_19252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19254 = 8'h9a == r_count_94_io_out ? io_r_154_b : _GEN_19253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19255 = 8'h9b == r_count_94_io_out ? io_r_155_b : _GEN_19254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19256 = 8'h9c == r_count_94_io_out ? io_r_156_b : _GEN_19255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19257 = 8'h9d == r_count_94_io_out ? io_r_157_b : _GEN_19256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19258 = 8'h9e == r_count_94_io_out ? io_r_158_b : _GEN_19257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19259 = 8'h9f == r_count_94_io_out ? io_r_159_b : _GEN_19258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19260 = 8'ha0 == r_count_94_io_out ? io_r_160_b : _GEN_19259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19261 = 8'ha1 == r_count_94_io_out ? io_r_161_b : _GEN_19260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19262 = 8'ha2 == r_count_94_io_out ? io_r_162_b : _GEN_19261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19263 = 8'ha3 == r_count_94_io_out ? io_r_163_b : _GEN_19262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19264 = 8'ha4 == r_count_94_io_out ? io_r_164_b : _GEN_19263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19265 = 8'ha5 == r_count_94_io_out ? io_r_165_b : _GEN_19264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19266 = 8'ha6 == r_count_94_io_out ? io_r_166_b : _GEN_19265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19267 = 8'ha7 == r_count_94_io_out ? io_r_167_b : _GEN_19266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19268 = 8'ha8 == r_count_94_io_out ? io_r_168_b : _GEN_19267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19269 = 8'ha9 == r_count_94_io_out ? io_r_169_b : _GEN_19268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19270 = 8'haa == r_count_94_io_out ? io_r_170_b : _GEN_19269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19271 = 8'hab == r_count_94_io_out ? io_r_171_b : _GEN_19270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19272 = 8'hac == r_count_94_io_out ? io_r_172_b : _GEN_19271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19273 = 8'had == r_count_94_io_out ? io_r_173_b : _GEN_19272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19274 = 8'hae == r_count_94_io_out ? io_r_174_b : _GEN_19273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19275 = 8'haf == r_count_94_io_out ? io_r_175_b : _GEN_19274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19276 = 8'hb0 == r_count_94_io_out ? io_r_176_b : _GEN_19275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19277 = 8'hb1 == r_count_94_io_out ? io_r_177_b : _GEN_19276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19278 = 8'hb2 == r_count_94_io_out ? io_r_178_b : _GEN_19277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19279 = 8'hb3 == r_count_94_io_out ? io_r_179_b : _GEN_19278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19280 = 8'hb4 == r_count_94_io_out ? io_r_180_b : _GEN_19279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19281 = 8'hb5 == r_count_94_io_out ? io_r_181_b : _GEN_19280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19282 = 8'hb6 == r_count_94_io_out ? io_r_182_b : _GEN_19281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19283 = 8'hb7 == r_count_94_io_out ? io_r_183_b : _GEN_19282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19284 = 8'hb8 == r_count_94_io_out ? io_r_184_b : _GEN_19283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19285 = 8'hb9 == r_count_94_io_out ? io_r_185_b : _GEN_19284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19286 = 8'hba == r_count_94_io_out ? io_r_186_b : _GEN_19285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19287 = 8'hbb == r_count_94_io_out ? io_r_187_b : _GEN_19286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19288 = 8'hbc == r_count_94_io_out ? io_r_188_b : _GEN_19287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19289 = 8'hbd == r_count_94_io_out ? io_r_189_b : _GEN_19288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19290 = 8'hbe == r_count_94_io_out ? io_r_190_b : _GEN_19289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19291 = 8'hbf == r_count_94_io_out ? io_r_191_b : _GEN_19290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19292 = 8'hc0 == r_count_94_io_out ? io_r_192_b : _GEN_19291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19293 = 8'hc1 == r_count_94_io_out ? io_r_193_b : _GEN_19292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19294 = 8'hc2 == r_count_94_io_out ? io_r_194_b : _GEN_19293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19295 = 8'hc3 == r_count_94_io_out ? io_r_195_b : _GEN_19294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19296 = 8'hc4 == r_count_94_io_out ? io_r_196_b : _GEN_19295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19297 = 8'hc5 == r_count_94_io_out ? io_r_197_b : _GEN_19296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19298 = 8'hc6 == r_count_94_io_out ? io_r_198_b : _GEN_19297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19301 = 8'h1 == r_count_95_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19302 = 8'h2 == r_count_95_io_out ? io_r_2_b : _GEN_19301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19303 = 8'h3 == r_count_95_io_out ? io_r_3_b : _GEN_19302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19304 = 8'h4 == r_count_95_io_out ? io_r_4_b : _GEN_19303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19305 = 8'h5 == r_count_95_io_out ? io_r_5_b : _GEN_19304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19306 = 8'h6 == r_count_95_io_out ? io_r_6_b : _GEN_19305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19307 = 8'h7 == r_count_95_io_out ? io_r_7_b : _GEN_19306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19308 = 8'h8 == r_count_95_io_out ? io_r_8_b : _GEN_19307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19309 = 8'h9 == r_count_95_io_out ? io_r_9_b : _GEN_19308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19310 = 8'ha == r_count_95_io_out ? io_r_10_b : _GEN_19309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19311 = 8'hb == r_count_95_io_out ? io_r_11_b : _GEN_19310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19312 = 8'hc == r_count_95_io_out ? io_r_12_b : _GEN_19311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19313 = 8'hd == r_count_95_io_out ? io_r_13_b : _GEN_19312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19314 = 8'he == r_count_95_io_out ? io_r_14_b : _GEN_19313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19315 = 8'hf == r_count_95_io_out ? io_r_15_b : _GEN_19314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19316 = 8'h10 == r_count_95_io_out ? io_r_16_b : _GEN_19315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19317 = 8'h11 == r_count_95_io_out ? io_r_17_b : _GEN_19316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19318 = 8'h12 == r_count_95_io_out ? io_r_18_b : _GEN_19317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19319 = 8'h13 == r_count_95_io_out ? io_r_19_b : _GEN_19318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19320 = 8'h14 == r_count_95_io_out ? io_r_20_b : _GEN_19319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19321 = 8'h15 == r_count_95_io_out ? io_r_21_b : _GEN_19320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19322 = 8'h16 == r_count_95_io_out ? io_r_22_b : _GEN_19321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19323 = 8'h17 == r_count_95_io_out ? io_r_23_b : _GEN_19322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19324 = 8'h18 == r_count_95_io_out ? io_r_24_b : _GEN_19323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19325 = 8'h19 == r_count_95_io_out ? io_r_25_b : _GEN_19324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19326 = 8'h1a == r_count_95_io_out ? io_r_26_b : _GEN_19325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19327 = 8'h1b == r_count_95_io_out ? io_r_27_b : _GEN_19326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19328 = 8'h1c == r_count_95_io_out ? io_r_28_b : _GEN_19327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19329 = 8'h1d == r_count_95_io_out ? io_r_29_b : _GEN_19328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19330 = 8'h1e == r_count_95_io_out ? io_r_30_b : _GEN_19329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19331 = 8'h1f == r_count_95_io_out ? io_r_31_b : _GEN_19330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19332 = 8'h20 == r_count_95_io_out ? io_r_32_b : _GEN_19331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19333 = 8'h21 == r_count_95_io_out ? io_r_33_b : _GEN_19332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19334 = 8'h22 == r_count_95_io_out ? io_r_34_b : _GEN_19333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19335 = 8'h23 == r_count_95_io_out ? io_r_35_b : _GEN_19334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19336 = 8'h24 == r_count_95_io_out ? io_r_36_b : _GEN_19335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19337 = 8'h25 == r_count_95_io_out ? io_r_37_b : _GEN_19336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19338 = 8'h26 == r_count_95_io_out ? io_r_38_b : _GEN_19337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19339 = 8'h27 == r_count_95_io_out ? io_r_39_b : _GEN_19338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19340 = 8'h28 == r_count_95_io_out ? io_r_40_b : _GEN_19339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19341 = 8'h29 == r_count_95_io_out ? io_r_41_b : _GEN_19340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19342 = 8'h2a == r_count_95_io_out ? io_r_42_b : _GEN_19341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19343 = 8'h2b == r_count_95_io_out ? io_r_43_b : _GEN_19342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19344 = 8'h2c == r_count_95_io_out ? io_r_44_b : _GEN_19343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19345 = 8'h2d == r_count_95_io_out ? io_r_45_b : _GEN_19344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19346 = 8'h2e == r_count_95_io_out ? io_r_46_b : _GEN_19345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19347 = 8'h2f == r_count_95_io_out ? io_r_47_b : _GEN_19346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19348 = 8'h30 == r_count_95_io_out ? io_r_48_b : _GEN_19347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19349 = 8'h31 == r_count_95_io_out ? io_r_49_b : _GEN_19348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19350 = 8'h32 == r_count_95_io_out ? io_r_50_b : _GEN_19349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19351 = 8'h33 == r_count_95_io_out ? io_r_51_b : _GEN_19350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19352 = 8'h34 == r_count_95_io_out ? io_r_52_b : _GEN_19351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19353 = 8'h35 == r_count_95_io_out ? io_r_53_b : _GEN_19352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19354 = 8'h36 == r_count_95_io_out ? io_r_54_b : _GEN_19353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19355 = 8'h37 == r_count_95_io_out ? io_r_55_b : _GEN_19354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19356 = 8'h38 == r_count_95_io_out ? io_r_56_b : _GEN_19355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19357 = 8'h39 == r_count_95_io_out ? io_r_57_b : _GEN_19356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19358 = 8'h3a == r_count_95_io_out ? io_r_58_b : _GEN_19357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19359 = 8'h3b == r_count_95_io_out ? io_r_59_b : _GEN_19358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19360 = 8'h3c == r_count_95_io_out ? io_r_60_b : _GEN_19359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19361 = 8'h3d == r_count_95_io_out ? io_r_61_b : _GEN_19360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19362 = 8'h3e == r_count_95_io_out ? io_r_62_b : _GEN_19361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19363 = 8'h3f == r_count_95_io_out ? io_r_63_b : _GEN_19362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19364 = 8'h40 == r_count_95_io_out ? io_r_64_b : _GEN_19363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19365 = 8'h41 == r_count_95_io_out ? io_r_65_b : _GEN_19364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19366 = 8'h42 == r_count_95_io_out ? io_r_66_b : _GEN_19365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19367 = 8'h43 == r_count_95_io_out ? io_r_67_b : _GEN_19366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19368 = 8'h44 == r_count_95_io_out ? io_r_68_b : _GEN_19367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19369 = 8'h45 == r_count_95_io_out ? io_r_69_b : _GEN_19368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19370 = 8'h46 == r_count_95_io_out ? io_r_70_b : _GEN_19369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19371 = 8'h47 == r_count_95_io_out ? io_r_71_b : _GEN_19370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19372 = 8'h48 == r_count_95_io_out ? io_r_72_b : _GEN_19371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19373 = 8'h49 == r_count_95_io_out ? io_r_73_b : _GEN_19372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19374 = 8'h4a == r_count_95_io_out ? io_r_74_b : _GEN_19373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19375 = 8'h4b == r_count_95_io_out ? io_r_75_b : _GEN_19374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19376 = 8'h4c == r_count_95_io_out ? io_r_76_b : _GEN_19375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19377 = 8'h4d == r_count_95_io_out ? io_r_77_b : _GEN_19376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19378 = 8'h4e == r_count_95_io_out ? io_r_78_b : _GEN_19377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19379 = 8'h4f == r_count_95_io_out ? io_r_79_b : _GEN_19378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19380 = 8'h50 == r_count_95_io_out ? io_r_80_b : _GEN_19379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19381 = 8'h51 == r_count_95_io_out ? io_r_81_b : _GEN_19380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19382 = 8'h52 == r_count_95_io_out ? io_r_82_b : _GEN_19381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19383 = 8'h53 == r_count_95_io_out ? io_r_83_b : _GEN_19382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19384 = 8'h54 == r_count_95_io_out ? io_r_84_b : _GEN_19383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19385 = 8'h55 == r_count_95_io_out ? io_r_85_b : _GEN_19384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19386 = 8'h56 == r_count_95_io_out ? io_r_86_b : _GEN_19385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19387 = 8'h57 == r_count_95_io_out ? io_r_87_b : _GEN_19386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19388 = 8'h58 == r_count_95_io_out ? io_r_88_b : _GEN_19387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19389 = 8'h59 == r_count_95_io_out ? io_r_89_b : _GEN_19388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19390 = 8'h5a == r_count_95_io_out ? io_r_90_b : _GEN_19389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19391 = 8'h5b == r_count_95_io_out ? io_r_91_b : _GEN_19390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19392 = 8'h5c == r_count_95_io_out ? io_r_92_b : _GEN_19391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19393 = 8'h5d == r_count_95_io_out ? io_r_93_b : _GEN_19392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19394 = 8'h5e == r_count_95_io_out ? io_r_94_b : _GEN_19393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19395 = 8'h5f == r_count_95_io_out ? io_r_95_b : _GEN_19394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19396 = 8'h60 == r_count_95_io_out ? io_r_96_b : _GEN_19395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19397 = 8'h61 == r_count_95_io_out ? io_r_97_b : _GEN_19396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19398 = 8'h62 == r_count_95_io_out ? io_r_98_b : _GEN_19397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19399 = 8'h63 == r_count_95_io_out ? io_r_99_b : _GEN_19398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19400 = 8'h64 == r_count_95_io_out ? io_r_100_b : _GEN_19399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19401 = 8'h65 == r_count_95_io_out ? io_r_101_b : _GEN_19400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19402 = 8'h66 == r_count_95_io_out ? io_r_102_b : _GEN_19401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19403 = 8'h67 == r_count_95_io_out ? io_r_103_b : _GEN_19402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19404 = 8'h68 == r_count_95_io_out ? io_r_104_b : _GEN_19403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19405 = 8'h69 == r_count_95_io_out ? io_r_105_b : _GEN_19404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19406 = 8'h6a == r_count_95_io_out ? io_r_106_b : _GEN_19405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19407 = 8'h6b == r_count_95_io_out ? io_r_107_b : _GEN_19406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19408 = 8'h6c == r_count_95_io_out ? io_r_108_b : _GEN_19407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19409 = 8'h6d == r_count_95_io_out ? io_r_109_b : _GEN_19408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19410 = 8'h6e == r_count_95_io_out ? io_r_110_b : _GEN_19409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19411 = 8'h6f == r_count_95_io_out ? io_r_111_b : _GEN_19410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19412 = 8'h70 == r_count_95_io_out ? io_r_112_b : _GEN_19411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19413 = 8'h71 == r_count_95_io_out ? io_r_113_b : _GEN_19412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19414 = 8'h72 == r_count_95_io_out ? io_r_114_b : _GEN_19413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19415 = 8'h73 == r_count_95_io_out ? io_r_115_b : _GEN_19414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19416 = 8'h74 == r_count_95_io_out ? io_r_116_b : _GEN_19415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19417 = 8'h75 == r_count_95_io_out ? io_r_117_b : _GEN_19416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19418 = 8'h76 == r_count_95_io_out ? io_r_118_b : _GEN_19417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19419 = 8'h77 == r_count_95_io_out ? io_r_119_b : _GEN_19418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19420 = 8'h78 == r_count_95_io_out ? io_r_120_b : _GEN_19419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19421 = 8'h79 == r_count_95_io_out ? io_r_121_b : _GEN_19420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19422 = 8'h7a == r_count_95_io_out ? io_r_122_b : _GEN_19421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19423 = 8'h7b == r_count_95_io_out ? io_r_123_b : _GEN_19422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19424 = 8'h7c == r_count_95_io_out ? io_r_124_b : _GEN_19423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19425 = 8'h7d == r_count_95_io_out ? io_r_125_b : _GEN_19424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19426 = 8'h7e == r_count_95_io_out ? io_r_126_b : _GEN_19425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19427 = 8'h7f == r_count_95_io_out ? io_r_127_b : _GEN_19426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19428 = 8'h80 == r_count_95_io_out ? io_r_128_b : _GEN_19427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19429 = 8'h81 == r_count_95_io_out ? io_r_129_b : _GEN_19428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19430 = 8'h82 == r_count_95_io_out ? io_r_130_b : _GEN_19429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19431 = 8'h83 == r_count_95_io_out ? io_r_131_b : _GEN_19430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19432 = 8'h84 == r_count_95_io_out ? io_r_132_b : _GEN_19431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19433 = 8'h85 == r_count_95_io_out ? io_r_133_b : _GEN_19432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19434 = 8'h86 == r_count_95_io_out ? io_r_134_b : _GEN_19433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19435 = 8'h87 == r_count_95_io_out ? io_r_135_b : _GEN_19434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19436 = 8'h88 == r_count_95_io_out ? io_r_136_b : _GEN_19435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19437 = 8'h89 == r_count_95_io_out ? io_r_137_b : _GEN_19436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19438 = 8'h8a == r_count_95_io_out ? io_r_138_b : _GEN_19437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19439 = 8'h8b == r_count_95_io_out ? io_r_139_b : _GEN_19438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19440 = 8'h8c == r_count_95_io_out ? io_r_140_b : _GEN_19439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19441 = 8'h8d == r_count_95_io_out ? io_r_141_b : _GEN_19440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19442 = 8'h8e == r_count_95_io_out ? io_r_142_b : _GEN_19441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19443 = 8'h8f == r_count_95_io_out ? io_r_143_b : _GEN_19442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19444 = 8'h90 == r_count_95_io_out ? io_r_144_b : _GEN_19443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19445 = 8'h91 == r_count_95_io_out ? io_r_145_b : _GEN_19444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19446 = 8'h92 == r_count_95_io_out ? io_r_146_b : _GEN_19445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19447 = 8'h93 == r_count_95_io_out ? io_r_147_b : _GEN_19446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19448 = 8'h94 == r_count_95_io_out ? io_r_148_b : _GEN_19447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19449 = 8'h95 == r_count_95_io_out ? io_r_149_b : _GEN_19448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19450 = 8'h96 == r_count_95_io_out ? io_r_150_b : _GEN_19449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19451 = 8'h97 == r_count_95_io_out ? io_r_151_b : _GEN_19450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19452 = 8'h98 == r_count_95_io_out ? io_r_152_b : _GEN_19451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19453 = 8'h99 == r_count_95_io_out ? io_r_153_b : _GEN_19452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19454 = 8'h9a == r_count_95_io_out ? io_r_154_b : _GEN_19453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19455 = 8'h9b == r_count_95_io_out ? io_r_155_b : _GEN_19454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19456 = 8'h9c == r_count_95_io_out ? io_r_156_b : _GEN_19455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19457 = 8'h9d == r_count_95_io_out ? io_r_157_b : _GEN_19456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19458 = 8'h9e == r_count_95_io_out ? io_r_158_b : _GEN_19457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19459 = 8'h9f == r_count_95_io_out ? io_r_159_b : _GEN_19458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19460 = 8'ha0 == r_count_95_io_out ? io_r_160_b : _GEN_19459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19461 = 8'ha1 == r_count_95_io_out ? io_r_161_b : _GEN_19460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19462 = 8'ha2 == r_count_95_io_out ? io_r_162_b : _GEN_19461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19463 = 8'ha3 == r_count_95_io_out ? io_r_163_b : _GEN_19462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19464 = 8'ha4 == r_count_95_io_out ? io_r_164_b : _GEN_19463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19465 = 8'ha5 == r_count_95_io_out ? io_r_165_b : _GEN_19464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19466 = 8'ha6 == r_count_95_io_out ? io_r_166_b : _GEN_19465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19467 = 8'ha7 == r_count_95_io_out ? io_r_167_b : _GEN_19466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19468 = 8'ha8 == r_count_95_io_out ? io_r_168_b : _GEN_19467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19469 = 8'ha9 == r_count_95_io_out ? io_r_169_b : _GEN_19468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19470 = 8'haa == r_count_95_io_out ? io_r_170_b : _GEN_19469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19471 = 8'hab == r_count_95_io_out ? io_r_171_b : _GEN_19470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19472 = 8'hac == r_count_95_io_out ? io_r_172_b : _GEN_19471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19473 = 8'had == r_count_95_io_out ? io_r_173_b : _GEN_19472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19474 = 8'hae == r_count_95_io_out ? io_r_174_b : _GEN_19473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19475 = 8'haf == r_count_95_io_out ? io_r_175_b : _GEN_19474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19476 = 8'hb0 == r_count_95_io_out ? io_r_176_b : _GEN_19475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19477 = 8'hb1 == r_count_95_io_out ? io_r_177_b : _GEN_19476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19478 = 8'hb2 == r_count_95_io_out ? io_r_178_b : _GEN_19477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19479 = 8'hb3 == r_count_95_io_out ? io_r_179_b : _GEN_19478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19480 = 8'hb4 == r_count_95_io_out ? io_r_180_b : _GEN_19479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19481 = 8'hb5 == r_count_95_io_out ? io_r_181_b : _GEN_19480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19482 = 8'hb6 == r_count_95_io_out ? io_r_182_b : _GEN_19481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19483 = 8'hb7 == r_count_95_io_out ? io_r_183_b : _GEN_19482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19484 = 8'hb8 == r_count_95_io_out ? io_r_184_b : _GEN_19483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19485 = 8'hb9 == r_count_95_io_out ? io_r_185_b : _GEN_19484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19486 = 8'hba == r_count_95_io_out ? io_r_186_b : _GEN_19485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19487 = 8'hbb == r_count_95_io_out ? io_r_187_b : _GEN_19486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19488 = 8'hbc == r_count_95_io_out ? io_r_188_b : _GEN_19487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19489 = 8'hbd == r_count_95_io_out ? io_r_189_b : _GEN_19488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19490 = 8'hbe == r_count_95_io_out ? io_r_190_b : _GEN_19489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19491 = 8'hbf == r_count_95_io_out ? io_r_191_b : _GEN_19490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19492 = 8'hc0 == r_count_95_io_out ? io_r_192_b : _GEN_19491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19493 = 8'hc1 == r_count_95_io_out ? io_r_193_b : _GEN_19492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19494 = 8'hc2 == r_count_95_io_out ? io_r_194_b : _GEN_19493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19495 = 8'hc3 == r_count_95_io_out ? io_r_195_b : _GEN_19494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19496 = 8'hc4 == r_count_95_io_out ? io_r_196_b : _GEN_19495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19497 = 8'hc5 == r_count_95_io_out ? io_r_197_b : _GEN_19496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19498 = 8'hc6 == r_count_95_io_out ? io_r_198_b : _GEN_19497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19501 = 8'h1 == r_count_96_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19502 = 8'h2 == r_count_96_io_out ? io_r_2_b : _GEN_19501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19503 = 8'h3 == r_count_96_io_out ? io_r_3_b : _GEN_19502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19504 = 8'h4 == r_count_96_io_out ? io_r_4_b : _GEN_19503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19505 = 8'h5 == r_count_96_io_out ? io_r_5_b : _GEN_19504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19506 = 8'h6 == r_count_96_io_out ? io_r_6_b : _GEN_19505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19507 = 8'h7 == r_count_96_io_out ? io_r_7_b : _GEN_19506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19508 = 8'h8 == r_count_96_io_out ? io_r_8_b : _GEN_19507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19509 = 8'h9 == r_count_96_io_out ? io_r_9_b : _GEN_19508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19510 = 8'ha == r_count_96_io_out ? io_r_10_b : _GEN_19509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19511 = 8'hb == r_count_96_io_out ? io_r_11_b : _GEN_19510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19512 = 8'hc == r_count_96_io_out ? io_r_12_b : _GEN_19511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19513 = 8'hd == r_count_96_io_out ? io_r_13_b : _GEN_19512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19514 = 8'he == r_count_96_io_out ? io_r_14_b : _GEN_19513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19515 = 8'hf == r_count_96_io_out ? io_r_15_b : _GEN_19514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19516 = 8'h10 == r_count_96_io_out ? io_r_16_b : _GEN_19515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19517 = 8'h11 == r_count_96_io_out ? io_r_17_b : _GEN_19516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19518 = 8'h12 == r_count_96_io_out ? io_r_18_b : _GEN_19517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19519 = 8'h13 == r_count_96_io_out ? io_r_19_b : _GEN_19518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19520 = 8'h14 == r_count_96_io_out ? io_r_20_b : _GEN_19519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19521 = 8'h15 == r_count_96_io_out ? io_r_21_b : _GEN_19520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19522 = 8'h16 == r_count_96_io_out ? io_r_22_b : _GEN_19521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19523 = 8'h17 == r_count_96_io_out ? io_r_23_b : _GEN_19522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19524 = 8'h18 == r_count_96_io_out ? io_r_24_b : _GEN_19523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19525 = 8'h19 == r_count_96_io_out ? io_r_25_b : _GEN_19524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19526 = 8'h1a == r_count_96_io_out ? io_r_26_b : _GEN_19525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19527 = 8'h1b == r_count_96_io_out ? io_r_27_b : _GEN_19526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19528 = 8'h1c == r_count_96_io_out ? io_r_28_b : _GEN_19527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19529 = 8'h1d == r_count_96_io_out ? io_r_29_b : _GEN_19528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19530 = 8'h1e == r_count_96_io_out ? io_r_30_b : _GEN_19529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19531 = 8'h1f == r_count_96_io_out ? io_r_31_b : _GEN_19530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19532 = 8'h20 == r_count_96_io_out ? io_r_32_b : _GEN_19531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19533 = 8'h21 == r_count_96_io_out ? io_r_33_b : _GEN_19532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19534 = 8'h22 == r_count_96_io_out ? io_r_34_b : _GEN_19533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19535 = 8'h23 == r_count_96_io_out ? io_r_35_b : _GEN_19534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19536 = 8'h24 == r_count_96_io_out ? io_r_36_b : _GEN_19535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19537 = 8'h25 == r_count_96_io_out ? io_r_37_b : _GEN_19536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19538 = 8'h26 == r_count_96_io_out ? io_r_38_b : _GEN_19537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19539 = 8'h27 == r_count_96_io_out ? io_r_39_b : _GEN_19538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19540 = 8'h28 == r_count_96_io_out ? io_r_40_b : _GEN_19539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19541 = 8'h29 == r_count_96_io_out ? io_r_41_b : _GEN_19540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19542 = 8'h2a == r_count_96_io_out ? io_r_42_b : _GEN_19541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19543 = 8'h2b == r_count_96_io_out ? io_r_43_b : _GEN_19542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19544 = 8'h2c == r_count_96_io_out ? io_r_44_b : _GEN_19543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19545 = 8'h2d == r_count_96_io_out ? io_r_45_b : _GEN_19544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19546 = 8'h2e == r_count_96_io_out ? io_r_46_b : _GEN_19545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19547 = 8'h2f == r_count_96_io_out ? io_r_47_b : _GEN_19546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19548 = 8'h30 == r_count_96_io_out ? io_r_48_b : _GEN_19547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19549 = 8'h31 == r_count_96_io_out ? io_r_49_b : _GEN_19548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19550 = 8'h32 == r_count_96_io_out ? io_r_50_b : _GEN_19549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19551 = 8'h33 == r_count_96_io_out ? io_r_51_b : _GEN_19550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19552 = 8'h34 == r_count_96_io_out ? io_r_52_b : _GEN_19551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19553 = 8'h35 == r_count_96_io_out ? io_r_53_b : _GEN_19552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19554 = 8'h36 == r_count_96_io_out ? io_r_54_b : _GEN_19553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19555 = 8'h37 == r_count_96_io_out ? io_r_55_b : _GEN_19554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19556 = 8'h38 == r_count_96_io_out ? io_r_56_b : _GEN_19555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19557 = 8'h39 == r_count_96_io_out ? io_r_57_b : _GEN_19556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19558 = 8'h3a == r_count_96_io_out ? io_r_58_b : _GEN_19557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19559 = 8'h3b == r_count_96_io_out ? io_r_59_b : _GEN_19558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19560 = 8'h3c == r_count_96_io_out ? io_r_60_b : _GEN_19559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19561 = 8'h3d == r_count_96_io_out ? io_r_61_b : _GEN_19560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19562 = 8'h3e == r_count_96_io_out ? io_r_62_b : _GEN_19561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19563 = 8'h3f == r_count_96_io_out ? io_r_63_b : _GEN_19562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19564 = 8'h40 == r_count_96_io_out ? io_r_64_b : _GEN_19563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19565 = 8'h41 == r_count_96_io_out ? io_r_65_b : _GEN_19564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19566 = 8'h42 == r_count_96_io_out ? io_r_66_b : _GEN_19565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19567 = 8'h43 == r_count_96_io_out ? io_r_67_b : _GEN_19566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19568 = 8'h44 == r_count_96_io_out ? io_r_68_b : _GEN_19567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19569 = 8'h45 == r_count_96_io_out ? io_r_69_b : _GEN_19568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19570 = 8'h46 == r_count_96_io_out ? io_r_70_b : _GEN_19569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19571 = 8'h47 == r_count_96_io_out ? io_r_71_b : _GEN_19570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19572 = 8'h48 == r_count_96_io_out ? io_r_72_b : _GEN_19571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19573 = 8'h49 == r_count_96_io_out ? io_r_73_b : _GEN_19572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19574 = 8'h4a == r_count_96_io_out ? io_r_74_b : _GEN_19573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19575 = 8'h4b == r_count_96_io_out ? io_r_75_b : _GEN_19574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19576 = 8'h4c == r_count_96_io_out ? io_r_76_b : _GEN_19575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19577 = 8'h4d == r_count_96_io_out ? io_r_77_b : _GEN_19576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19578 = 8'h4e == r_count_96_io_out ? io_r_78_b : _GEN_19577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19579 = 8'h4f == r_count_96_io_out ? io_r_79_b : _GEN_19578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19580 = 8'h50 == r_count_96_io_out ? io_r_80_b : _GEN_19579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19581 = 8'h51 == r_count_96_io_out ? io_r_81_b : _GEN_19580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19582 = 8'h52 == r_count_96_io_out ? io_r_82_b : _GEN_19581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19583 = 8'h53 == r_count_96_io_out ? io_r_83_b : _GEN_19582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19584 = 8'h54 == r_count_96_io_out ? io_r_84_b : _GEN_19583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19585 = 8'h55 == r_count_96_io_out ? io_r_85_b : _GEN_19584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19586 = 8'h56 == r_count_96_io_out ? io_r_86_b : _GEN_19585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19587 = 8'h57 == r_count_96_io_out ? io_r_87_b : _GEN_19586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19588 = 8'h58 == r_count_96_io_out ? io_r_88_b : _GEN_19587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19589 = 8'h59 == r_count_96_io_out ? io_r_89_b : _GEN_19588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19590 = 8'h5a == r_count_96_io_out ? io_r_90_b : _GEN_19589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19591 = 8'h5b == r_count_96_io_out ? io_r_91_b : _GEN_19590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19592 = 8'h5c == r_count_96_io_out ? io_r_92_b : _GEN_19591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19593 = 8'h5d == r_count_96_io_out ? io_r_93_b : _GEN_19592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19594 = 8'h5e == r_count_96_io_out ? io_r_94_b : _GEN_19593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19595 = 8'h5f == r_count_96_io_out ? io_r_95_b : _GEN_19594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19596 = 8'h60 == r_count_96_io_out ? io_r_96_b : _GEN_19595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19597 = 8'h61 == r_count_96_io_out ? io_r_97_b : _GEN_19596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19598 = 8'h62 == r_count_96_io_out ? io_r_98_b : _GEN_19597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19599 = 8'h63 == r_count_96_io_out ? io_r_99_b : _GEN_19598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19600 = 8'h64 == r_count_96_io_out ? io_r_100_b : _GEN_19599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19601 = 8'h65 == r_count_96_io_out ? io_r_101_b : _GEN_19600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19602 = 8'h66 == r_count_96_io_out ? io_r_102_b : _GEN_19601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19603 = 8'h67 == r_count_96_io_out ? io_r_103_b : _GEN_19602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19604 = 8'h68 == r_count_96_io_out ? io_r_104_b : _GEN_19603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19605 = 8'h69 == r_count_96_io_out ? io_r_105_b : _GEN_19604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19606 = 8'h6a == r_count_96_io_out ? io_r_106_b : _GEN_19605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19607 = 8'h6b == r_count_96_io_out ? io_r_107_b : _GEN_19606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19608 = 8'h6c == r_count_96_io_out ? io_r_108_b : _GEN_19607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19609 = 8'h6d == r_count_96_io_out ? io_r_109_b : _GEN_19608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19610 = 8'h6e == r_count_96_io_out ? io_r_110_b : _GEN_19609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19611 = 8'h6f == r_count_96_io_out ? io_r_111_b : _GEN_19610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19612 = 8'h70 == r_count_96_io_out ? io_r_112_b : _GEN_19611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19613 = 8'h71 == r_count_96_io_out ? io_r_113_b : _GEN_19612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19614 = 8'h72 == r_count_96_io_out ? io_r_114_b : _GEN_19613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19615 = 8'h73 == r_count_96_io_out ? io_r_115_b : _GEN_19614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19616 = 8'h74 == r_count_96_io_out ? io_r_116_b : _GEN_19615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19617 = 8'h75 == r_count_96_io_out ? io_r_117_b : _GEN_19616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19618 = 8'h76 == r_count_96_io_out ? io_r_118_b : _GEN_19617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19619 = 8'h77 == r_count_96_io_out ? io_r_119_b : _GEN_19618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19620 = 8'h78 == r_count_96_io_out ? io_r_120_b : _GEN_19619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19621 = 8'h79 == r_count_96_io_out ? io_r_121_b : _GEN_19620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19622 = 8'h7a == r_count_96_io_out ? io_r_122_b : _GEN_19621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19623 = 8'h7b == r_count_96_io_out ? io_r_123_b : _GEN_19622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19624 = 8'h7c == r_count_96_io_out ? io_r_124_b : _GEN_19623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19625 = 8'h7d == r_count_96_io_out ? io_r_125_b : _GEN_19624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19626 = 8'h7e == r_count_96_io_out ? io_r_126_b : _GEN_19625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19627 = 8'h7f == r_count_96_io_out ? io_r_127_b : _GEN_19626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19628 = 8'h80 == r_count_96_io_out ? io_r_128_b : _GEN_19627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19629 = 8'h81 == r_count_96_io_out ? io_r_129_b : _GEN_19628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19630 = 8'h82 == r_count_96_io_out ? io_r_130_b : _GEN_19629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19631 = 8'h83 == r_count_96_io_out ? io_r_131_b : _GEN_19630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19632 = 8'h84 == r_count_96_io_out ? io_r_132_b : _GEN_19631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19633 = 8'h85 == r_count_96_io_out ? io_r_133_b : _GEN_19632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19634 = 8'h86 == r_count_96_io_out ? io_r_134_b : _GEN_19633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19635 = 8'h87 == r_count_96_io_out ? io_r_135_b : _GEN_19634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19636 = 8'h88 == r_count_96_io_out ? io_r_136_b : _GEN_19635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19637 = 8'h89 == r_count_96_io_out ? io_r_137_b : _GEN_19636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19638 = 8'h8a == r_count_96_io_out ? io_r_138_b : _GEN_19637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19639 = 8'h8b == r_count_96_io_out ? io_r_139_b : _GEN_19638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19640 = 8'h8c == r_count_96_io_out ? io_r_140_b : _GEN_19639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19641 = 8'h8d == r_count_96_io_out ? io_r_141_b : _GEN_19640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19642 = 8'h8e == r_count_96_io_out ? io_r_142_b : _GEN_19641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19643 = 8'h8f == r_count_96_io_out ? io_r_143_b : _GEN_19642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19644 = 8'h90 == r_count_96_io_out ? io_r_144_b : _GEN_19643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19645 = 8'h91 == r_count_96_io_out ? io_r_145_b : _GEN_19644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19646 = 8'h92 == r_count_96_io_out ? io_r_146_b : _GEN_19645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19647 = 8'h93 == r_count_96_io_out ? io_r_147_b : _GEN_19646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19648 = 8'h94 == r_count_96_io_out ? io_r_148_b : _GEN_19647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19649 = 8'h95 == r_count_96_io_out ? io_r_149_b : _GEN_19648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19650 = 8'h96 == r_count_96_io_out ? io_r_150_b : _GEN_19649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19651 = 8'h97 == r_count_96_io_out ? io_r_151_b : _GEN_19650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19652 = 8'h98 == r_count_96_io_out ? io_r_152_b : _GEN_19651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19653 = 8'h99 == r_count_96_io_out ? io_r_153_b : _GEN_19652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19654 = 8'h9a == r_count_96_io_out ? io_r_154_b : _GEN_19653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19655 = 8'h9b == r_count_96_io_out ? io_r_155_b : _GEN_19654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19656 = 8'h9c == r_count_96_io_out ? io_r_156_b : _GEN_19655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19657 = 8'h9d == r_count_96_io_out ? io_r_157_b : _GEN_19656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19658 = 8'h9e == r_count_96_io_out ? io_r_158_b : _GEN_19657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19659 = 8'h9f == r_count_96_io_out ? io_r_159_b : _GEN_19658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19660 = 8'ha0 == r_count_96_io_out ? io_r_160_b : _GEN_19659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19661 = 8'ha1 == r_count_96_io_out ? io_r_161_b : _GEN_19660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19662 = 8'ha2 == r_count_96_io_out ? io_r_162_b : _GEN_19661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19663 = 8'ha3 == r_count_96_io_out ? io_r_163_b : _GEN_19662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19664 = 8'ha4 == r_count_96_io_out ? io_r_164_b : _GEN_19663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19665 = 8'ha5 == r_count_96_io_out ? io_r_165_b : _GEN_19664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19666 = 8'ha6 == r_count_96_io_out ? io_r_166_b : _GEN_19665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19667 = 8'ha7 == r_count_96_io_out ? io_r_167_b : _GEN_19666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19668 = 8'ha8 == r_count_96_io_out ? io_r_168_b : _GEN_19667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19669 = 8'ha9 == r_count_96_io_out ? io_r_169_b : _GEN_19668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19670 = 8'haa == r_count_96_io_out ? io_r_170_b : _GEN_19669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19671 = 8'hab == r_count_96_io_out ? io_r_171_b : _GEN_19670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19672 = 8'hac == r_count_96_io_out ? io_r_172_b : _GEN_19671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19673 = 8'had == r_count_96_io_out ? io_r_173_b : _GEN_19672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19674 = 8'hae == r_count_96_io_out ? io_r_174_b : _GEN_19673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19675 = 8'haf == r_count_96_io_out ? io_r_175_b : _GEN_19674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19676 = 8'hb0 == r_count_96_io_out ? io_r_176_b : _GEN_19675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19677 = 8'hb1 == r_count_96_io_out ? io_r_177_b : _GEN_19676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19678 = 8'hb2 == r_count_96_io_out ? io_r_178_b : _GEN_19677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19679 = 8'hb3 == r_count_96_io_out ? io_r_179_b : _GEN_19678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19680 = 8'hb4 == r_count_96_io_out ? io_r_180_b : _GEN_19679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19681 = 8'hb5 == r_count_96_io_out ? io_r_181_b : _GEN_19680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19682 = 8'hb6 == r_count_96_io_out ? io_r_182_b : _GEN_19681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19683 = 8'hb7 == r_count_96_io_out ? io_r_183_b : _GEN_19682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19684 = 8'hb8 == r_count_96_io_out ? io_r_184_b : _GEN_19683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19685 = 8'hb9 == r_count_96_io_out ? io_r_185_b : _GEN_19684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19686 = 8'hba == r_count_96_io_out ? io_r_186_b : _GEN_19685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19687 = 8'hbb == r_count_96_io_out ? io_r_187_b : _GEN_19686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19688 = 8'hbc == r_count_96_io_out ? io_r_188_b : _GEN_19687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19689 = 8'hbd == r_count_96_io_out ? io_r_189_b : _GEN_19688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19690 = 8'hbe == r_count_96_io_out ? io_r_190_b : _GEN_19689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19691 = 8'hbf == r_count_96_io_out ? io_r_191_b : _GEN_19690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19692 = 8'hc0 == r_count_96_io_out ? io_r_192_b : _GEN_19691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19693 = 8'hc1 == r_count_96_io_out ? io_r_193_b : _GEN_19692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19694 = 8'hc2 == r_count_96_io_out ? io_r_194_b : _GEN_19693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19695 = 8'hc3 == r_count_96_io_out ? io_r_195_b : _GEN_19694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19696 = 8'hc4 == r_count_96_io_out ? io_r_196_b : _GEN_19695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19697 = 8'hc5 == r_count_96_io_out ? io_r_197_b : _GEN_19696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19698 = 8'hc6 == r_count_96_io_out ? io_r_198_b : _GEN_19697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19701 = 8'h1 == r_count_97_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19702 = 8'h2 == r_count_97_io_out ? io_r_2_b : _GEN_19701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19703 = 8'h3 == r_count_97_io_out ? io_r_3_b : _GEN_19702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19704 = 8'h4 == r_count_97_io_out ? io_r_4_b : _GEN_19703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19705 = 8'h5 == r_count_97_io_out ? io_r_5_b : _GEN_19704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19706 = 8'h6 == r_count_97_io_out ? io_r_6_b : _GEN_19705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19707 = 8'h7 == r_count_97_io_out ? io_r_7_b : _GEN_19706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19708 = 8'h8 == r_count_97_io_out ? io_r_8_b : _GEN_19707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19709 = 8'h9 == r_count_97_io_out ? io_r_9_b : _GEN_19708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19710 = 8'ha == r_count_97_io_out ? io_r_10_b : _GEN_19709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19711 = 8'hb == r_count_97_io_out ? io_r_11_b : _GEN_19710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19712 = 8'hc == r_count_97_io_out ? io_r_12_b : _GEN_19711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19713 = 8'hd == r_count_97_io_out ? io_r_13_b : _GEN_19712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19714 = 8'he == r_count_97_io_out ? io_r_14_b : _GEN_19713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19715 = 8'hf == r_count_97_io_out ? io_r_15_b : _GEN_19714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19716 = 8'h10 == r_count_97_io_out ? io_r_16_b : _GEN_19715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19717 = 8'h11 == r_count_97_io_out ? io_r_17_b : _GEN_19716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19718 = 8'h12 == r_count_97_io_out ? io_r_18_b : _GEN_19717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19719 = 8'h13 == r_count_97_io_out ? io_r_19_b : _GEN_19718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19720 = 8'h14 == r_count_97_io_out ? io_r_20_b : _GEN_19719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19721 = 8'h15 == r_count_97_io_out ? io_r_21_b : _GEN_19720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19722 = 8'h16 == r_count_97_io_out ? io_r_22_b : _GEN_19721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19723 = 8'h17 == r_count_97_io_out ? io_r_23_b : _GEN_19722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19724 = 8'h18 == r_count_97_io_out ? io_r_24_b : _GEN_19723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19725 = 8'h19 == r_count_97_io_out ? io_r_25_b : _GEN_19724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19726 = 8'h1a == r_count_97_io_out ? io_r_26_b : _GEN_19725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19727 = 8'h1b == r_count_97_io_out ? io_r_27_b : _GEN_19726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19728 = 8'h1c == r_count_97_io_out ? io_r_28_b : _GEN_19727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19729 = 8'h1d == r_count_97_io_out ? io_r_29_b : _GEN_19728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19730 = 8'h1e == r_count_97_io_out ? io_r_30_b : _GEN_19729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19731 = 8'h1f == r_count_97_io_out ? io_r_31_b : _GEN_19730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19732 = 8'h20 == r_count_97_io_out ? io_r_32_b : _GEN_19731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19733 = 8'h21 == r_count_97_io_out ? io_r_33_b : _GEN_19732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19734 = 8'h22 == r_count_97_io_out ? io_r_34_b : _GEN_19733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19735 = 8'h23 == r_count_97_io_out ? io_r_35_b : _GEN_19734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19736 = 8'h24 == r_count_97_io_out ? io_r_36_b : _GEN_19735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19737 = 8'h25 == r_count_97_io_out ? io_r_37_b : _GEN_19736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19738 = 8'h26 == r_count_97_io_out ? io_r_38_b : _GEN_19737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19739 = 8'h27 == r_count_97_io_out ? io_r_39_b : _GEN_19738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19740 = 8'h28 == r_count_97_io_out ? io_r_40_b : _GEN_19739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19741 = 8'h29 == r_count_97_io_out ? io_r_41_b : _GEN_19740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19742 = 8'h2a == r_count_97_io_out ? io_r_42_b : _GEN_19741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19743 = 8'h2b == r_count_97_io_out ? io_r_43_b : _GEN_19742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19744 = 8'h2c == r_count_97_io_out ? io_r_44_b : _GEN_19743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19745 = 8'h2d == r_count_97_io_out ? io_r_45_b : _GEN_19744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19746 = 8'h2e == r_count_97_io_out ? io_r_46_b : _GEN_19745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19747 = 8'h2f == r_count_97_io_out ? io_r_47_b : _GEN_19746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19748 = 8'h30 == r_count_97_io_out ? io_r_48_b : _GEN_19747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19749 = 8'h31 == r_count_97_io_out ? io_r_49_b : _GEN_19748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19750 = 8'h32 == r_count_97_io_out ? io_r_50_b : _GEN_19749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19751 = 8'h33 == r_count_97_io_out ? io_r_51_b : _GEN_19750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19752 = 8'h34 == r_count_97_io_out ? io_r_52_b : _GEN_19751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19753 = 8'h35 == r_count_97_io_out ? io_r_53_b : _GEN_19752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19754 = 8'h36 == r_count_97_io_out ? io_r_54_b : _GEN_19753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19755 = 8'h37 == r_count_97_io_out ? io_r_55_b : _GEN_19754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19756 = 8'h38 == r_count_97_io_out ? io_r_56_b : _GEN_19755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19757 = 8'h39 == r_count_97_io_out ? io_r_57_b : _GEN_19756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19758 = 8'h3a == r_count_97_io_out ? io_r_58_b : _GEN_19757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19759 = 8'h3b == r_count_97_io_out ? io_r_59_b : _GEN_19758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19760 = 8'h3c == r_count_97_io_out ? io_r_60_b : _GEN_19759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19761 = 8'h3d == r_count_97_io_out ? io_r_61_b : _GEN_19760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19762 = 8'h3e == r_count_97_io_out ? io_r_62_b : _GEN_19761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19763 = 8'h3f == r_count_97_io_out ? io_r_63_b : _GEN_19762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19764 = 8'h40 == r_count_97_io_out ? io_r_64_b : _GEN_19763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19765 = 8'h41 == r_count_97_io_out ? io_r_65_b : _GEN_19764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19766 = 8'h42 == r_count_97_io_out ? io_r_66_b : _GEN_19765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19767 = 8'h43 == r_count_97_io_out ? io_r_67_b : _GEN_19766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19768 = 8'h44 == r_count_97_io_out ? io_r_68_b : _GEN_19767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19769 = 8'h45 == r_count_97_io_out ? io_r_69_b : _GEN_19768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19770 = 8'h46 == r_count_97_io_out ? io_r_70_b : _GEN_19769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19771 = 8'h47 == r_count_97_io_out ? io_r_71_b : _GEN_19770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19772 = 8'h48 == r_count_97_io_out ? io_r_72_b : _GEN_19771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19773 = 8'h49 == r_count_97_io_out ? io_r_73_b : _GEN_19772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19774 = 8'h4a == r_count_97_io_out ? io_r_74_b : _GEN_19773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19775 = 8'h4b == r_count_97_io_out ? io_r_75_b : _GEN_19774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19776 = 8'h4c == r_count_97_io_out ? io_r_76_b : _GEN_19775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19777 = 8'h4d == r_count_97_io_out ? io_r_77_b : _GEN_19776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19778 = 8'h4e == r_count_97_io_out ? io_r_78_b : _GEN_19777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19779 = 8'h4f == r_count_97_io_out ? io_r_79_b : _GEN_19778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19780 = 8'h50 == r_count_97_io_out ? io_r_80_b : _GEN_19779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19781 = 8'h51 == r_count_97_io_out ? io_r_81_b : _GEN_19780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19782 = 8'h52 == r_count_97_io_out ? io_r_82_b : _GEN_19781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19783 = 8'h53 == r_count_97_io_out ? io_r_83_b : _GEN_19782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19784 = 8'h54 == r_count_97_io_out ? io_r_84_b : _GEN_19783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19785 = 8'h55 == r_count_97_io_out ? io_r_85_b : _GEN_19784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19786 = 8'h56 == r_count_97_io_out ? io_r_86_b : _GEN_19785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19787 = 8'h57 == r_count_97_io_out ? io_r_87_b : _GEN_19786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19788 = 8'h58 == r_count_97_io_out ? io_r_88_b : _GEN_19787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19789 = 8'h59 == r_count_97_io_out ? io_r_89_b : _GEN_19788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19790 = 8'h5a == r_count_97_io_out ? io_r_90_b : _GEN_19789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19791 = 8'h5b == r_count_97_io_out ? io_r_91_b : _GEN_19790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19792 = 8'h5c == r_count_97_io_out ? io_r_92_b : _GEN_19791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19793 = 8'h5d == r_count_97_io_out ? io_r_93_b : _GEN_19792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19794 = 8'h5e == r_count_97_io_out ? io_r_94_b : _GEN_19793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19795 = 8'h5f == r_count_97_io_out ? io_r_95_b : _GEN_19794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19796 = 8'h60 == r_count_97_io_out ? io_r_96_b : _GEN_19795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19797 = 8'h61 == r_count_97_io_out ? io_r_97_b : _GEN_19796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19798 = 8'h62 == r_count_97_io_out ? io_r_98_b : _GEN_19797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19799 = 8'h63 == r_count_97_io_out ? io_r_99_b : _GEN_19798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19800 = 8'h64 == r_count_97_io_out ? io_r_100_b : _GEN_19799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19801 = 8'h65 == r_count_97_io_out ? io_r_101_b : _GEN_19800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19802 = 8'h66 == r_count_97_io_out ? io_r_102_b : _GEN_19801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19803 = 8'h67 == r_count_97_io_out ? io_r_103_b : _GEN_19802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19804 = 8'h68 == r_count_97_io_out ? io_r_104_b : _GEN_19803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19805 = 8'h69 == r_count_97_io_out ? io_r_105_b : _GEN_19804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19806 = 8'h6a == r_count_97_io_out ? io_r_106_b : _GEN_19805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19807 = 8'h6b == r_count_97_io_out ? io_r_107_b : _GEN_19806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19808 = 8'h6c == r_count_97_io_out ? io_r_108_b : _GEN_19807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19809 = 8'h6d == r_count_97_io_out ? io_r_109_b : _GEN_19808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19810 = 8'h6e == r_count_97_io_out ? io_r_110_b : _GEN_19809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19811 = 8'h6f == r_count_97_io_out ? io_r_111_b : _GEN_19810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19812 = 8'h70 == r_count_97_io_out ? io_r_112_b : _GEN_19811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19813 = 8'h71 == r_count_97_io_out ? io_r_113_b : _GEN_19812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19814 = 8'h72 == r_count_97_io_out ? io_r_114_b : _GEN_19813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19815 = 8'h73 == r_count_97_io_out ? io_r_115_b : _GEN_19814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19816 = 8'h74 == r_count_97_io_out ? io_r_116_b : _GEN_19815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19817 = 8'h75 == r_count_97_io_out ? io_r_117_b : _GEN_19816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19818 = 8'h76 == r_count_97_io_out ? io_r_118_b : _GEN_19817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19819 = 8'h77 == r_count_97_io_out ? io_r_119_b : _GEN_19818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19820 = 8'h78 == r_count_97_io_out ? io_r_120_b : _GEN_19819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19821 = 8'h79 == r_count_97_io_out ? io_r_121_b : _GEN_19820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19822 = 8'h7a == r_count_97_io_out ? io_r_122_b : _GEN_19821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19823 = 8'h7b == r_count_97_io_out ? io_r_123_b : _GEN_19822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19824 = 8'h7c == r_count_97_io_out ? io_r_124_b : _GEN_19823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19825 = 8'h7d == r_count_97_io_out ? io_r_125_b : _GEN_19824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19826 = 8'h7e == r_count_97_io_out ? io_r_126_b : _GEN_19825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19827 = 8'h7f == r_count_97_io_out ? io_r_127_b : _GEN_19826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19828 = 8'h80 == r_count_97_io_out ? io_r_128_b : _GEN_19827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19829 = 8'h81 == r_count_97_io_out ? io_r_129_b : _GEN_19828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19830 = 8'h82 == r_count_97_io_out ? io_r_130_b : _GEN_19829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19831 = 8'h83 == r_count_97_io_out ? io_r_131_b : _GEN_19830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19832 = 8'h84 == r_count_97_io_out ? io_r_132_b : _GEN_19831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19833 = 8'h85 == r_count_97_io_out ? io_r_133_b : _GEN_19832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19834 = 8'h86 == r_count_97_io_out ? io_r_134_b : _GEN_19833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19835 = 8'h87 == r_count_97_io_out ? io_r_135_b : _GEN_19834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19836 = 8'h88 == r_count_97_io_out ? io_r_136_b : _GEN_19835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19837 = 8'h89 == r_count_97_io_out ? io_r_137_b : _GEN_19836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19838 = 8'h8a == r_count_97_io_out ? io_r_138_b : _GEN_19837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19839 = 8'h8b == r_count_97_io_out ? io_r_139_b : _GEN_19838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19840 = 8'h8c == r_count_97_io_out ? io_r_140_b : _GEN_19839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19841 = 8'h8d == r_count_97_io_out ? io_r_141_b : _GEN_19840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19842 = 8'h8e == r_count_97_io_out ? io_r_142_b : _GEN_19841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19843 = 8'h8f == r_count_97_io_out ? io_r_143_b : _GEN_19842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19844 = 8'h90 == r_count_97_io_out ? io_r_144_b : _GEN_19843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19845 = 8'h91 == r_count_97_io_out ? io_r_145_b : _GEN_19844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19846 = 8'h92 == r_count_97_io_out ? io_r_146_b : _GEN_19845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19847 = 8'h93 == r_count_97_io_out ? io_r_147_b : _GEN_19846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19848 = 8'h94 == r_count_97_io_out ? io_r_148_b : _GEN_19847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19849 = 8'h95 == r_count_97_io_out ? io_r_149_b : _GEN_19848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19850 = 8'h96 == r_count_97_io_out ? io_r_150_b : _GEN_19849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19851 = 8'h97 == r_count_97_io_out ? io_r_151_b : _GEN_19850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19852 = 8'h98 == r_count_97_io_out ? io_r_152_b : _GEN_19851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19853 = 8'h99 == r_count_97_io_out ? io_r_153_b : _GEN_19852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19854 = 8'h9a == r_count_97_io_out ? io_r_154_b : _GEN_19853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19855 = 8'h9b == r_count_97_io_out ? io_r_155_b : _GEN_19854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19856 = 8'h9c == r_count_97_io_out ? io_r_156_b : _GEN_19855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19857 = 8'h9d == r_count_97_io_out ? io_r_157_b : _GEN_19856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19858 = 8'h9e == r_count_97_io_out ? io_r_158_b : _GEN_19857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19859 = 8'h9f == r_count_97_io_out ? io_r_159_b : _GEN_19858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19860 = 8'ha0 == r_count_97_io_out ? io_r_160_b : _GEN_19859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19861 = 8'ha1 == r_count_97_io_out ? io_r_161_b : _GEN_19860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19862 = 8'ha2 == r_count_97_io_out ? io_r_162_b : _GEN_19861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19863 = 8'ha3 == r_count_97_io_out ? io_r_163_b : _GEN_19862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19864 = 8'ha4 == r_count_97_io_out ? io_r_164_b : _GEN_19863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19865 = 8'ha5 == r_count_97_io_out ? io_r_165_b : _GEN_19864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19866 = 8'ha6 == r_count_97_io_out ? io_r_166_b : _GEN_19865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19867 = 8'ha7 == r_count_97_io_out ? io_r_167_b : _GEN_19866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19868 = 8'ha8 == r_count_97_io_out ? io_r_168_b : _GEN_19867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19869 = 8'ha9 == r_count_97_io_out ? io_r_169_b : _GEN_19868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19870 = 8'haa == r_count_97_io_out ? io_r_170_b : _GEN_19869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19871 = 8'hab == r_count_97_io_out ? io_r_171_b : _GEN_19870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19872 = 8'hac == r_count_97_io_out ? io_r_172_b : _GEN_19871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19873 = 8'had == r_count_97_io_out ? io_r_173_b : _GEN_19872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19874 = 8'hae == r_count_97_io_out ? io_r_174_b : _GEN_19873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19875 = 8'haf == r_count_97_io_out ? io_r_175_b : _GEN_19874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19876 = 8'hb0 == r_count_97_io_out ? io_r_176_b : _GEN_19875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19877 = 8'hb1 == r_count_97_io_out ? io_r_177_b : _GEN_19876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19878 = 8'hb2 == r_count_97_io_out ? io_r_178_b : _GEN_19877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19879 = 8'hb3 == r_count_97_io_out ? io_r_179_b : _GEN_19878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19880 = 8'hb4 == r_count_97_io_out ? io_r_180_b : _GEN_19879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19881 = 8'hb5 == r_count_97_io_out ? io_r_181_b : _GEN_19880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19882 = 8'hb6 == r_count_97_io_out ? io_r_182_b : _GEN_19881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19883 = 8'hb7 == r_count_97_io_out ? io_r_183_b : _GEN_19882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19884 = 8'hb8 == r_count_97_io_out ? io_r_184_b : _GEN_19883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19885 = 8'hb9 == r_count_97_io_out ? io_r_185_b : _GEN_19884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19886 = 8'hba == r_count_97_io_out ? io_r_186_b : _GEN_19885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19887 = 8'hbb == r_count_97_io_out ? io_r_187_b : _GEN_19886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19888 = 8'hbc == r_count_97_io_out ? io_r_188_b : _GEN_19887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19889 = 8'hbd == r_count_97_io_out ? io_r_189_b : _GEN_19888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19890 = 8'hbe == r_count_97_io_out ? io_r_190_b : _GEN_19889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19891 = 8'hbf == r_count_97_io_out ? io_r_191_b : _GEN_19890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19892 = 8'hc0 == r_count_97_io_out ? io_r_192_b : _GEN_19891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19893 = 8'hc1 == r_count_97_io_out ? io_r_193_b : _GEN_19892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19894 = 8'hc2 == r_count_97_io_out ? io_r_194_b : _GEN_19893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19895 = 8'hc3 == r_count_97_io_out ? io_r_195_b : _GEN_19894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19896 = 8'hc4 == r_count_97_io_out ? io_r_196_b : _GEN_19895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19897 = 8'hc5 == r_count_97_io_out ? io_r_197_b : _GEN_19896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19898 = 8'hc6 == r_count_97_io_out ? io_r_198_b : _GEN_19897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19901 = 8'h1 == r_count_98_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19902 = 8'h2 == r_count_98_io_out ? io_r_2_b : _GEN_19901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19903 = 8'h3 == r_count_98_io_out ? io_r_3_b : _GEN_19902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19904 = 8'h4 == r_count_98_io_out ? io_r_4_b : _GEN_19903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19905 = 8'h5 == r_count_98_io_out ? io_r_5_b : _GEN_19904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19906 = 8'h6 == r_count_98_io_out ? io_r_6_b : _GEN_19905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19907 = 8'h7 == r_count_98_io_out ? io_r_7_b : _GEN_19906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19908 = 8'h8 == r_count_98_io_out ? io_r_8_b : _GEN_19907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19909 = 8'h9 == r_count_98_io_out ? io_r_9_b : _GEN_19908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19910 = 8'ha == r_count_98_io_out ? io_r_10_b : _GEN_19909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19911 = 8'hb == r_count_98_io_out ? io_r_11_b : _GEN_19910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19912 = 8'hc == r_count_98_io_out ? io_r_12_b : _GEN_19911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19913 = 8'hd == r_count_98_io_out ? io_r_13_b : _GEN_19912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19914 = 8'he == r_count_98_io_out ? io_r_14_b : _GEN_19913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19915 = 8'hf == r_count_98_io_out ? io_r_15_b : _GEN_19914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19916 = 8'h10 == r_count_98_io_out ? io_r_16_b : _GEN_19915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19917 = 8'h11 == r_count_98_io_out ? io_r_17_b : _GEN_19916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19918 = 8'h12 == r_count_98_io_out ? io_r_18_b : _GEN_19917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19919 = 8'h13 == r_count_98_io_out ? io_r_19_b : _GEN_19918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19920 = 8'h14 == r_count_98_io_out ? io_r_20_b : _GEN_19919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19921 = 8'h15 == r_count_98_io_out ? io_r_21_b : _GEN_19920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19922 = 8'h16 == r_count_98_io_out ? io_r_22_b : _GEN_19921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19923 = 8'h17 == r_count_98_io_out ? io_r_23_b : _GEN_19922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19924 = 8'h18 == r_count_98_io_out ? io_r_24_b : _GEN_19923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19925 = 8'h19 == r_count_98_io_out ? io_r_25_b : _GEN_19924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19926 = 8'h1a == r_count_98_io_out ? io_r_26_b : _GEN_19925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19927 = 8'h1b == r_count_98_io_out ? io_r_27_b : _GEN_19926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19928 = 8'h1c == r_count_98_io_out ? io_r_28_b : _GEN_19927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19929 = 8'h1d == r_count_98_io_out ? io_r_29_b : _GEN_19928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19930 = 8'h1e == r_count_98_io_out ? io_r_30_b : _GEN_19929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19931 = 8'h1f == r_count_98_io_out ? io_r_31_b : _GEN_19930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19932 = 8'h20 == r_count_98_io_out ? io_r_32_b : _GEN_19931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19933 = 8'h21 == r_count_98_io_out ? io_r_33_b : _GEN_19932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19934 = 8'h22 == r_count_98_io_out ? io_r_34_b : _GEN_19933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19935 = 8'h23 == r_count_98_io_out ? io_r_35_b : _GEN_19934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19936 = 8'h24 == r_count_98_io_out ? io_r_36_b : _GEN_19935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19937 = 8'h25 == r_count_98_io_out ? io_r_37_b : _GEN_19936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19938 = 8'h26 == r_count_98_io_out ? io_r_38_b : _GEN_19937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19939 = 8'h27 == r_count_98_io_out ? io_r_39_b : _GEN_19938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19940 = 8'h28 == r_count_98_io_out ? io_r_40_b : _GEN_19939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19941 = 8'h29 == r_count_98_io_out ? io_r_41_b : _GEN_19940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19942 = 8'h2a == r_count_98_io_out ? io_r_42_b : _GEN_19941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19943 = 8'h2b == r_count_98_io_out ? io_r_43_b : _GEN_19942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19944 = 8'h2c == r_count_98_io_out ? io_r_44_b : _GEN_19943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19945 = 8'h2d == r_count_98_io_out ? io_r_45_b : _GEN_19944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19946 = 8'h2e == r_count_98_io_out ? io_r_46_b : _GEN_19945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19947 = 8'h2f == r_count_98_io_out ? io_r_47_b : _GEN_19946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19948 = 8'h30 == r_count_98_io_out ? io_r_48_b : _GEN_19947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19949 = 8'h31 == r_count_98_io_out ? io_r_49_b : _GEN_19948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19950 = 8'h32 == r_count_98_io_out ? io_r_50_b : _GEN_19949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19951 = 8'h33 == r_count_98_io_out ? io_r_51_b : _GEN_19950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19952 = 8'h34 == r_count_98_io_out ? io_r_52_b : _GEN_19951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19953 = 8'h35 == r_count_98_io_out ? io_r_53_b : _GEN_19952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19954 = 8'h36 == r_count_98_io_out ? io_r_54_b : _GEN_19953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19955 = 8'h37 == r_count_98_io_out ? io_r_55_b : _GEN_19954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19956 = 8'h38 == r_count_98_io_out ? io_r_56_b : _GEN_19955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19957 = 8'h39 == r_count_98_io_out ? io_r_57_b : _GEN_19956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19958 = 8'h3a == r_count_98_io_out ? io_r_58_b : _GEN_19957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19959 = 8'h3b == r_count_98_io_out ? io_r_59_b : _GEN_19958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19960 = 8'h3c == r_count_98_io_out ? io_r_60_b : _GEN_19959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19961 = 8'h3d == r_count_98_io_out ? io_r_61_b : _GEN_19960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19962 = 8'h3e == r_count_98_io_out ? io_r_62_b : _GEN_19961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19963 = 8'h3f == r_count_98_io_out ? io_r_63_b : _GEN_19962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19964 = 8'h40 == r_count_98_io_out ? io_r_64_b : _GEN_19963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19965 = 8'h41 == r_count_98_io_out ? io_r_65_b : _GEN_19964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19966 = 8'h42 == r_count_98_io_out ? io_r_66_b : _GEN_19965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19967 = 8'h43 == r_count_98_io_out ? io_r_67_b : _GEN_19966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19968 = 8'h44 == r_count_98_io_out ? io_r_68_b : _GEN_19967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19969 = 8'h45 == r_count_98_io_out ? io_r_69_b : _GEN_19968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19970 = 8'h46 == r_count_98_io_out ? io_r_70_b : _GEN_19969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19971 = 8'h47 == r_count_98_io_out ? io_r_71_b : _GEN_19970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19972 = 8'h48 == r_count_98_io_out ? io_r_72_b : _GEN_19971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19973 = 8'h49 == r_count_98_io_out ? io_r_73_b : _GEN_19972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19974 = 8'h4a == r_count_98_io_out ? io_r_74_b : _GEN_19973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19975 = 8'h4b == r_count_98_io_out ? io_r_75_b : _GEN_19974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19976 = 8'h4c == r_count_98_io_out ? io_r_76_b : _GEN_19975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19977 = 8'h4d == r_count_98_io_out ? io_r_77_b : _GEN_19976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19978 = 8'h4e == r_count_98_io_out ? io_r_78_b : _GEN_19977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19979 = 8'h4f == r_count_98_io_out ? io_r_79_b : _GEN_19978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19980 = 8'h50 == r_count_98_io_out ? io_r_80_b : _GEN_19979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19981 = 8'h51 == r_count_98_io_out ? io_r_81_b : _GEN_19980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19982 = 8'h52 == r_count_98_io_out ? io_r_82_b : _GEN_19981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19983 = 8'h53 == r_count_98_io_out ? io_r_83_b : _GEN_19982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19984 = 8'h54 == r_count_98_io_out ? io_r_84_b : _GEN_19983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19985 = 8'h55 == r_count_98_io_out ? io_r_85_b : _GEN_19984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19986 = 8'h56 == r_count_98_io_out ? io_r_86_b : _GEN_19985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19987 = 8'h57 == r_count_98_io_out ? io_r_87_b : _GEN_19986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19988 = 8'h58 == r_count_98_io_out ? io_r_88_b : _GEN_19987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19989 = 8'h59 == r_count_98_io_out ? io_r_89_b : _GEN_19988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19990 = 8'h5a == r_count_98_io_out ? io_r_90_b : _GEN_19989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19991 = 8'h5b == r_count_98_io_out ? io_r_91_b : _GEN_19990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19992 = 8'h5c == r_count_98_io_out ? io_r_92_b : _GEN_19991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19993 = 8'h5d == r_count_98_io_out ? io_r_93_b : _GEN_19992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19994 = 8'h5e == r_count_98_io_out ? io_r_94_b : _GEN_19993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19995 = 8'h5f == r_count_98_io_out ? io_r_95_b : _GEN_19994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19996 = 8'h60 == r_count_98_io_out ? io_r_96_b : _GEN_19995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19997 = 8'h61 == r_count_98_io_out ? io_r_97_b : _GEN_19996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19998 = 8'h62 == r_count_98_io_out ? io_r_98_b : _GEN_19997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_19999 = 8'h63 == r_count_98_io_out ? io_r_99_b : _GEN_19998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20000 = 8'h64 == r_count_98_io_out ? io_r_100_b : _GEN_19999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20001 = 8'h65 == r_count_98_io_out ? io_r_101_b : _GEN_20000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20002 = 8'h66 == r_count_98_io_out ? io_r_102_b : _GEN_20001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20003 = 8'h67 == r_count_98_io_out ? io_r_103_b : _GEN_20002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20004 = 8'h68 == r_count_98_io_out ? io_r_104_b : _GEN_20003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20005 = 8'h69 == r_count_98_io_out ? io_r_105_b : _GEN_20004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20006 = 8'h6a == r_count_98_io_out ? io_r_106_b : _GEN_20005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20007 = 8'h6b == r_count_98_io_out ? io_r_107_b : _GEN_20006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20008 = 8'h6c == r_count_98_io_out ? io_r_108_b : _GEN_20007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20009 = 8'h6d == r_count_98_io_out ? io_r_109_b : _GEN_20008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20010 = 8'h6e == r_count_98_io_out ? io_r_110_b : _GEN_20009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20011 = 8'h6f == r_count_98_io_out ? io_r_111_b : _GEN_20010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20012 = 8'h70 == r_count_98_io_out ? io_r_112_b : _GEN_20011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20013 = 8'h71 == r_count_98_io_out ? io_r_113_b : _GEN_20012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20014 = 8'h72 == r_count_98_io_out ? io_r_114_b : _GEN_20013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20015 = 8'h73 == r_count_98_io_out ? io_r_115_b : _GEN_20014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20016 = 8'h74 == r_count_98_io_out ? io_r_116_b : _GEN_20015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20017 = 8'h75 == r_count_98_io_out ? io_r_117_b : _GEN_20016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20018 = 8'h76 == r_count_98_io_out ? io_r_118_b : _GEN_20017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20019 = 8'h77 == r_count_98_io_out ? io_r_119_b : _GEN_20018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20020 = 8'h78 == r_count_98_io_out ? io_r_120_b : _GEN_20019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20021 = 8'h79 == r_count_98_io_out ? io_r_121_b : _GEN_20020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20022 = 8'h7a == r_count_98_io_out ? io_r_122_b : _GEN_20021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20023 = 8'h7b == r_count_98_io_out ? io_r_123_b : _GEN_20022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20024 = 8'h7c == r_count_98_io_out ? io_r_124_b : _GEN_20023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20025 = 8'h7d == r_count_98_io_out ? io_r_125_b : _GEN_20024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20026 = 8'h7e == r_count_98_io_out ? io_r_126_b : _GEN_20025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20027 = 8'h7f == r_count_98_io_out ? io_r_127_b : _GEN_20026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20028 = 8'h80 == r_count_98_io_out ? io_r_128_b : _GEN_20027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20029 = 8'h81 == r_count_98_io_out ? io_r_129_b : _GEN_20028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20030 = 8'h82 == r_count_98_io_out ? io_r_130_b : _GEN_20029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20031 = 8'h83 == r_count_98_io_out ? io_r_131_b : _GEN_20030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20032 = 8'h84 == r_count_98_io_out ? io_r_132_b : _GEN_20031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20033 = 8'h85 == r_count_98_io_out ? io_r_133_b : _GEN_20032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20034 = 8'h86 == r_count_98_io_out ? io_r_134_b : _GEN_20033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20035 = 8'h87 == r_count_98_io_out ? io_r_135_b : _GEN_20034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20036 = 8'h88 == r_count_98_io_out ? io_r_136_b : _GEN_20035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20037 = 8'h89 == r_count_98_io_out ? io_r_137_b : _GEN_20036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20038 = 8'h8a == r_count_98_io_out ? io_r_138_b : _GEN_20037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20039 = 8'h8b == r_count_98_io_out ? io_r_139_b : _GEN_20038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20040 = 8'h8c == r_count_98_io_out ? io_r_140_b : _GEN_20039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20041 = 8'h8d == r_count_98_io_out ? io_r_141_b : _GEN_20040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20042 = 8'h8e == r_count_98_io_out ? io_r_142_b : _GEN_20041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20043 = 8'h8f == r_count_98_io_out ? io_r_143_b : _GEN_20042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20044 = 8'h90 == r_count_98_io_out ? io_r_144_b : _GEN_20043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20045 = 8'h91 == r_count_98_io_out ? io_r_145_b : _GEN_20044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20046 = 8'h92 == r_count_98_io_out ? io_r_146_b : _GEN_20045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20047 = 8'h93 == r_count_98_io_out ? io_r_147_b : _GEN_20046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20048 = 8'h94 == r_count_98_io_out ? io_r_148_b : _GEN_20047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20049 = 8'h95 == r_count_98_io_out ? io_r_149_b : _GEN_20048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20050 = 8'h96 == r_count_98_io_out ? io_r_150_b : _GEN_20049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20051 = 8'h97 == r_count_98_io_out ? io_r_151_b : _GEN_20050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20052 = 8'h98 == r_count_98_io_out ? io_r_152_b : _GEN_20051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20053 = 8'h99 == r_count_98_io_out ? io_r_153_b : _GEN_20052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20054 = 8'h9a == r_count_98_io_out ? io_r_154_b : _GEN_20053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20055 = 8'h9b == r_count_98_io_out ? io_r_155_b : _GEN_20054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20056 = 8'h9c == r_count_98_io_out ? io_r_156_b : _GEN_20055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20057 = 8'h9d == r_count_98_io_out ? io_r_157_b : _GEN_20056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20058 = 8'h9e == r_count_98_io_out ? io_r_158_b : _GEN_20057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20059 = 8'h9f == r_count_98_io_out ? io_r_159_b : _GEN_20058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20060 = 8'ha0 == r_count_98_io_out ? io_r_160_b : _GEN_20059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20061 = 8'ha1 == r_count_98_io_out ? io_r_161_b : _GEN_20060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20062 = 8'ha2 == r_count_98_io_out ? io_r_162_b : _GEN_20061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20063 = 8'ha3 == r_count_98_io_out ? io_r_163_b : _GEN_20062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20064 = 8'ha4 == r_count_98_io_out ? io_r_164_b : _GEN_20063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20065 = 8'ha5 == r_count_98_io_out ? io_r_165_b : _GEN_20064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20066 = 8'ha6 == r_count_98_io_out ? io_r_166_b : _GEN_20065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20067 = 8'ha7 == r_count_98_io_out ? io_r_167_b : _GEN_20066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20068 = 8'ha8 == r_count_98_io_out ? io_r_168_b : _GEN_20067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20069 = 8'ha9 == r_count_98_io_out ? io_r_169_b : _GEN_20068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20070 = 8'haa == r_count_98_io_out ? io_r_170_b : _GEN_20069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20071 = 8'hab == r_count_98_io_out ? io_r_171_b : _GEN_20070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20072 = 8'hac == r_count_98_io_out ? io_r_172_b : _GEN_20071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20073 = 8'had == r_count_98_io_out ? io_r_173_b : _GEN_20072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20074 = 8'hae == r_count_98_io_out ? io_r_174_b : _GEN_20073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20075 = 8'haf == r_count_98_io_out ? io_r_175_b : _GEN_20074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20076 = 8'hb0 == r_count_98_io_out ? io_r_176_b : _GEN_20075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20077 = 8'hb1 == r_count_98_io_out ? io_r_177_b : _GEN_20076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20078 = 8'hb2 == r_count_98_io_out ? io_r_178_b : _GEN_20077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20079 = 8'hb3 == r_count_98_io_out ? io_r_179_b : _GEN_20078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20080 = 8'hb4 == r_count_98_io_out ? io_r_180_b : _GEN_20079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20081 = 8'hb5 == r_count_98_io_out ? io_r_181_b : _GEN_20080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20082 = 8'hb6 == r_count_98_io_out ? io_r_182_b : _GEN_20081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20083 = 8'hb7 == r_count_98_io_out ? io_r_183_b : _GEN_20082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20084 = 8'hb8 == r_count_98_io_out ? io_r_184_b : _GEN_20083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20085 = 8'hb9 == r_count_98_io_out ? io_r_185_b : _GEN_20084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20086 = 8'hba == r_count_98_io_out ? io_r_186_b : _GEN_20085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20087 = 8'hbb == r_count_98_io_out ? io_r_187_b : _GEN_20086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20088 = 8'hbc == r_count_98_io_out ? io_r_188_b : _GEN_20087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20089 = 8'hbd == r_count_98_io_out ? io_r_189_b : _GEN_20088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20090 = 8'hbe == r_count_98_io_out ? io_r_190_b : _GEN_20089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20091 = 8'hbf == r_count_98_io_out ? io_r_191_b : _GEN_20090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20092 = 8'hc0 == r_count_98_io_out ? io_r_192_b : _GEN_20091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20093 = 8'hc1 == r_count_98_io_out ? io_r_193_b : _GEN_20092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20094 = 8'hc2 == r_count_98_io_out ? io_r_194_b : _GEN_20093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20095 = 8'hc3 == r_count_98_io_out ? io_r_195_b : _GEN_20094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20096 = 8'hc4 == r_count_98_io_out ? io_r_196_b : _GEN_20095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20097 = 8'hc5 == r_count_98_io_out ? io_r_197_b : _GEN_20096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20098 = 8'hc6 == r_count_98_io_out ? io_r_198_b : _GEN_20097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20101 = 8'h1 == r_count_99_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20102 = 8'h2 == r_count_99_io_out ? io_r_2_b : _GEN_20101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20103 = 8'h3 == r_count_99_io_out ? io_r_3_b : _GEN_20102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20104 = 8'h4 == r_count_99_io_out ? io_r_4_b : _GEN_20103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20105 = 8'h5 == r_count_99_io_out ? io_r_5_b : _GEN_20104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20106 = 8'h6 == r_count_99_io_out ? io_r_6_b : _GEN_20105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20107 = 8'h7 == r_count_99_io_out ? io_r_7_b : _GEN_20106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20108 = 8'h8 == r_count_99_io_out ? io_r_8_b : _GEN_20107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20109 = 8'h9 == r_count_99_io_out ? io_r_9_b : _GEN_20108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20110 = 8'ha == r_count_99_io_out ? io_r_10_b : _GEN_20109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20111 = 8'hb == r_count_99_io_out ? io_r_11_b : _GEN_20110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20112 = 8'hc == r_count_99_io_out ? io_r_12_b : _GEN_20111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20113 = 8'hd == r_count_99_io_out ? io_r_13_b : _GEN_20112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20114 = 8'he == r_count_99_io_out ? io_r_14_b : _GEN_20113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20115 = 8'hf == r_count_99_io_out ? io_r_15_b : _GEN_20114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20116 = 8'h10 == r_count_99_io_out ? io_r_16_b : _GEN_20115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20117 = 8'h11 == r_count_99_io_out ? io_r_17_b : _GEN_20116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20118 = 8'h12 == r_count_99_io_out ? io_r_18_b : _GEN_20117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20119 = 8'h13 == r_count_99_io_out ? io_r_19_b : _GEN_20118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20120 = 8'h14 == r_count_99_io_out ? io_r_20_b : _GEN_20119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20121 = 8'h15 == r_count_99_io_out ? io_r_21_b : _GEN_20120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20122 = 8'h16 == r_count_99_io_out ? io_r_22_b : _GEN_20121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20123 = 8'h17 == r_count_99_io_out ? io_r_23_b : _GEN_20122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20124 = 8'h18 == r_count_99_io_out ? io_r_24_b : _GEN_20123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20125 = 8'h19 == r_count_99_io_out ? io_r_25_b : _GEN_20124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20126 = 8'h1a == r_count_99_io_out ? io_r_26_b : _GEN_20125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20127 = 8'h1b == r_count_99_io_out ? io_r_27_b : _GEN_20126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20128 = 8'h1c == r_count_99_io_out ? io_r_28_b : _GEN_20127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20129 = 8'h1d == r_count_99_io_out ? io_r_29_b : _GEN_20128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20130 = 8'h1e == r_count_99_io_out ? io_r_30_b : _GEN_20129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20131 = 8'h1f == r_count_99_io_out ? io_r_31_b : _GEN_20130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20132 = 8'h20 == r_count_99_io_out ? io_r_32_b : _GEN_20131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20133 = 8'h21 == r_count_99_io_out ? io_r_33_b : _GEN_20132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20134 = 8'h22 == r_count_99_io_out ? io_r_34_b : _GEN_20133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20135 = 8'h23 == r_count_99_io_out ? io_r_35_b : _GEN_20134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20136 = 8'h24 == r_count_99_io_out ? io_r_36_b : _GEN_20135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20137 = 8'h25 == r_count_99_io_out ? io_r_37_b : _GEN_20136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20138 = 8'h26 == r_count_99_io_out ? io_r_38_b : _GEN_20137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20139 = 8'h27 == r_count_99_io_out ? io_r_39_b : _GEN_20138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20140 = 8'h28 == r_count_99_io_out ? io_r_40_b : _GEN_20139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20141 = 8'h29 == r_count_99_io_out ? io_r_41_b : _GEN_20140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20142 = 8'h2a == r_count_99_io_out ? io_r_42_b : _GEN_20141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20143 = 8'h2b == r_count_99_io_out ? io_r_43_b : _GEN_20142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20144 = 8'h2c == r_count_99_io_out ? io_r_44_b : _GEN_20143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20145 = 8'h2d == r_count_99_io_out ? io_r_45_b : _GEN_20144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20146 = 8'h2e == r_count_99_io_out ? io_r_46_b : _GEN_20145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20147 = 8'h2f == r_count_99_io_out ? io_r_47_b : _GEN_20146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20148 = 8'h30 == r_count_99_io_out ? io_r_48_b : _GEN_20147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20149 = 8'h31 == r_count_99_io_out ? io_r_49_b : _GEN_20148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20150 = 8'h32 == r_count_99_io_out ? io_r_50_b : _GEN_20149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20151 = 8'h33 == r_count_99_io_out ? io_r_51_b : _GEN_20150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20152 = 8'h34 == r_count_99_io_out ? io_r_52_b : _GEN_20151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20153 = 8'h35 == r_count_99_io_out ? io_r_53_b : _GEN_20152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20154 = 8'h36 == r_count_99_io_out ? io_r_54_b : _GEN_20153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20155 = 8'h37 == r_count_99_io_out ? io_r_55_b : _GEN_20154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20156 = 8'h38 == r_count_99_io_out ? io_r_56_b : _GEN_20155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20157 = 8'h39 == r_count_99_io_out ? io_r_57_b : _GEN_20156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20158 = 8'h3a == r_count_99_io_out ? io_r_58_b : _GEN_20157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20159 = 8'h3b == r_count_99_io_out ? io_r_59_b : _GEN_20158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20160 = 8'h3c == r_count_99_io_out ? io_r_60_b : _GEN_20159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20161 = 8'h3d == r_count_99_io_out ? io_r_61_b : _GEN_20160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20162 = 8'h3e == r_count_99_io_out ? io_r_62_b : _GEN_20161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20163 = 8'h3f == r_count_99_io_out ? io_r_63_b : _GEN_20162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20164 = 8'h40 == r_count_99_io_out ? io_r_64_b : _GEN_20163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20165 = 8'h41 == r_count_99_io_out ? io_r_65_b : _GEN_20164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20166 = 8'h42 == r_count_99_io_out ? io_r_66_b : _GEN_20165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20167 = 8'h43 == r_count_99_io_out ? io_r_67_b : _GEN_20166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20168 = 8'h44 == r_count_99_io_out ? io_r_68_b : _GEN_20167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20169 = 8'h45 == r_count_99_io_out ? io_r_69_b : _GEN_20168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20170 = 8'h46 == r_count_99_io_out ? io_r_70_b : _GEN_20169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20171 = 8'h47 == r_count_99_io_out ? io_r_71_b : _GEN_20170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20172 = 8'h48 == r_count_99_io_out ? io_r_72_b : _GEN_20171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20173 = 8'h49 == r_count_99_io_out ? io_r_73_b : _GEN_20172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20174 = 8'h4a == r_count_99_io_out ? io_r_74_b : _GEN_20173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20175 = 8'h4b == r_count_99_io_out ? io_r_75_b : _GEN_20174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20176 = 8'h4c == r_count_99_io_out ? io_r_76_b : _GEN_20175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20177 = 8'h4d == r_count_99_io_out ? io_r_77_b : _GEN_20176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20178 = 8'h4e == r_count_99_io_out ? io_r_78_b : _GEN_20177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20179 = 8'h4f == r_count_99_io_out ? io_r_79_b : _GEN_20178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20180 = 8'h50 == r_count_99_io_out ? io_r_80_b : _GEN_20179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20181 = 8'h51 == r_count_99_io_out ? io_r_81_b : _GEN_20180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20182 = 8'h52 == r_count_99_io_out ? io_r_82_b : _GEN_20181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20183 = 8'h53 == r_count_99_io_out ? io_r_83_b : _GEN_20182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20184 = 8'h54 == r_count_99_io_out ? io_r_84_b : _GEN_20183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20185 = 8'h55 == r_count_99_io_out ? io_r_85_b : _GEN_20184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20186 = 8'h56 == r_count_99_io_out ? io_r_86_b : _GEN_20185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20187 = 8'h57 == r_count_99_io_out ? io_r_87_b : _GEN_20186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20188 = 8'h58 == r_count_99_io_out ? io_r_88_b : _GEN_20187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20189 = 8'h59 == r_count_99_io_out ? io_r_89_b : _GEN_20188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20190 = 8'h5a == r_count_99_io_out ? io_r_90_b : _GEN_20189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20191 = 8'h5b == r_count_99_io_out ? io_r_91_b : _GEN_20190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20192 = 8'h5c == r_count_99_io_out ? io_r_92_b : _GEN_20191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20193 = 8'h5d == r_count_99_io_out ? io_r_93_b : _GEN_20192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20194 = 8'h5e == r_count_99_io_out ? io_r_94_b : _GEN_20193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20195 = 8'h5f == r_count_99_io_out ? io_r_95_b : _GEN_20194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20196 = 8'h60 == r_count_99_io_out ? io_r_96_b : _GEN_20195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20197 = 8'h61 == r_count_99_io_out ? io_r_97_b : _GEN_20196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20198 = 8'h62 == r_count_99_io_out ? io_r_98_b : _GEN_20197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20199 = 8'h63 == r_count_99_io_out ? io_r_99_b : _GEN_20198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20200 = 8'h64 == r_count_99_io_out ? io_r_100_b : _GEN_20199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20201 = 8'h65 == r_count_99_io_out ? io_r_101_b : _GEN_20200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20202 = 8'h66 == r_count_99_io_out ? io_r_102_b : _GEN_20201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20203 = 8'h67 == r_count_99_io_out ? io_r_103_b : _GEN_20202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20204 = 8'h68 == r_count_99_io_out ? io_r_104_b : _GEN_20203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20205 = 8'h69 == r_count_99_io_out ? io_r_105_b : _GEN_20204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20206 = 8'h6a == r_count_99_io_out ? io_r_106_b : _GEN_20205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20207 = 8'h6b == r_count_99_io_out ? io_r_107_b : _GEN_20206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20208 = 8'h6c == r_count_99_io_out ? io_r_108_b : _GEN_20207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20209 = 8'h6d == r_count_99_io_out ? io_r_109_b : _GEN_20208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20210 = 8'h6e == r_count_99_io_out ? io_r_110_b : _GEN_20209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20211 = 8'h6f == r_count_99_io_out ? io_r_111_b : _GEN_20210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20212 = 8'h70 == r_count_99_io_out ? io_r_112_b : _GEN_20211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20213 = 8'h71 == r_count_99_io_out ? io_r_113_b : _GEN_20212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20214 = 8'h72 == r_count_99_io_out ? io_r_114_b : _GEN_20213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20215 = 8'h73 == r_count_99_io_out ? io_r_115_b : _GEN_20214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20216 = 8'h74 == r_count_99_io_out ? io_r_116_b : _GEN_20215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20217 = 8'h75 == r_count_99_io_out ? io_r_117_b : _GEN_20216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20218 = 8'h76 == r_count_99_io_out ? io_r_118_b : _GEN_20217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20219 = 8'h77 == r_count_99_io_out ? io_r_119_b : _GEN_20218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20220 = 8'h78 == r_count_99_io_out ? io_r_120_b : _GEN_20219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20221 = 8'h79 == r_count_99_io_out ? io_r_121_b : _GEN_20220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20222 = 8'h7a == r_count_99_io_out ? io_r_122_b : _GEN_20221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20223 = 8'h7b == r_count_99_io_out ? io_r_123_b : _GEN_20222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20224 = 8'h7c == r_count_99_io_out ? io_r_124_b : _GEN_20223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20225 = 8'h7d == r_count_99_io_out ? io_r_125_b : _GEN_20224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20226 = 8'h7e == r_count_99_io_out ? io_r_126_b : _GEN_20225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20227 = 8'h7f == r_count_99_io_out ? io_r_127_b : _GEN_20226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20228 = 8'h80 == r_count_99_io_out ? io_r_128_b : _GEN_20227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20229 = 8'h81 == r_count_99_io_out ? io_r_129_b : _GEN_20228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20230 = 8'h82 == r_count_99_io_out ? io_r_130_b : _GEN_20229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20231 = 8'h83 == r_count_99_io_out ? io_r_131_b : _GEN_20230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20232 = 8'h84 == r_count_99_io_out ? io_r_132_b : _GEN_20231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20233 = 8'h85 == r_count_99_io_out ? io_r_133_b : _GEN_20232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20234 = 8'h86 == r_count_99_io_out ? io_r_134_b : _GEN_20233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20235 = 8'h87 == r_count_99_io_out ? io_r_135_b : _GEN_20234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20236 = 8'h88 == r_count_99_io_out ? io_r_136_b : _GEN_20235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20237 = 8'h89 == r_count_99_io_out ? io_r_137_b : _GEN_20236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20238 = 8'h8a == r_count_99_io_out ? io_r_138_b : _GEN_20237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20239 = 8'h8b == r_count_99_io_out ? io_r_139_b : _GEN_20238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20240 = 8'h8c == r_count_99_io_out ? io_r_140_b : _GEN_20239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20241 = 8'h8d == r_count_99_io_out ? io_r_141_b : _GEN_20240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20242 = 8'h8e == r_count_99_io_out ? io_r_142_b : _GEN_20241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20243 = 8'h8f == r_count_99_io_out ? io_r_143_b : _GEN_20242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20244 = 8'h90 == r_count_99_io_out ? io_r_144_b : _GEN_20243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20245 = 8'h91 == r_count_99_io_out ? io_r_145_b : _GEN_20244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20246 = 8'h92 == r_count_99_io_out ? io_r_146_b : _GEN_20245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20247 = 8'h93 == r_count_99_io_out ? io_r_147_b : _GEN_20246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20248 = 8'h94 == r_count_99_io_out ? io_r_148_b : _GEN_20247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20249 = 8'h95 == r_count_99_io_out ? io_r_149_b : _GEN_20248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20250 = 8'h96 == r_count_99_io_out ? io_r_150_b : _GEN_20249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20251 = 8'h97 == r_count_99_io_out ? io_r_151_b : _GEN_20250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20252 = 8'h98 == r_count_99_io_out ? io_r_152_b : _GEN_20251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20253 = 8'h99 == r_count_99_io_out ? io_r_153_b : _GEN_20252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20254 = 8'h9a == r_count_99_io_out ? io_r_154_b : _GEN_20253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20255 = 8'h9b == r_count_99_io_out ? io_r_155_b : _GEN_20254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20256 = 8'h9c == r_count_99_io_out ? io_r_156_b : _GEN_20255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20257 = 8'h9d == r_count_99_io_out ? io_r_157_b : _GEN_20256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20258 = 8'h9e == r_count_99_io_out ? io_r_158_b : _GEN_20257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20259 = 8'h9f == r_count_99_io_out ? io_r_159_b : _GEN_20258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20260 = 8'ha0 == r_count_99_io_out ? io_r_160_b : _GEN_20259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20261 = 8'ha1 == r_count_99_io_out ? io_r_161_b : _GEN_20260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20262 = 8'ha2 == r_count_99_io_out ? io_r_162_b : _GEN_20261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20263 = 8'ha3 == r_count_99_io_out ? io_r_163_b : _GEN_20262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20264 = 8'ha4 == r_count_99_io_out ? io_r_164_b : _GEN_20263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20265 = 8'ha5 == r_count_99_io_out ? io_r_165_b : _GEN_20264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20266 = 8'ha6 == r_count_99_io_out ? io_r_166_b : _GEN_20265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20267 = 8'ha7 == r_count_99_io_out ? io_r_167_b : _GEN_20266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20268 = 8'ha8 == r_count_99_io_out ? io_r_168_b : _GEN_20267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20269 = 8'ha9 == r_count_99_io_out ? io_r_169_b : _GEN_20268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20270 = 8'haa == r_count_99_io_out ? io_r_170_b : _GEN_20269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20271 = 8'hab == r_count_99_io_out ? io_r_171_b : _GEN_20270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20272 = 8'hac == r_count_99_io_out ? io_r_172_b : _GEN_20271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20273 = 8'had == r_count_99_io_out ? io_r_173_b : _GEN_20272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20274 = 8'hae == r_count_99_io_out ? io_r_174_b : _GEN_20273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20275 = 8'haf == r_count_99_io_out ? io_r_175_b : _GEN_20274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20276 = 8'hb0 == r_count_99_io_out ? io_r_176_b : _GEN_20275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20277 = 8'hb1 == r_count_99_io_out ? io_r_177_b : _GEN_20276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20278 = 8'hb2 == r_count_99_io_out ? io_r_178_b : _GEN_20277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20279 = 8'hb3 == r_count_99_io_out ? io_r_179_b : _GEN_20278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20280 = 8'hb4 == r_count_99_io_out ? io_r_180_b : _GEN_20279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20281 = 8'hb5 == r_count_99_io_out ? io_r_181_b : _GEN_20280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20282 = 8'hb6 == r_count_99_io_out ? io_r_182_b : _GEN_20281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20283 = 8'hb7 == r_count_99_io_out ? io_r_183_b : _GEN_20282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20284 = 8'hb8 == r_count_99_io_out ? io_r_184_b : _GEN_20283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20285 = 8'hb9 == r_count_99_io_out ? io_r_185_b : _GEN_20284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20286 = 8'hba == r_count_99_io_out ? io_r_186_b : _GEN_20285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20287 = 8'hbb == r_count_99_io_out ? io_r_187_b : _GEN_20286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20288 = 8'hbc == r_count_99_io_out ? io_r_188_b : _GEN_20287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20289 = 8'hbd == r_count_99_io_out ? io_r_189_b : _GEN_20288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20290 = 8'hbe == r_count_99_io_out ? io_r_190_b : _GEN_20289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20291 = 8'hbf == r_count_99_io_out ? io_r_191_b : _GEN_20290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20292 = 8'hc0 == r_count_99_io_out ? io_r_192_b : _GEN_20291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20293 = 8'hc1 == r_count_99_io_out ? io_r_193_b : _GEN_20292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20294 = 8'hc2 == r_count_99_io_out ? io_r_194_b : _GEN_20293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20295 = 8'hc3 == r_count_99_io_out ? io_r_195_b : _GEN_20294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20296 = 8'hc4 == r_count_99_io_out ? io_r_196_b : _GEN_20295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20297 = 8'hc5 == r_count_99_io_out ? io_r_197_b : _GEN_20296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_20298 = 8'hc6 == r_count_99_io_out ? io_r_198_b : _GEN_20297; // @[SWChisel.scala 221:{19,19}]
  SWCell array_0 ( // @[SWChisel.scala 170:39]
    .io_q(array_0_io_q),
    .io_r(array_0_io_r),
    .io_e_i(array_0_io_e_i),
    .io_f_i(array_0_io_f_i),
    .io_ve_i(array_0_io_ve_i),
    .io_vf_i(array_0_io_vf_i),
    .io_vv_i(array_0_io_vv_i),
    .io_e_o(array_0_io_e_o),
    .io_f_o(array_0_io_f_o),
    .io_v_o(array_0_io_v_o)
  );
  SWCell array_1 ( // @[SWChisel.scala 170:39]
    .io_q(array_1_io_q),
    .io_r(array_1_io_r),
    .io_e_i(array_1_io_e_i),
    .io_f_i(array_1_io_f_i),
    .io_ve_i(array_1_io_ve_i),
    .io_vf_i(array_1_io_vf_i),
    .io_vv_i(array_1_io_vv_i),
    .io_e_o(array_1_io_e_o),
    .io_f_o(array_1_io_f_o),
    .io_v_o(array_1_io_v_o)
  );
  SWCell array_2 ( // @[SWChisel.scala 170:39]
    .io_q(array_2_io_q),
    .io_r(array_2_io_r),
    .io_e_i(array_2_io_e_i),
    .io_f_i(array_2_io_f_i),
    .io_ve_i(array_2_io_ve_i),
    .io_vf_i(array_2_io_vf_i),
    .io_vv_i(array_2_io_vv_i),
    .io_e_o(array_2_io_e_o),
    .io_f_o(array_2_io_f_o),
    .io_v_o(array_2_io_v_o)
  );
  SWCell array_3 ( // @[SWChisel.scala 170:39]
    .io_q(array_3_io_q),
    .io_r(array_3_io_r),
    .io_e_i(array_3_io_e_i),
    .io_f_i(array_3_io_f_i),
    .io_ve_i(array_3_io_ve_i),
    .io_vf_i(array_3_io_vf_i),
    .io_vv_i(array_3_io_vv_i),
    .io_e_o(array_3_io_e_o),
    .io_f_o(array_3_io_f_o),
    .io_v_o(array_3_io_v_o)
  );
  SWCell array_4 ( // @[SWChisel.scala 170:39]
    .io_q(array_4_io_q),
    .io_r(array_4_io_r),
    .io_e_i(array_4_io_e_i),
    .io_f_i(array_4_io_f_i),
    .io_ve_i(array_4_io_ve_i),
    .io_vf_i(array_4_io_vf_i),
    .io_vv_i(array_4_io_vv_i),
    .io_e_o(array_4_io_e_o),
    .io_f_o(array_4_io_f_o),
    .io_v_o(array_4_io_v_o)
  );
  SWCell array_5 ( // @[SWChisel.scala 170:39]
    .io_q(array_5_io_q),
    .io_r(array_5_io_r),
    .io_e_i(array_5_io_e_i),
    .io_f_i(array_5_io_f_i),
    .io_ve_i(array_5_io_ve_i),
    .io_vf_i(array_5_io_vf_i),
    .io_vv_i(array_5_io_vv_i),
    .io_e_o(array_5_io_e_o),
    .io_f_o(array_5_io_f_o),
    .io_v_o(array_5_io_v_o)
  );
  SWCell array_6 ( // @[SWChisel.scala 170:39]
    .io_q(array_6_io_q),
    .io_r(array_6_io_r),
    .io_e_i(array_6_io_e_i),
    .io_f_i(array_6_io_f_i),
    .io_ve_i(array_6_io_ve_i),
    .io_vf_i(array_6_io_vf_i),
    .io_vv_i(array_6_io_vv_i),
    .io_e_o(array_6_io_e_o),
    .io_f_o(array_6_io_f_o),
    .io_v_o(array_6_io_v_o)
  );
  SWCell array_7 ( // @[SWChisel.scala 170:39]
    .io_q(array_7_io_q),
    .io_r(array_7_io_r),
    .io_e_i(array_7_io_e_i),
    .io_f_i(array_7_io_f_i),
    .io_ve_i(array_7_io_ve_i),
    .io_vf_i(array_7_io_vf_i),
    .io_vv_i(array_7_io_vv_i),
    .io_e_o(array_7_io_e_o),
    .io_f_o(array_7_io_f_o),
    .io_v_o(array_7_io_v_o)
  );
  SWCell array_8 ( // @[SWChisel.scala 170:39]
    .io_q(array_8_io_q),
    .io_r(array_8_io_r),
    .io_e_i(array_8_io_e_i),
    .io_f_i(array_8_io_f_i),
    .io_ve_i(array_8_io_ve_i),
    .io_vf_i(array_8_io_vf_i),
    .io_vv_i(array_8_io_vv_i),
    .io_e_o(array_8_io_e_o),
    .io_f_o(array_8_io_f_o),
    .io_v_o(array_8_io_v_o)
  );
  SWCell array_9 ( // @[SWChisel.scala 170:39]
    .io_q(array_9_io_q),
    .io_r(array_9_io_r),
    .io_e_i(array_9_io_e_i),
    .io_f_i(array_9_io_f_i),
    .io_ve_i(array_9_io_ve_i),
    .io_vf_i(array_9_io_vf_i),
    .io_vv_i(array_9_io_vv_i),
    .io_e_o(array_9_io_e_o),
    .io_f_o(array_9_io_f_o),
    .io_v_o(array_9_io_v_o)
  );
  SWCell array_10 ( // @[SWChisel.scala 170:39]
    .io_q(array_10_io_q),
    .io_r(array_10_io_r),
    .io_e_i(array_10_io_e_i),
    .io_f_i(array_10_io_f_i),
    .io_ve_i(array_10_io_ve_i),
    .io_vf_i(array_10_io_vf_i),
    .io_vv_i(array_10_io_vv_i),
    .io_e_o(array_10_io_e_o),
    .io_f_o(array_10_io_f_o),
    .io_v_o(array_10_io_v_o)
  );
  SWCell array_11 ( // @[SWChisel.scala 170:39]
    .io_q(array_11_io_q),
    .io_r(array_11_io_r),
    .io_e_i(array_11_io_e_i),
    .io_f_i(array_11_io_f_i),
    .io_ve_i(array_11_io_ve_i),
    .io_vf_i(array_11_io_vf_i),
    .io_vv_i(array_11_io_vv_i),
    .io_e_o(array_11_io_e_o),
    .io_f_o(array_11_io_f_o),
    .io_v_o(array_11_io_v_o)
  );
  SWCell array_12 ( // @[SWChisel.scala 170:39]
    .io_q(array_12_io_q),
    .io_r(array_12_io_r),
    .io_e_i(array_12_io_e_i),
    .io_f_i(array_12_io_f_i),
    .io_ve_i(array_12_io_ve_i),
    .io_vf_i(array_12_io_vf_i),
    .io_vv_i(array_12_io_vv_i),
    .io_e_o(array_12_io_e_o),
    .io_f_o(array_12_io_f_o),
    .io_v_o(array_12_io_v_o)
  );
  SWCell array_13 ( // @[SWChisel.scala 170:39]
    .io_q(array_13_io_q),
    .io_r(array_13_io_r),
    .io_e_i(array_13_io_e_i),
    .io_f_i(array_13_io_f_i),
    .io_ve_i(array_13_io_ve_i),
    .io_vf_i(array_13_io_vf_i),
    .io_vv_i(array_13_io_vv_i),
    .io_e_o(array_13_io_e_o),
    .io_f_o(array_13_io_f_o),
    .io_v_o(array_13_io_v_o)
  );
  SWCell array_14 ( // @[SWChisel.scala 170:39]
    .io_q(array_14_io_q),
    .io_r(array_14_io_r),
    .io_e_i(array_14_io_e_i),
    .io_f_i(array_14_io_f_i),
    .io_ve_i(array_14_io_ve_i),
    .io_vf_i(array_14_io_vf_i),
    .io_vv_i(array_14_io_vv_i),
    .io_e_o(array_14_io_e_o),
    .io_f_o(array_14_io_f_o),
    .io_v_o(array_14_io_v_o)
  );
  SWCell array_15 ( // @[SWChisel.scala 170:39]
    .io_q(array_15_io_q),
    .io_r(array_15_io_r),
    .io_e_i(array_15_io_e_i),
    .io_f_i(array_15_io_f_i),
    .io_ve_i(array_15_io_ve_i),
    .io_vf_i(array_15_io_vf_i),
    .io_vv_i(array_15_io_vv_i),
    .io_e_o(array_15_io_e_o),
    .io_f_o(array_15_io_f_o),
    .io_v_o(array_15_io_v_o)
  );
  SWCell array_16 ( // @[SWChisel.scala 170:39]
    .io_q(array_16_io_q),
    .io_r(array_16_io_r),
    .io_e_i(array_16_io_e_i),
    .io_f_i(array_16_io_f_i),
    .io_ve_i(array_16_io_ve_i),
    .io_vf_i(array_16_io_vf_i),
    .io_vv_i(array_16_io_vv_i),
    .io_e_o(array_16_io_e_o),
    .io_f_o(array_16_io_f_o),
    .io_v_o(array_16_io_v_o)
  );
  SWCell array_17 ( // @[SWChisel.scala 170:39]
    .io_q(array_17_io_q),
    .io_r(array_17_io_r),
    .io_e_i(array_17_io_e_i),
    .io_f_i(array_17_io_f_i),
    .io_ve_i(array_17_io_ve_i),
    .io_vf_i(array_17_io_vf_i),
    .io_vv_i(array_17_io_vv_i),
    .io_e_o(array_17_io_e_o),
    .io_f_o(array_17_io_f_o),
    .io_v_o(array_17_io_v_o)
  );
  SWCell array_18 ( // @[SWChisel.scala 170:39]
    .io_q(array_18_io_q),
    .io_r(array_18_io_r),
    .io_e_i(array_18_io_e_i),
    .io_f_i(array_18_io_f_i),
    .io_ve_i(array_18_io_ve_i),
    .io_vf_i(array_18_io_vf_i),
    .io_vv_i(array_18_io_vv_i),
    .io_e_o(array_18_io_e_o),
    .io_f_o(array_18_io_f_o),
    .io_v_o(array_18_io_v_o)
  );
  SWCell array_19 ( // @[SWChisel.scala 170:39]
    .io_q(array_19_io_q),
    .io_r(array_19_io_r),
    .io_e_i(array_19_io_e_i),
    .io_f_i(array_19_io_f_i),
    .io_ve_i(array_19_io_ve_i),
    .io_vf_i(array_19_io_vf_i),
    .io_vv_i(array_19_io_vv_i),
    .io_e_o(array_19_io_e_o),
    .io_f_o(array_19_io_f_o),
    .io_v_o(array_19_io_v_o)
  );
  SWCell array_20 ( // @[SWChisel.scala 170:39]
    .io_q(array_20_io_q),
    .io_r(array_20_io_r),
    .io_e_i(array_20_io_e_i),
    .io_f_i(array_20_io_f_i),
    .io_ve_i(array_20_io_ve_i),
    .io_vf_i(array_20_io_vf_i),
    .io_vv_i(array_20_io_vv_i),
    .io_e_o(array_20_io_e_o),
    .io_f_o(array_20_io_f_o),
    .io_v_o(array_20_io_v_o)
  );
  SWCell array_21 ( // @[SWChisel.scala 170:39]
    .io_q(array_21_io_q),
    .io_r(array_21_io_r),
    .io_e_i(array_21_io_e_i),
    .io_f_i(array_21_io_f_i),
    .io_ve_i(array_21_io_ve_i),
    .io_vf_i(array_21_io_vf_i),
    .io_vv_i(array_21_io_vv_i),
    .io_e_o(array_21_io_e_o),
    .io_f_o(array_21_io_f_o),
    .io_v_o(array_21_io_v_o)
  );
  SWCell array_22 ( // @[SWChisel.scala 170:39]
    .io_q(array_22_io_q),
    .io_r(array_22_io_r),
    .io_e_i(array_22_io_e_i),
    .io_f_i(array_22_io_f_i),
    .io_ve_i(array_22_io_ve_i),
    .io_vf_i(array_22_io_vf_i),
    .io_vv_i(array_22_io_vv_i),
    .io_e_o(array_22_io_e_o),
    .io_f_o(array_22_io_f_o),
    .io_v_o(array_22_io_v_o)
  );
  SWCell array_23 ( // @[SWChisel.scala 170:39]
    .io_q(array_23_io_q),
    .io_r(array_23_io_r),
    .io_e_i(array_23_io_e_i),
    .io_f_i(array_23_io_f_i),
    .io_ve_i(array_23_io_ve_i),
    .io_vf_i(array_23_io_vf_i),
    .io_vv_i(array_23_io_vv_i),
    .io_e_o(array_23_io_e_o),
    .io_f_o(array_23_io_f_o),
    .io_v_o(array_23_io_v_o)
  );
  SWCell array_24 ( // @[SWChisel.scala 170:39]
    .io_q(array_24_io_q),
    .io_r(array_24_io_r),
    .io_e_i(array_24_io_e_i),
    .io_f_i(array_24_io_f_i),
    .io_ve_i(array_24_io_ve_i),
    .io_vf_i(array_24_io_vf_i),
    .io_vv_i(array_24_io_vv_i),
    .io_e_o(array_24_io_e_o),
    .io_f_o(array_24_io_f_o),
    .io_v_o(array_24_io_v_o)
  );
  SWCell array_25 ( // @[SWChisel.scala 170:39]
    .io_q(array_25_io_q),
    .io_r(array_25_io_r),
    .io_e_i(array_25_io_e_i),
    .io_f_i(array_25_io_f_i),
    .io_ve_i(array_25_io_ve_i),
    .io_vf_i(array_25_io_vf_i),
    .io_vv_i(array_25_io_vv_i),
    .io_e_o(array_25_io_e_o),
    .io_f_o(array_25_io_f_o),
    .io_v_o(array_25_io_v_o)
  );
  SWCell array_26 ( // @[SWChisel.scala 170:39]
    .io_q(array_26_io_q),
    .io_r(array_26_io_r),
    .io_e_i(array_26_io_e_i),
    .io_f_i(array_26_io_f_i),
    .io_ve_i(array_26_io_ve_i),
    .io_vf_i(array_26_io_vf_i),
    .io_vv_i(array_26_io_vv_i),
    .io_e_o(array_26_io_e_o),
    .io_f_o(array_26_io_f_o),
    .io_v_o(array_26_io_v_o)
  );
  SWCell array_27 ( // @[SWChisel.scala 170:39]
    .io_q(array_27_io_q),
    .io_r(array_27_io_r),
    .io_e_i(array_27_io_e_i),
    .io_f_i(array_27_io_f_i),
    .io_ve_i(array_27_io_ve_i),
    .io_vf_i(array_27_io_vf_i),
    .io_vv_i(array_27_io_vv_i),
    .io_e_o(array_27_io_e_o),
    .io_f_o(array_27_io_f_o),
    .io_v_o(array_27_io_v_o)
  );
  SWCell array_28 ( // @[SWChisel.scala 170:39]
    .io_q(array_28_io_q),
    .io_r(array_28_io_r),
    .io_e_i(array_28_io_e_i),
    .io_f_i(array_28_io_f_i),
    .io_ve_i(array_28_io_ve_i),
    .io_vf_i(array_28_io_vf_i),
    .io_vv_i(array_28_io_vv_i),
    .io_e_o(array_28_io_e_o),
    .io_f_o(array_28_io_f_o),
    .io_v_o(array_28_io_v_o)
  );
  SWCell array_29 ( // @[SWChisel.scala 170:39]
    .io_q(array_29_io_q),
    .io_r(array_29_io_r),
    .io_e_i(array_29_io_e_i),
    .io_f_i(array_29_io_f_i),
    .io_ve_i(array_29_io_ve_i),
    .io_vf_i(array_29_io_vf_i),
    .io_vv_i(array_29_io_vv_i),
    .io_e_o(array_29_io_e_o),
    .io_f_o(array_29_io_f_o),
    .io_v_o(array_29_io_v_o)
  );
  SWCell array_30 ( // @[SWChisel.scala 170:39]
    .io_q(array_30_io_q),
    .io_r(array_30_io_r),
    .io_e_i(array_30_io_e_i),
    .io_f_i(array_30_io_f_i),
    .io_ve_i(array_30_io_ve_i),
    .io_vf_i(array_30_io_vf_i),
    .io_vv_i(array_30_io_vv_i),
    .io_e_o(array_30_io_e_o),
    .io_f_o(array_30_io_f_o),
    .io_v_o(array_30_io_v_o)
  );
  SWCell array_31 ( // @[SWChisel.scala 170:39]
    .io_q(array_31_io_q),
    .io_r(array_31_io_r),
    .io_e_i(array_31_io_e_i),
    .io_f_i(array_31_io_f_i),
    .io_ve_i(array_31_io_ve_i),
    .io_vf_i(array_31_io_vf_i),
    .io_vv_i(array_31_io_vv_i),
    .io_e_o(array_31_io_e_o),
    .io_f_o(array_31_io_f_o),
    .io_v_o(array_31_io_v_o)
  );
  SWCell array_32 ( // @[SWChisel.scala 170:39]
    .io_q(array_32_io_q),
    .io_r(array_32_io_r),
    .io_e_i(array_32_io_e_i),
    .io_f_i(array_32_io_f_i),
    .io_ve_i(array_32_io_ve_i),
    .io_vf_i(array_32_io_vf_i),
    .io_vv_i(array_32_io_vv_i),
    .io_e_o(array_32_io_e_o),
    .io_f_o(array_32_io_f_o),
    .io_v_o(array_32_io_v_o)
  );
  SWCell array_33 ( // @[SWChisel.scala 170:39]
    .io_q(array_33_io_q),
    .io_r(array_33_io_r),
    .io_e_i(array_33_io_e_i),
    .io_f_i(array_33_io_f_i),
    .io_ve_i(array_33_io_ve_i),
    .io_vf_i(array_33_io_vf_i),
    .io_vv_i(array_33_io_vv_i),
    .io_e_o(array_33_io_e_o),
    .io_f_o(array_33_io_f_o),
    .io_v_o(array_33_io_v_o)
  );
  SWCell array_34 ( // @[SWChisel.scala 170:39]
    .io_q(array_34_io_q),
    .io_r(array_34_io_r),
    .io_e_i(array_34_io_e_i),
    .io_f_i(array_34_io_f_i),
    .io_ve_i(array_34_io_ve_i),
    .io_vf_i(array_34_io_vf_i),
    .io_vv_i(array_34_io_vv_i),
    .io_e_o(array_34_io_e_o),
    .io_f_o(array_34_io_f_o),
    .io_v_o(array_34_io_v_o)
  );
  SWCell array_35 ( // @[SWChisel.scala 170:39]
    .io_q(array_35_io_q),
    .io_r(array_35_io_r),
    .io_e_i(array_35_io_e_i),
    .io_f_i(array_35_io_f_i),
    .io_ve_i(array_35_io_ve_i),
    .io_vf_i(array_35_io_vf_i),
    .io_vv_i(array_35_io_vv_i),
    .io_e_o(array_35_io_e_o),
    .io_f_o(array_35_io_f_o),
    .io_v_o(array_35_io_v_o)
  );
  SWCell array_36 ( // @[SWChisel.scala 170:39]
    .io_q(array_36_io_q),
    .io_r(array_36_io_r),
    .io_e_i(array_36_io_e_i),
    .io_f_i(array_36_io_f_i),
    .io_ve_i(array_36_io_ve_i),
    .io_vf_i(array_36_io_vf_i),
    .io_vv_i(array_36_io_vv_i),
    .io_e_o(array_36_io_e_o),
    .io_f_o(array_36_io_f_o),
    .io_v_o(array_36_io_v_o)
  );
  SWCell array_37 ( // @[SWChisel.scala 170:39]
    .io_q(array_37_io_q),
    .io_r(array_37_io_r),
    .io_e_i(array_37_io_e_i),
    .io_f_i(array_37_io_f_i),
    .io_ve_i(array_37_io_ve_i),
    .io_vf_i(array_37_io_vf_i),
    .io_vv_i(array_37_io_vv_i),
    .io_e_o(array_37_io_e_o),
    .io_f_o(array_37_io_f_o),
    .io_v_o(array_37_io_v_o)
  );
  SWCell array_38 ( // @[SWChisel.scala 170:39]
    .io_q(array_38_io_q),
    .io_r(array_38_io_r),
    .io_e_i(array_38_io_e_i),
    .io_f_i(array_38_io_f_i),
    .io_ve_i(array_38_io_ve_i),
    .io_vf_i(array_38_io_vf_i),
    .io_vv_i(array_38_io_vv_i),
    .io_e_o(array_38_io_e_o),
    .io_f_o(array_38_io_f_o),
    .io_v_o(array_38_io_v_o)
  );
  SWCell array_39 ( // @[SWChisel.scala 170:39]
    .io_q(array_39_io_q),
    .io_r(array_39_io_r),
    .io_e_i(array_39_io_e_i),
    .io_f_i(array_39_io_f_i),
    .io_ve_i(array_39_io_ve_i),
    .io_vf_i(array_39_io_vf_i),
    .io_vv_i(array_39_io_vv_i),
    .io_e_o(array_39_io_e_o),
    .io_f_o(array_39_io_f_o),
    .io_v_o(array_39_io_v_o)
  );
  SWCell array_40 ( // @[SWChisel.scala 170:39]
    .io_q(array_40_io_q),
    .io_r(array_40_io_r),
    .io_e_i(array_40_io_e_i),
    .io_f_i(array_40_io_f_i),
    .io_ve_i(array_40_io_ve_i),
    .io_vf_i(array_40_io_vf_i),
    .io_vv_i(array_40_io_vv_i),
    .io_e_o(array_40_io_e_o),
    .io_f_o(array_40_io_f_o),
    .io_v_o(array_40_io_v_o)
  );
  SWCell array_41 ( // @[SWChisel.scala 170:39]
    .io_q(array_41_io_q),
    .io_r(array_41_io_r),
    .io_e_i(array_41_io_e_i),
    .io_f_i(array_41_io_f_i),
    .io_ve_i(array_41_io_ve_i),
    .io_vf_i(array_41_io_vf_i),
    .io_vv_i(array_41_io_vv_i),
    .io_e_o(array_41_io_e_o),
    .io_f_o(array_41_io_f_o),
    .io_v_o(array_41_io_v_o)
  );
  SWCell array_42 ( // @[SWChisel.scala 170:39]
    .io_q(array_42_io_q),
    .io_r(array_42_io_r),
    .io_e_i(array_42_io_e_i),
    .io_f_i(array_42_io_f_i),
    .io_ve_i(array_42_io_ve_i),
    .io_vf_i(array_42_io_vf_i),
    .io_vv_i(array_42_io_vv_i),
    .io_e_o(array_42_io_e_o),
    .io_f_o(array_42_io_f_o),
    .io_v_o(array_42_io_v_o)
  );
  SWCell array_43 ( // @[SWChisel.scala 170:39]
    .io_q(array_43_io_q),
    .io_r(array_43_io_r),
    .io_e_i(array_43_io_e_i),
    .io_f_i(array_43_io_f_i),
    .io_ve_i(array_43_io_ve_i),
    .io_vf_i(array_43_io_vf_i),
    .io_vv_i(array_43_io_vv_i),
    .io_e_o(array_43_io_e_o),
    .io_f_o(array_43_io_f_o),
    .io_v_o(array_43_io_v_o)
  );
  SWCell array_44 ( // @[SWChisel.scala 170:39]
    .io_q(array_44_io_q),
    .io_r(array_44_io_r),
    .io_e_i(array_44_io_e_i),
    .io_f_i(array_44_io_f_i),
    .io_ve_i(array_44_io_ve_i),
    .io_vf_i(array_44_io_vf_i),
    .io_vv_i(array_44_io_vv_i),
    .io_e_o(array_44_io_e_o),
    .io_f_o(array_44_io_f_o),
    .io_v_o(array_44_io_v_o)
  );
  SWCell array_45 ( // @[SWChisel.scala 170:39]
    .io_q(array_45_io_q),
    .io_r(array_45_io_r),
    .io_e_i(array_45_io_e_i),
    .io_f_i(array_45_io_f_i),
    .io_ve_i(array_45_io_ve_i),
    .io_vf_i(array_45_io_vf_i),
    .io_vv_i(array_45_io_vv_i),
    .io_e_o(array_45_io_e_o),
    .io_f_o(array_45_io_f_o),
    .io_v_o(array_45_io_v_o)
  );
  SWCell array_46 ( // @[SWChisel.scala 170:39]
    .io_q(array_46_io_q),
    .io_r(array_46_io_r),
    .io_e_i(array_46_io_e_i),
    .io_f_i(array_46_io_f_i),
    .io_ve_i(array_46_io_ve_i),
    .io_vf_i(array_46_io_vf_i),
    .io_vv_i(array_46_io_vv_i),
    .io_e_o(array_46_io_e_o),
    .io_f_o(array_46_io_f_o),
    .io_v_o(array_46_io_v_o)
  );
  SWCell array_47 ( // @[SWChisel.scala 170:39]
    .io_q(array_47_io_q),
    .io_r(array_47_io_r),
    .io_e_i(array_47_io_e_i),
    .io_f_i(array_47_io_f_i),
    .io_ve_i(array_47_io_ve_i),
    .io_vf_i(array_47_io_vf_i),
    .io_vv_i(array_47_io_vv_i),
    .io_e_o(array_47_io_e_o),
    .io_f_o(array_47_io_f_o),
    .io_v_o(array_47_io_v_o)
  );
  SWCell array_48 ( // @[SWChisel.scala 170:39]
    .io_q(array_48_io_q),
    .io_r(array_48_io_r),
    .io_e_i(array_48_io_e_i),
    .io_f_i(array_48_io_f_i),
    .io_ve_i(array_48_io_ve_i),
    .io_vf_i(array_48_io_vf_i),
    .io_vv_i(array_48_io_vv_i),
    .io_e_o(array_48_io_e_o),
    .io_f_o(array_48_io_f_o),
    .io_v_o(array_48_io_v_o)
  );
  SWCell array_49 ( // @[SWChisel.scala 170:39]
    .io_q(array_49_io_q),
    .io_r(array_49_io_r),
    .io_e_i(array_49_io_e_i),
    .io_f_i(array_49_io_f_i),
    .io_ve_i(array_49_io_ve_i),
    .io_vf_i(array_49_io_vf_i),
    .io_vv_i(array_49_io_vv_i),
    .io_e_o(array_49_io_e_o),
    .io_f_o(array_49_io_f_o),
    .io_v_o(array_49_io_v_o)
  );
  SWCell array_50 ( // @[SWChisel.scala 170:39]
    .io_q(array_50_io_q),
    .io_r(array_50_io_r),
    .io_e_i(array_50_io_e_i),
    .io_f_i(array_50_io_f_i),
    .io_ve_i(array_50_io_ve_i),
    .io_vf_i(array_50_io_vf_i),
    .io_vv_i(array_50_io_vv_i),
    .io_e_o(array_50_io_e_o),
    .io_f_o(array_50_io_f_o),
    .io_v_o(array_50_io_v_o)
  );
  SWCell array_51 ( // @[SWChisel.scala 170:39]
    .io_q(array_51_io_q),
    .io_r(array_51_io_r),
    .io_e_i(array_51_io_e_i),
    .io_f_i(array_51_io_f_i),
    .io_ve_i(array_51_io_ve_i),
    .io_vf_i(array_51_io_vf_i),
    .io_vv_i(array_51_io_vv_i),
    .io_e_o(array_51_io_e_o),
    .io_f_o(array_51_io_f_o),
    .io_v_o(array_51_io_v_o)
  );
  SWCell array_52 ( // @[SWChisel.scala 170:39]
    .io_q(array_52_io_q),
    .io_r(array_52_io_r),
    .io_e_i(array_52_io_e_i),
    .io_f_i(array_52_io_f_i),
    .io_ve_i(array_52_io_ve_i),
    .io_vf_i(array_52_io_vf_i),
    .io_vv_i(array_52_io_vv_i),
    .io_e_o(array_52_io_e_o),
    .io_f_o(array_52_io_f_o),
    .io_v_o(array_52_io_v_o)
  );
  SWCell array_53 ( // @[SWChisel.scala 170:39]
    .io_q(array_53_io_q),
    .io_r(array_53_io_r),
    .io_e_i(array_53_io_e_i),
    .io_f_i(array_53_io_f_i),
    .io_ve_i(array_53_io_ve_i),
    .io_vf_i(array_53_io_vf_i),
    .io_vv_i(array_53_io_vv_i),
    .io_e_o(array_53_io_e_o),
    .io_f_o(array_53_io_f_o),
    .io_v_o(array_53_io_v_o)
  );
  SWCell array_54 ( // @[SWChisel.scala 170:39]
    .io_q(array_54_io_q),
    .io_r(array_54_io_r),
    .io_e_i(array_54_io_e_i),
    .io_f_i(array_54_io_f_i),
    .io_ve_i(array_54_io_ve_i),
    .io_vf_i(array_54_io_vf_i),
    .io_vv_i(array_54_io_vv_i),
    .io_e_o(array_54_io_e_o),
    .io_f_o(array_54_io_f_o),
    .io_v_o(array_54_io_v_o)
  );
  SWCell array_55 ( // @[SWChisel.scala 170:39]
    .io_q(array_55_io_q),
    .io_r(array_55_io_r),
    .io_e_i(array_55_io_e_i),
    .io_f_i(array_55_io_f_i),
    .io_ve_i(array_55_io_ve_i),
    .io_vf_i(array_55_io_vf_i),
    .io_vv_i(array_55_io_vv_i),
    .io_e_o(array_55_io_e_o),
    .io_f_o(array_55_io_f_o),
    .io_v_o(array_55_io_v_o)
  );
  SWCell array_56 ( // @[SWChisel.scala 170:39]
    .io_q(array_56_io_q),
    .io_r(array_56_io_r),
    .io_e_i(array_56_io_e_i),
    .io_f_i(array_56_io_f_i),
    .io_ve_i(array_56_io_ve_i),
    .io_vf_i(array_56_io_vf_i),
    .io_vv_i(array_56_io_vv_i),
    .io_e_o(array_56_io_e_o),
    .io_f_o(array_56_io_f_o),
    .io_v_o(array_56_io_v_o)
  );
  SWCell array_57 ( // @[SWChisel.scala 170:39]
    .io_q(array_57_io_q),
    .io_r(array_57_io_r),
    .io_e_i(array_57_io_e_i),
    .io_f_i(array_57_io_f_i),
    .io_ve_i(array_57_io_ve_i),
    .io_vf_i(array_57_io_vf_i),
    .io_vv_i(array_57_io_vv_i),
    .io_e_o(array_57_io_e_o),
    .io_f_o(array_57_io_f_o),
    .io_v_o(array_57_io_v_o)
  );
  SWCell array_58 ( // @[SWChisel.scala 170:39]
    .io_q(array_58_io_q),
    .io_r(array_58_io_r),
    .io_e_i(array_58_io_e_i),
    .io_f_i(array_58_io_f_i),
    .io_ve_i(array_58_io_ve_i),
    .io_vf_i(array_58_io_vf_i),
    .io_vv_i(array_58_io_vv_i),
    .io_e_o(array_58_io_e_o),
    .io_f_o(array_58_io_f_o),
    .io_v_o(array_58_io_v_o)
  );
  SWCell array_59 ( // @[SWChisel.scala 170:39]
    .io_q(array_59_io_q),
    .io_r(array_59_io_r),
    .io_e_i(array_59_io_e_i),
    .io_f_i(array_59_io_f_i),
    .io_ve_i(array_59_io_ve_i),
    .io_vf_i(array_59_io_vf_i),
    .io_vv_i(array_59_io_vv_i),
    .io_e_o(array_59_io_e_o),
    .io_f_o(array_59_io_f_o),
    .io_v_o(array_59_io_v_o)
  );
  SWCell array_60 ( // @[SWChisel.scala 170:39]
    .io_q(array_60_io_q),
    .io_r(array_60_io_r),
    .io_e_i(array_60_io_e_i),
    .io_f_i(array_60_io_f_i),
    .io_ve_i(array_60_io_ve_i),
    .io_vf_i(array_60_io_vf_i),
    .io_vv_i(array_60_io_vv_i),
    .io_e_o(array_60_io_e_o),
    .io_f_o(array_60_io_f_o),
    .io_v_o(array_60_io_v_o)
  );
  SWCell array_61 ( // @[SWChisel.scala 170:39]
    .io_q(array_61_io_q),
    .io_r(array_61_io_r),
    .io_e_i(array_61_io_e_i),
    .io_f_i(array_61_io_f_i),
    .io_ve_i(array_61_io_ve_i),
    .io_vf_i(array_61_io_vf_i),
    .io_vv_i(array_61_io_vv_i),
    .io_e_o(array_61_io_e_o),
    .io_f_o(array_61_io_f_o),
    .io_v_o(array_61_io_v_o)
  );
  SWCell array_62 ( // @[SWChisel.scala 170:39]
    .io_q(array_62_io_q),
    .io_r(array_62_io_r),
    .io_e_i(array_62_io_e_i),
    .io_f_i(array_62_io_f_i),
    .io_ve_i(array_62_io_ve_i),
    .io_vf_i(array_62_io_vf_i),
    .io_vv_i(array_62_io_vv_i),
    .io_e_o(array_62_io_e_o),
    .io_f_o(array_62_io_f_o),
    .io_v_o(array_62_io_v_o)
  );
  SWCell array_63 ( // @[SWChisel.scala 170:39]
    .io_q(array_63_io_q),
    .io_r(array_63_io_r),
    .io_e_i(array_63_io_e_i),
    .io_f_i(array_63_io_f_i),
    .io_ve_i(array_63_io_ve_i),
    .io_vf_i(array_63_io_vf_i),
    .io_vv_i(array_63_io_vv_i),
    .io_e_o(array_63_io_e_o),
    .io_f_o(array_63_io_f_o),
    .io_v_o(array_63_io_v_o)
  );
  SWCell array_64 ( // @[SWChisel.scala 170:39]
    .io_q(array_64_io_q),
    .io_r(array_64_io_r),
    .io_e_i(array_64_io_e_i),
    .io_f_i(array_64_io_f_i),
    .io_ve_i(array_64_io_ve_i),
    .io_vf_i(array_64_io_vf_i),
    .io_vv_i(array_64_io_vv_i),
    .io_e_o(array_64_io_e_o),
    .io_f_o(array_64_io_f_o),
    .io_v_o(array_64_io_v_o)
  );
  SWCell array_65 ( // @[SWChisel.scala 170:39]
    .io_q(array_65_io_q),
    .io_r(array_65_io_r),
    .io_e_i(array_65_io_e_i),
    .io_f_i(array_65_io_f_i),
    .io_ve_i(array_65_io_ve_i),
    .io_vf_i(array_65_io_vf_i),
    .io_vv_i(array_65_io_vv_i),
    .io_e_o(array_65_io_e_o),
    .io_f_o(array_65_io_f_o),
    .io_v_o(array_65_io_v_o)
  );
  SWCell array_66 ( // @[SWChisel.scala 170:39]
    .io_q(array_66_io_q),
    .io_r(array_66_io_r),
    .io_e_i(array_66_io_e_i),
    .io_f_i(array_66_io_f_i),
    .io_ve_i(array_66_io_ve_i),
    .io_vf_i(array_66_io_vf_i),
    .io_vv_i(array_66_io_vv_i),
    .io_e_o(array_66_io_e_o),
    .io_f_o(array_66_io_f_o),
    .io_v_o(array_66_io_v_o)
  );
  SWCell array_67 ( // @[SWChisel.scala 170:39]
    .io_q(array_67_io_q),
    .io_r(array_67_io_r),
    .io_e_i(array_67_io_e_i),
    .io_f_i(array_67_io_f_i),
    .io_ve_i(array_67_io_ve_i),
    .io_vf_i(array_67_io_vf_i),
    .io_vv_i(array_67_io_vv_i),
    .io_e_o(array_67_io_e_o),
    .io_f_o(array_67_io_f_o),
    .io_v_o(array_67_io_v_o)
  );
  SWCell array_68 ( // @[SWChisel.scala 170:39]
    .io_q(array_68_io_q),
    .io_r(array_68_io_r),
    .io_e_i(array_68_io_e_i),
    .io_f_i(array_68_io_f_i),
    .io_ve_i(array_68_io_ve_i),
    .io_vf_i(array_68_io_vf_i),
    .io_vv_i(array_68_io_vv_i),
    .io_e_o(array_68_io_e_o),
    .io_f_o(array_68_io_f_o),
    .io_v_o(array_68_io_v_o)
  );
  SWCell array_69 ( // @[SWChisel.scala 170:39]
    .io_q(array_69_io_q),
    .io_r(array_69_io_r),
    .io_e_i(array_69_io_e_i),
    .io_f_i(array_69_io_f_i),
    .io_ve_i(array_69_io_ve_i),
    .io_vf_i(array_69_io_vf_i),
    .io_vv_i(array_69_io_vv_i),
    .io_e_o(array_69_io_e_o),
    .io_f_o(array_69_io_f_o),
    .io_v_o(array_69_io_v_o)
  );
  SWCell array_70 ( // @[SWChisel.scala 170:39]
    .io_q(array_70_io_q),
    .io_r(array_70_io_r),
    .io_e_i(array_70_io_e_i),
    .io_f_i(array_70_io_f_i),
    .io_ve_i(array_70_io_ve_i),
    .io_vf_i(array_70_io_vf_i),
    .io_vv_i(array_70_io_vv_i),
    .io_e_o(array_70_io_e_o),
    .io_f_o(array_70_io_f_o),
    .io_v_o(array_70_io_v_o)
  );
  SWCell array_71 ( // @[SWChisel.scala 170:39]
    .io_q(array_71_io_q),
    .io_r(array_71_io_r),
    .io_e_i(array_71_io_e_i),
    .io_f_i(array_71_io_f_i),
    .io_ve_i(array_71_io_ve_i),
    .io_vf_i(array_71_io_vf_i),
    .io_vv_i(array_71_io_vv_i),
    .io_e_o(array_71_io_e_o),
    .io_f_o(array_71_io_f_o),
    .io_v_o(array_71_io_v_o)
  );
  SWCell array_72 ( // @[SWChisel.scala 170:39]
    .io_q(array_72_io_q),
    .io_r(array_72_io_r),
    .io_e_i(array_72_io_e_i),
    .io_f_i(array_72_io_f_i),
    .io_ve_i(array_72_io_ve_i),
    .io_vf_i(array_72_io_vf_i),
    .io_vv_i(array_72_io_vv_i),
    .io_e_o(array_72_io_e_o),
    .io_f_o(array_72_io_f_o),
    .io_v_o(array_72_io_v_o)
  );
  SWCell array_73 ( // @[SWChisel.scala 170:39]
    .io_q(array_73_io_q),
    .io_r(array_73_io_r),
    .io_e_i(array_73_io_e_i),
    .io_f_i(array_73_io_f_i),
    .io_ve_i(array_73_io_ve_i),
    .io_vf_i(array_73_io_vf_i),
    .io_vv_i(array_73_io_vv_i),
    .io_e_o(array_73_io_e_o),
    .io_f_o(array_73_io_f_o),
    .io_v_o(array_73_io_v_o)
  );
  SWCell array_74 ( // @[SWChisel.scala 170:39]
    .io_q(array_74_io_q),
    .io_r(array_74_io_r),
    .io_e_i(array_74_io_e_i),
    .io_f_i(array_74_io_f_i),
    .io_ve_i(array_74_io_ve_i),
    .io_vf_i(array_74_io_vf_i),
    .io_vv_i(array_74_io_vv_i),
    .io_e_o(array_74_io_e_o),
    .io_f_o(array_74_io_f_o),
    .io_v_o(array_74_io_v_o)
  );
  SWCell array_75 ( // @[SWChisel.scala 170:39]
    .io_q(array_75_io_q),
    .io_r(array_75_io_r),
    .io_e_i(array_75_io_e_i),
    .io_f_i(array_75_io_f_i),
    .io_ve_i(array_75_io_ve_i),
    .io_vf_i(array_75_io_vf_i),
    .io_vv_i(array_75_io_vv_i),
    .io_e_o(array_75_io_e_o),
    .io_f_o(array_75_io_f_o),
    .io_v_o(array_75_io_v_o)
  );
  SWCell array_76 ( // @[SWChisel.scala 170:39]
    .io_q(array_76_io_q),
    .io_r(array_76_io_r),
    .io_e_i(array_76_io_e_i),
    .io_f_i(array_76_io_f_i),
    .io_ve_i(array_76_io_ve_i),
    .io_vf_i(array_76_io_vf_i),
    .io_vv_i(array_76_io_vv_i),
    .io_e_o(array_76_io_e_o),
    .io_f_o(array_76_io_f_o),
    .io_v_o(array_76_io_v_o)
  );
  SWCell array_77 ( // @[SWChisel.scala 170:39]
    .io_q(array_77_io_q),
    .io_r(array_77_io_r),
    .io_e_i(array_77_io_e_i),
    .io_f_i(array_77_io_f_i),
    .io_ve_i(array_77_io_ve_i),
    .io_vf_i(array_77_io_vf_i),
    .io_vv_i(array_77_io_vv_i),
    .io_e_o(array_77_io_e_o),
    .io_f_o(array_77_io_f_o),
    .io_v_o(array_77_io_v_o)
  );
  SWCell array_78 ( // @[SWChisel.scala 170:39]
    .io_q(array_78_io_q),
    .io_r(array_78_io_r),
    .io_e_i(array_78_io_e_i),
    .io_f_i(array_78_io_f_i),
    .io_ve_i(array_78_io_ve_i),
    .io_vf_i(array_78_io_vf_i),
    .io_vv_i(array_78_io_vv_i),
    .io_e_o(array_78_io_e_o),
    .io_f_o(array_78_io_f_o),
    .io_v_o(array_78_io_v_o)
  );
  SWCell array_79 ( // @[SWChisel.scala 170:39]
    .io_q(array_79_io_q),
    .io_r(array_79_io_r),
    .io_e_i(array_79_io_e_i),
    .io_f_i(array_79_io_f_i),
    .io_ve_i(array_79_io_ve_i),
    .io_vf_i(array_79_io_vf_i),
    .io_vv_i(array_79_io_vv_i),
    .io_e_o(array_79_io_e_o),
    .io_f_o(array_79_io_f_o),
    .io_v_o(array_79_io_v_o)
  );
  SWCell array_80 ( // @[SWChisel.scala 170:39]
    .io_q(array_80_io_q),
    .io_r(array_80_io_r),
    .io_e_i(array_80_io_e_i),
    .io_f_i(array_80_io_f_i),
    .io_ve_i(array_80_io_ve_i),
    .io_vf_i(array_80_io_vf_i),
    .io_vv_i(array_80_io_vv_i),
    .io_e_o(array_80_io_e_o),
    .io_f_o(array_80_io_f_o),
    .io_v_o(array_80_io_v_o)
  );
  SWCell array_81 ( // @[SWChisel.scala 170:39]
    .io_q(array_81_io_q),
    .io_r(array_81_io_r),
    .io_e_i(array_81_io_e_i),
    .io_f_i(array_81_io_f_i),
    .io_ve_i(array_81_io_ve_i),
    .io_vf_i(array_81_io_vf_i),
    .io_vv_i(array_81_io_vv_i),
    .io_e_o(array_81_io_e_o),
    .io_f_o(array_81_io_f_o),
    .io_v_o(array_81_io_v_o)
  );
  SWCell array_82 ( // @[SWChisel.scala 170:39]
    .io_q(array_82_io_q),
    .io_r(array_82_io_r),
    .io_e_i(array_82_io_e_i),
    .io_f_i(array_82_io_f_i),
    .io_ve_i(array_82_io_ve_i),
    .io_vf_i(array_82_io_vf_i),
    .io_vv_i(array_82_io_vv_i),
    .io_e_o(array_82_io_e_o),
    .io_f_o(array_82_io_f_o),
    .io_v_o(array_82_io_v_o)
  );
  SWCell array_83 ( // @[SWChisel.scala 170:39]
    .io_q(array_83_io_q),
    .io_r(array_83_io_r),
    .io_e_i(array_83_io_e_i),
    .io_f_i(array_83_io_f_i),
    .io_ve_i(array_83_io_ve_i),
    .io_vf_i(array_83_io_vf_i),
    .io_vv_i(array_83_io_vv_i),
    .io_e_o(array_83_io_e_o),
    .io_f_o(array_83_io_f_o),
    .io_v_o(array_83_io_v_o)
  );
  SWCell array_84 ( // @[SWChisel.scala 170:39]
    .io_q(array_84_io_q),
    .io_r(array_84_io_r),
    .io_e_i(array_84_io_e_i),
    .io_f_i(array_84_io_f_i),
    .io_ve_i(array_84_io_ve_i),
    .io_vf_i(array_84_io_vf_i),
    .io_vv_i(array_84_io_vv_i),
    .io_e_o(array_84_io_e_o),
    .io_f_o(array_84_io_f_o),
    .io_v_o(array_84_io_v_o)
  );
  SWCell array_85 ( // @[SWChisel.scala 170:39]
    .io_q(array_85_io_q),
    .io_r(array_85_io_r),
    .io_e_i(array_85_io_e_i),
    .io_f_i(array_85_io_f_i),
    .io_ve_i(array_85_io_ve_i),
    .io_vf_i(array_85_io_vf_i),
    .io_vv_i(array_85_io_vv_i),
    .io_e_o(array_85_io_e_o),
    .io_f_o(array_85_io_f_o),
    .io_v_o(array_85_io_v_o)
  );
  SWCell array_86 ( // @[SWChisel.scala 170:39]
    .io_q(array_86_io_q),
    .io_r(array_86_io_r),
    .io_e_i(array_86_io_e_i),
    .io_f_i(array_86_io_f_i),
    .io_ve_i(array_86_io_ve_i),
    .io_vf_i(array_86_io_vf_i),
    .io_vv_i(array_86_io_vv_i),
    .io_e_o(array_86_io_e_o),
    .io_f_o(array_86_io_f_o),
    .io_v_o(array_86_io_v_o)
  );
  SWCell array_87 ( // @[SWChisel.scala 170:39]
    .io_q(array_87_io_q),
    .io_r(array_87_io_r),
    .io_e_i(array_87_io_e_i),
    .io_f_i(array_87_io_f_i),
    .io_ve_i(array_87_io_ve_i),
    .io_vf_i(array_87_io_vf_i),
    .io_vv_i(array_87_io_vv_i),
    .io_e_o(array_87_io_e_o),
    .io_f_o(array_87_io_f_o),
    .io_v_o(array_87_io_v_o)
  );
  SWCell array_88 ( // @[SWChisel.scala 170:39]
    .io_q(array_88_io_q),
    .io_r(array_88_io_r),
    .io_e_i(array_88_io_e_i),
    .io_f_i(array_88_io_f_i),
    .io_ve_i(array_88_io_ve_i),
    .io_vf_i(array_88_io_vf_i),
    .io_vv_i(array_88_io_vv_i),
    .io_e_o(array_88_io_e_o),
    .io_f_o(array_88_io_f_o),
    .io_v_o(array_88_io_v_o)
  );
  SWCell array_89 ( // @[SWChisel.scala 170:39]
    .io_q(array_89_io_q),
    .io_r(array_89_io_r),
    .io_e_i(array_89_io_e_i),
    .io_f_i(array_89_io_f_i),
    .io_ve_i(array_89_io_ve_i),
    .io_vf_i(array_89_io_vf_i),
    .io_vv_i(array_89_io_vv_i),
    .io_e_o(array_89_io_e_o),
    .io_f_o(array_89_io_f_o),
    .io_v_o(array_89_io_v_o)
  );
  SWCell array_90 ( // @[SWChisel.scala 170:39]
    .io_q(array_90_io_q),
    .io_r(array_90_io_r),
    .io_e_i(array_90_io_e_i),
    .io_f_i(array_90_io_f_i),
    .io_ve_i(array_90_io_ve_i),
    .io_vf_i(array_90_io_vf_i),
    .io_vv_i(array_90_io_vv_i),
    .io_e_o(array_90_io_e_o),
    .io_f_o(array_90_io_f_o),
    .io_v_o(array_90_io_v_o)
  );
  SWCell array_91 ( // @[SWChisel.scala 170:39]
    .io_q(array_91_io_q),
    .io_r(array_91_io_r),
    .io_e_i(array_91_io_e_i),
    .io_f_i(array_91_io_f_i),
    .io_ve_i(array_91_io_ve_i),
    .io_vf_i(array_91_io_vf_i),
    .io_vv_i(array_91_io_vv_i),
    .io_e_o(array_91_io_e_o),
    .io_f_o(array_91_io_f_o),
    .io_v_o(array_91_io_v_o)
  );
  SWCell array_92 ( // @[SWChisel.scala 170:39]
    .io_q(array_92_io_q),
    .io_r(array_92_io_r),
    .io_e_i(array_92_io_e_i),
    .io_f_i(array_92_io_f_i),
    .io_ve_i(array_92_io_ve_i),
    .io_vf_i(array_92_io_vf_i),
    .io_vv_i(array_92_io_vv_i),
    .io_e_o(array_92_io_e_o),
    .io_f_o(array_92_io_f_o),
    .io_v_o(array_92_io_v_o)
  );
  SWCell array_93 ( // @[SWChisel.scala 170:39]
    .io_q(array_93_io_q),
    .io_r(array_93_io_r),
    .io_e_i(array_93_io_e_i),
    .io_f_i(array_93_io_f_i),
    .io_ve_i(array_93_io_ve_i),
    .io_vf_i(array_93_io_vf_i),
    .io_vv_i(array_93_io_vv_i),
    .io_e_o(array_93_io_e_o),
    .io_f_o(array_93_io_f_o),
    .io_v_o(array_93_io_v_o)
  );
  SWCell array_94 ( // @[SWChisel.scala 170:39]
    .io_q(array_94_io_q),
    .io_r(array_94_io_r),
    .io_e_i(array_94_io_e_i),
    .io_f_i(array_94_io_f_i),
    .io_ve_i(array_94_io_ve_i),
    .io_vf_i(array_94_io_vf_i),
    .io_vv_i(array_94_io_vv_i),
    .io_e_o(array_94_io_e_o),
    .io_f_o(array_94_io_f_o),
    .io_v_o(array_94_io_v_o)
  );
  SWCell array_95 ( // @[SWChisel.scala 170:39]
    .io_q(array_95_io_q),
    .io_r(array_95_io_r),
    .io_e_i(array_95_io_e_i),
    .io_f_i(array_95_io_f_i),
    .io_ve_i(array_95_io_ve_i),
    .io_vf_i(array_95_io_vf_i),
    .io_vv_i(array_95_io_vv_i),
    .io_e_o(array_95_io_e_o),
    .io_f_o(array_95_io_f_o),
    .io_v_o(array_95_io_v_o)
  );
  SWCell array_96 ( // @[SWChisel.scala 170:39]
    .io_q(array_96_io_q),
    .io_r(array_96_io_r),
    .io_e_i(array_96_io_e_i),
    .io_f_i(array_96_io_f_i),
    .io_ve_i(array_96_io_ve_i),
    .io_vf_i(array_96_io_vf_i),
    .io_vv_i(array_96_io_vv_i),
    .io_e_o(array_96_io_e_o),
    .io_f_o(array_96_io_f_o),
    .io_v_o(array_96_io_v_o)
  );
  SWCell array_97 ( // @[SWChisel.scala 170:39]
    .io_q(array_97_io_q),
    .io_r(array_97_io_r),
    .io_e_i(array_97_io_e_i),
    .io_f_i(array_97_io_f_i),
    .io_ve_i(array_97_io_ve_i),
    .io_vf_i(array_97_io_vf_i),
    .io_vv_i(array_97_io_vv_i),
    .io_e_o(array_97_io_e_o),
    .io_f_o(array_97_io_f_o),
    .io_v_o(array_97_io_v_o)
  );
  SWCell array_98 ( // @[SWChisel.scala 170:39]
    .io_q(array_98_io_q),
    .io_r(array_98_io_r),
    .io_e_i(array_98_io_e_i),
    .io_f_i(array_98_io_f_i),
    .io_ve_i(array_98_io_ve_i),
    .io_vf_i(array_98_io_vf_i),
    .io_vv_i(array_98_io_vv_i),
    .io_e_o(array_98_io_e_o),
    .io_f_o(array_98_io_f_o),
    .io_v_o(array_98_io_v_o)
  );
  SWCell array_99 ( // @[SWChisel.scala 170:39]
    .io_q(array_99_io_q),
    .io_r(array_99_io_r),
    .io_e_i(array_99_io_e_i),
    .io_f_i(array_99_io_f_i),
    .io_ve_i(array_99_io_ve_i),
    .io_vf_i(array_99_io_vf_i),
    .io_vv_i(array_99_io_vv_i),
    .io_e_o(array_99_io_e_o),
    .io_f_o(array_99_io_f_o),
    .io_v_o(array_99_io_v_o)
  );
  MyCounter r_count_0 ( // @[SWChisel.scala 171:41]
    .clock(r_count_0_clock),
    .reset(r_count_0_reset),
    .io_en(r_count_0_io_en),
    .io_out(r_count_0_io_out)
  );
  MyCounter r_count_1 ( // @[SWChisel.scala 171:41]
    .clock(r_count_1_clock),
    .reset(r_count_1_reset),
    .io_en(r_count_1_io_en),
    .io_out(r_count_1_io_out)
  );
  MyCounter r_count_2 ( // @[SWChisel.scala 171:41]
    .clock(r_count_2_clock),
    .reset(r_count_2_reset),
    .io_en(r_count_2_io_en),
    .io_out(r_count_2_io_out)
  );
  MyCounter r_count_3 ( // @[SWChisel.scala 171:41]
    .clock(r_count_3_clock),
    .reset(r_count_3_reset),
    .io_en(r_count_3_io_en),
    .io_out(r_count_3_io_out)
  );
  MyCounter r_count_4 ( // @[SWChisel.scala 171:41]
    .clock(r_count_4_clock),
    .reset(r_count_4_reset),
    .io_en(r_count_4_io_en),
    .io_out(r_count_4_io_out)
  );
  MyCounter r_count_5 ( // @[SWChisel.scala 171:41]
    .clock(r_count_5_clock),
    .reset(r_count_5_reset),
    .io_en(r_count_5_io_en),
    .io_out(r_count_5_io_out)
  );
  MyCounter r_count_6 ( // @[SWChisel.scala 171:41]
    .clock(r_count_6_clock),
    .reset(r_count_6_reset),
    .io_en(r_count_6_io_en),
    .io_out(r_count_6_io_out)
  );
  MyCounter r_count_7 ( // @[SWChisel.scala 171:41]
    .clock(r_count_7_clock),
    .reset(r_count_7_reset),
    .io_en(r_count_7_io_en),
    .io_out(r_count_7_io_out)
  );
  MyCounter r_count_8 ( // @[SWChisel.scala 171:41]
    .clock(r_count_8_clock),
    .reset(r_count_8_reset),
    .io_en(r_count_8_io_en),
    .io_out(r_count_8_io_out)
  );
  MyCounter r_count_9 ( // @[SWChisel.scala 171:41]
    .clock(r_count_9_clock),
    .reset(r_count_9_reset),
    .io_en(r_count_9_io_en),
    .io_out(r_count_9_io_out)
  );
  MyCounter r_count_10 ( // @[SWChisel.scala 171:41]
    .clock(r_count_10_clock),
    .reset(r_count_10_reset),
    .io_en(r_count_10_io_en),
    .io_out(r_count_10_io_out)
  );
  MyCounter r_count_11 ( // @[SWChisel.scala 171:41]
    .clock(r_count_11_clock),
    .reset(r_count_11_reset),
    .io_en(r_count_11_io_en),
    .io_out(r_count_11_io_out)
  );
  MyCounter r_count_12 ( // @[SWChisel.scala 171:41]
    .clock(r_count_12_clock),
    .reset(r_count_12_reset),
    .io_en(r_count_12_io_en),
    .io_out(r_count_12_io_out)
  );
  MyCounter r_count_13 ( // @[SWChisel.scala 171:41]
    .clock(r_count_13_clock),
    .reset(r_count_13_reset),
    .io_en(r_count_13_io_en),
    .io_out(r_count_13_io_out)
  );
  MyCounter r_count_14 ( // @[SWChisel.scala 171:41]
    .clock(r_count_14_clock),
    .reset(r_count_14_reset),
    .io_en(r_count_14_io_en),
    .io_out(r_count_14_io_out)
  );
  MyCounter r_count_15 ( // @[SWChisel.scala 171:41]
    .clock(r_count_15_clock),
    .reset(r_count_15_reset),
    .io_en(r_count_15_io_en),
    .io_out(r_count_15_io_out)
  );
  MyCounter r_count_16 ( // @[SWChisel.scala 171:41]
    .clock(r_count_16_clock),
    .reset(r_count_16_reset),
    .io_en(r_count_16_io_en),
    .io_out(r_count_16_io_out)
  );
  MyCounter r_count_17 ( // @[SWChisel.scala 171:41]
    .clock(r_count_17_clock),
    .reset(r_count_17_reset),
    .io_en(r_count_17_io_en),
    .io_out(r_count_17_io_out)
  );
  MyCounter r_count_18 ( // @[SWChisel.scala 171:41]
    .clock(r_count_18_clock),
    .reset(r_count_18_reset),
    .io_en(r_count_18_io_en),
    .io_out(r_count_18_io_out)
  );
  MyCounter r_count_19 ( // @[SWChisel.scala 171:41]
    .clock(r_count_19_clock),
    .reset(r_count_19_reset),
    .io_en(r_count_19_io_en),
    .io_out(r_count_19_io_out)
  );
  MyCounter r_count_20 ( // @[SWChisel.scala 171:41]
    .clock(r_count_20_clock),
    .reset(r_count_20_reset),
    .io_en(r_count_20_io_en),
    .io_out(r_count_20_io_out)
  );
  MyCounter r_count_21 ( // @[SWChisel.scala 171:41]
    .clock(r_count_21_clock),
    .reset(r_count_21_reset),
    .io_en(r_count_21_io_en),
    .io_out(r_count_21_io_out)
  );
  MyCounter r_count_22 ( // @[SWChisel.scala 171:41]
    .clock(r_count_22_clock),
    .reset(r_count_22_reset),
    .io_en(r_count_22_io_en),
    .io_out(r_count_22_io_out)
  );
  MyCounter r_count_23 ( // @[SWChisel.scala 171:41]
    .clock(r_count_23_clock),
    .reset(r_count_23_reset),
    .io_en(r_count_23_io_en),
    .io_out(r_count_23_io_out)
  );
  MyCounter r_count_24 ( // @[SWChisel.scala 171:41]
    .clock(r_count_24_clock),
    .reset(r_count_24_reset),
    .io_en(r_count_24_io_en),
    .io_out(r_count_24_io_out)
  );
  MyCounter r_count_25 ( // @[SWChisel.scala 171:41]
    .clock(r_count_25_clock),
    .reset(r_count_25_reset),
    .io_en(r_count_25_io_en),
    .io_out(r_count_25_io_out)
  );
  MyCounter r_count_26 ( // @[SWChisel.scala 171:41]
    .clock(r_count_26_clock),
    .reset(r_count_26_reset),
    .io_en(r_count_26_io_en),
    .io_out(r_count_26_io_out)
  );
  MyCounter r_count_27 ( // @[SWChisel.scala 171:41]
    .clock(r_count_27_clock),
    .reset(r_count_27_reset),
    .io_en(r_count_27_io_en),
    .io_out(r_count_27_io_out)
  );
  MyCounter r_count_28 ( // @[SWChisel.scala 171:41]
    .clock(r_count_28_clock),
    .reset(r_count_28_reset),
    .io_en(r_count_28_io_en),
    .io_out(r_count_28_io_out)
  );
  MyCounter r_count_29 ( // @[SWChisel.scala 171:41]
    .clock(r_count_29_clock),
    .reset(r_count_29_reset),
    .io_en(r_count_29_io_en),
    .io_out(r_count_29_io_out)
  );
  MyCounter r_count_30 ( // @[SWChisel.scala 171:41]
    .clock(r_count_30_clock),
    .reset(r_count_30_reset),
    .io_en(r_count_30_io_en),
    .io_out(r_count_30_io_out)
  );
  MyCounter r_count_31 ( // @[SWChisel.scala 171:41]
    .clock(r_count_31_clock),
    .reset(r_count_31_reset),
    .io_en(r_count_31_io_en),
    .io_out(r_count_31_io_out)
  );
  MyCounter r_count_32 ( // @[SWChisel.scala 171:41]
    .clock(r_count_32_clock),
    .reset(r_count_32_reset),
    .io_en(r_count_32_io_en),
    .io_out(r_count_32_io_out)
  );
  MyCounter r_count_33 ( // @[SWChisel.scala 171:41]
    .clock(r_count_33_clock),
    .reset(r_count_33_reset),
    .io_en(r_count_33_io_en),
    .io_out(r_count_33_io_out)
  );
  MyCounter r_count_34 ( // @[SWChisel.scala 171:41]
    .clock(r_count_34_clock),
    .reset(r_count_34_reset),
    .io_en(r_count_34_io_en),
    .io_out(r_count_34_io_out)
  );
  MyCounter r_count_35 ( // @[SWChisel.scala 171:41]
    .clock(r_count_35_clock),
    .reset(r_count_35_reset),
    .io_en(r_count_35_io_en),
    .io_out(r_count_35_io_out)
  );
  MyCounter r_count_36 ( // @[SWChisel.scala 171:41]
    .clock(r_count_36_clock),
    .reset(r_count_36_reset),
    .io_en(r_count_36_io_en),
    .io_out(r_count_36_io_out)
  );
  MyCounter r_count_37 ( // @[SWChisel.scala 171:41]
    .clock(r_count_37_clock),
    .reset(r_count_37_reset),
    .io_en(r_count_37_io_en),
    .io_out(r_count_37_io_out)
  );
  MyCounter r_count_38 ( // @[SWChisel.scala 171:41]
    .clock(r_count_38_clock),
    .reset(r_count_38_reset),
    .io_en(r_count_38_io_en),
    .io_out(r_count_38_io_out)
  );
  MyCounter r_count_39 ( // @[SWChisel.scala 171:41]
    .clock(r_count_39_clock),
    .reset(r_count_39_reset),
    .io_en(r_count_39_io_en),
    .io_out(r_count_39_io_out)
  );
  MyCounter r_count_40 ( // @[SWChisel.scala 171:41]
    .clock(r_count_40_clock),
    .reset(r_count_40_reset),
    .io_en(r_count_40_io_en),
    .io_out(r_count_40_io_out)
  );
  MyCounter r_count_41 ( // @[SWChisel.scala 171:41]
    .clock(r_count_41_clock),
    .reset(r_count_41_reset),
    .io_en(r_count_41_io_en),
    .io_out(r_count_41_io_out)
  );
  MyCounter r_count_42 ( // @[SWChisel.scala 171:41]
    .clock(r_count_42_clock),
    .reset(r_count_42_reset),
    .io_en(r_count_42_io_en),
    .io_out(r_count_42_io_out)
  );
  MyCounter r_count_43 ( // @[SWChisel.scala 171:41]
    .clock(r_count_43_clock),
    .reset(r_count_43_reset),
    .io_en(r_count_43_io_en),
    .io_out(r_count_43_io_out)
  );
  MyCounter r_count_44 ( // @[SWChisel.scala 171:41]
    .clock(r_count_44_clock),
    .reset(r_count_44_reset),
    .io_en(r_count_44_io_en),
    .io_out(r_count_44_io_out)
  );
  MyCounter r_count_45 ( // @[SWChisel.scala 171:41]
    .clock(r_count_45_clock),
    .reset(r_count_45_reset),
    .io_en(r_count_45_io_en),
    .io_out(r_count_45_io_out)
  );
  MyCounter r_count_46 ( // @[SWChisel.scala 171:41]
    .clock(r_count_46_clock),
    .reset(r_count_46_reset),
    .io_en(r_count_46_io_en),
    .io_out(r_count_46_io_out)
  );
  MyCounter r_count_47 ( // @[SWChisel.scala 171:41]
    .clock(r_count_47_clock),
    .reset(r_count_47_reset),
    .io_en(r_count_47_io_en),
    .io_out(r_count_47_io_out)
  );
  MyCounter r_count_48 ( // @[SWChisel.scala 171:41]
    .clock(r_count_48_clock),
    .reset(r_count_48_reset),
    .io_en(r_count_48_io_en),
    .io_out(r_count_48_io_out)
  );
  MyCounter r_count_49 ( // @[SWChisel.scala 171:41]
    .clock(r_count_49_clock),
    .reset(r_count_49_reset),
    .io_en(r_count_49_io_en),
    .io_out(r_count_49_io_out)
  );
  MyCounter r_count_50 ( // @[SWChisel.scala 171:41]
    .clock(r_count_50_clock),
    .reset(r_count_50_reset),
    .io_en(r_count_50_io_en),
    .io_out(r_count_50_io_out)
  );
  MyCounter r_count_51 ( // @[SWChisel.scala 171:41]
    .clock(r_count_51_clock),
    .reset(r_count_51_reset),
    .io_en(r_count_51_io_en),
    .io_out(r_count_51_io_out)
  );
  MyCounter r_count_52 ( // @[SWChisel.scala 171:41]
    .clock(r_count_52_clock),
    .reset(r_count_52_reset),
    .io_en(r_count_52_io_en),
    .io_out(r_count_52_io_out)
  );
  MyCounter r_count_53 ( // @[SWChisel.scala 171:41]
    .clock(r_count_53_clock),
    .reset(r_count_53_reset),
    .io_en(r_count_53_io_en),
    .io_out(r_count_53_io_out)
  );
  MyCounter r_count_54 ( // @[SWChisel.scala 171:41]
    .clock(r_count_54_clock),
    .reset(r_count_54_reset),
    .io_en(r_count_54_io_en),
    .io_out(r_count_54_io_out)
  );
  MyCounter r_count_55 ( // @[SWChisel.scala 171:41]
    .clock(r_count_55_clock),
    .reset(r_count_55_reset),
    .io_en(r_count_55_io_en),
    .io_out(r_count_55_io_out)
  );
  MyCounter r_count_56 ( // @[SWChisel.scala 171:41]
    .clock(r_count_56_clock),
    .reset(r_count_56_reset),
    .io_en(r_count_56_io_en),
    .io_out(r_count_56_io_out)
  );
  MyCounter r_count_57 ( // @[SWChisel.scala 171:41]
    .clock(r_count_57_clock),
    .reset(r_count_57_reset),
    .io_en(r_count_57_io_en),
    .io_out(r_count_57_io_out)
  );
  MyCounter r_count_58 ( // @[SWChisel.scala 171:41]
    .clock(r_count_58_clock),
    .reset(r_count_58_reset),
    .io_en(r_count_58_io_en),
    .io_out(r_count_58_io_out)
  );
  MyCounter r_count_59 ( // @[SWChisel.scala 171:41]
    .clock(r_count_59_clock),
    .reset(r_count_59_reset),
    .io_en(r_count_59_io_en),
    .io_out(r_count_59_io_out)
  );
  MyCounter r_count_60 ( // @[SWChisel.scala 171:41]
    .clock(r_count_60_clock),
    .reset(r_count_60_reset),
    .io_en(r_count_60_io_en),
    .io_out(r_count_60_io_out)
  );
  MyCounter r_count_61 ( // @[SWChisel.scala 171:41]
    .clock(r_count_61_clock),
    .reset(r_count_61_reset),
    .io_en(r_count_61_io_en),
    .io_out(r_count_61_io_out)
  );
  MyCounter r_count_62 ( // @[SWChisel.scala 171:41]
    .clock(r_count_62_clock),
    .reset(r_count_62_reset),
    .io_en(r_count_62_io_en),
    .io_out(r_count_62_io_out)
  );
  MyCounter r_count_63 ( // @[SWChisel.scala 171:41]
    .clock(r_count_63_clock),
    .reset(r_count_63_reset),
    .io_en(r_count_63_io_en),
    .io_out(r_count_63_io_out)
  );
  MyCounter r_count_64 ( // @[SWChisel.scala 171:41]
    .clock(r_count_64_clock),
    .reset(r_count_64_reset),
    .io_en(r_count_64_io_en),
    .io_out(r_count_64_io_out)
  );
  MyCounter r_count_65 ( // @[SWChisel.scala 171:41]
    .clock(r_count_65_clock),
    .reset(r_count_65_reset),
    .io_en(r_count_65_io_en),
    .io_out(r_count_65_io_out)
  );
  MyCounter r_count_66 ( // @[SWChisel.scala 171:41]
    .clock(r_count_66_clock),
    .reset(r_count_66_reset),
    .io_en(r_count_66_io_en),
    .io_out(r_count_66_io_out)
  );
  MyCounter r_count_67 ( // @[SWChisel.scala 171:41]
    .clock(r_count_67_clock),
    .reset(r_count_67_reset),
    .io_en(r_count_67_io_en),
    .io_out(r_count_67_io_out)
  );
  MyCounter r_count_68 ( // @[SWChisel.scala 171:41]
    .clock(r_count_68_clock),
    .reset(r_count_68_reset),
    .io_en(r_count_68_io_en),
    .io_out(r_count_68_io_out)
  );
  MyCounter r_count_69 ( // @[SWChisel.scala 171:41]
    .clock(r_count_69_clock),
    .reset(r_count_69_reset),
    .io_en(r_count_69_io_en),
    .io_out(r_count_69_io_out)
  );
  MyCounter r_count_70 ( // @[SWChisel.scala 171:41]
    .clock(r_count_70_clock),
    .reset(r_count_70_reset),
    .io_en(r_count_70_io_en),
    .io_out(r_count_70_io_out)
  );
  MyCounter r_count_71 ( // @[SWChisel.scala 171:41]
    .clock(r_count_71_clock),
    .reset(r_count_71_reset),
    .io_en(r_count_71_io_en),
    .io_out(r_count_71_io_out)
  );
  MyCounter r_count_72 ( // @[SWChisel.scala 171:41]
    .clock(r_count_72_clock),
    .reset(r_count_72_reset),
    .io_en(r_count_72_io_en),
    .io_out(r_count_72_io_out)
  );
  MyCounter r_count_73 ( // @[SWChisel.scala 171:41]
    .clock(r_count_73_clock),
    .reset(r_count_73_reset),
    .io_en(r_count_73_io_en),
    .io_out(r_count_73_io_out)
  );
  MyCounter r_count_74 ( // @[SWChisel.scala 171:41]
    .clock(r_count_74_clock),
    .reset(r_count_74_reset),
    .io_en(r_count_74_io_en),
    .io_out(r_count_74_io_out)
  );
  MyCounter r_count_75 ( // @[SWChisel.scala 171:41]
    .clock(r_count_75_clock),
    .reset(r_count_75_reset),
    .io_en(r_count_75_io_en),
    .io_out(r_count_75_io_out)
  );
  MyCounter r_count_76 ( // @[SWChisel.scala 171:41]
    .clock(r_count_76_clock),
    .reset(r_count_76_reset),
    .io_en(r_count_76_io_en),
    .io_out(r_count_76_io_out)
  );
  MyCounter r_count_77 ( // @[SWChisel.scala 171:41]
    .clock(r_count_77_clock),
    .reset(r_count_77_reset),
    .io_en(r_count_77_io_en),
    .io_out(r_count_77_io_out)
  );
  MyCounter r_count_78 ( // @[SWChisel.scala 171:41]
    .clock(r_count_78_clock),
    .reset(r_count_78_reset),
    .io_en(r_count_78_io_en),
    .io_out(r_count_78_io_out)
  );
  MyCounter r_count_79 ( // @[SWChisel.scala 171:41]
    .clock(r_count_79_clock),
    .reset(r_count_79_reset),
    .io_en(r_count_79_io_en),
    .io_out(r_count_79_io_out)
  );
  MyCounter r_count_80 ( // @[SWChisel.scala 171:41]
    .clock(r_count_80_clock),
    .reset(r_count_80_reset),
    .io_en(r_count_80_io_en),
    .io_out(r_count_80_io_out)
  );
  MyCounter r_count_81 ( // @[SWChisel.scala 171:41]
    .clock(r_count_81_clock),
    .reset(r_count_81_reset),
    .io_en(r_count_81_io_en),
    .io_out(r_count_81_io_out)
  );
  MyCounter r_count_82 ( // @[SWChisel.scala 171:41]
    .clock(r_count_82_clock),
    .reset(r_count_82_reset),
    .io_en(r_count_82_io_en),
    .io_out(r_count_82_io_out)
  );
  MyCounter r_count_83 ( // @[SWChisel.scala 171:41]
    .clock(r_count_83_clock),
    .reset(r_count_83_reset),
    .io_en(r_count_83_io_en),
    .io_out(r_count_83_io_out)
  );
  MyCounter r_count_84 ( // @[SWChisel.scala 171:41]
    .clock(r_count_84_clock),
    .reset(r_count_84_reset),
    .io_en(r_count_84_io_en),
    .io_out(r_count_84_io_out)
  );
  MyCounter r_count_85 ( // @[SWChisel.scala 171:41]
    .clock(r_count_85_clock),
    .reset(r_count_85_reset),
    .io_en(r_count_85_io_en),
    .io_out(r_count_85_io_out)
  );
  MyCounter r_count_86 ( // @[SWChisel.scala 171:41]
    .clock(r_count_86_clock),
    .reset(r_count_86_reset),
    .io_en(r_count_86_io_en),
    .io_out(r_count_86_io_out)
  );
  MyCounter r_count_87 ( // @[SWChisel.scala 171:41]
    .clock(r_count_87_clock),
    .reset(r_count_87_reset),
    .io_en(r_count_87_io_en),
    .io_out(r_count_87_io_out)
  );
  MyCounter r_count_88 ( // @[SWChisel.scala 171:41]
    .clock(r_count_88_clock),
    .reset(r_count_88_reset),
    .io_en(r_count_88_io_en),
    .io_out(r_count_88_io_out)
  );
  MyCounter r_count_89 ( // @[SWChisel.scala 171:41]
    .clock(r_count_89_clock),
    .reset(r_count_89_reset),
    .io_en(r_count_89_io_en),
    .io_out(r_count_89_io_out)
  );
  MyCounter r_count_90 ( // @[SWChisel.scala 171:41]
    .clock(r_count_90_clock),
    .reset(r_count_90_reset),
    .io_en(r_count_90_io_en),
    .io_out(r_count_90_io_out)
  );
  MyCounter r_count_91 ( // @[SWChisel.scala 171:41]
    .clock(r_count_91_clock),
    .reset(r_count_91_reset),
    .io_en(r_count_91_io_en),
    .io_out(r_count_91_io_out)
  );
  MyCounter r_count_92 ( // @[SWChisel.scala 171:41]
    .clock(r_count_92_clock),
    .reset(r_count_92_reset),
    .io_en(r_count_92_io_en),
    .io_out(r_count_92_io_out)
  );
  MyCounter r_count_93 ( // @[SWChisel.scala 171:41]
    .clock(r_count_93_clock),
    .reset(r_count_93_reset),
    .io_en(r_count_93_io_en),
    .io_out(r_count_93_io_out)
  );
  MyCounter r_count_94 ( // @[SWChisel.scala 171:41]
    .clock(r_count_94_clock),
    .reset(r_count_94_reset),
    .io_en(r_count_94_io_en),
    .io_out(r_count_94_io_out)
  );
  MyCounter r_count_95 ( // @[SWChisel.scala 171:41]
    .clock(r_count_95_clock),
    .reset(r_count_95_reset),
    .io_en(r_count_95_io_en),
    .io_out(r_count_95_io_out)
  );
  MyCounter r_count_96 ( // @[SWChisel.scala 171:41]
    .clock(r_count_96_clock),
    .reset(r_count_96_reset),
    .io_en(r_count_96_io_en),
    .io_out(r_count_96_io_out)
  );
  MyCounter r_count_97 ( // @[SWChisel.scala 171:41]
    .clock(r_count_97_clock),
    .reset(r_count_97_reset),
    .io_en(r_count_97_io_en),
    .io_out(r_count_97_io_out)
  );
  MyCounter r_count_98 ( // @[SWChisel.scala 171:41]
    .clock(r_count_98_clock),
    .reset(r_count_98_reset),
    .io_en(r_count_98_io_en),
    .io_out(r_count_98_io_out)
  );
  MyCounter r_count_99 ( // @[SWChisel.scala 171:41]
    .clock(r_count_99_clock),
    .reset(r_count_99_reset),
    .io_en(r_count_99_io_en),
    .io_out(r_count_99_io_out)
  );
  MAX max ( // @[SWChisel.scala 174:19]
    .clock(max_clock),
    .reset(max_reset),
    .io_start(max_io_start),
    .io_in(max_io_in),
    .io_done(max_io_done),
    .io_out(max_io_out)
  );
  assign io_result = max_io_out; // @[SWChisel.scala 181:13]
  assign io_done = max_io_done; // @[SWChisel.scala 182:11]
  assign array_0_io_q = io_q_0_b; // @[SWChisel.scala 220:19]
  assign array_0_io_r = 8'hc7 == r_count_0_io_out ? io_r_199_b : _GEN_498; // @[SWChisel.scala 221:{19,19}]
  assign array_0_io_e_i = E_0; // @[SWChisel.scala 196:21]
  assign array_0_io_f_i = 16'sh0; // @[SWChisel.scala 198:21]
  assign array_0_io_ve_i = V1_1; // @[SWChisel.scala 197:22]
  assign array_0_io_vf_i = V1_0; // @[SWChisel.scala 199:22]
  assign array_0_io_vv_i = V2_0; // @[SWChisel.scala 200:22]
  assign array_1_io_q = io_q_1_b; // @[SWChisel.scala 220:19]
  assign array_1_io_r = 8'hc7 == r_count_1_io_out ? io_r_199_b : _GEN_698; // @[SWChisel.scala 221:{19,19}]
  assign array_1_io_e_i = E_1; // @[SWChisel.scala 196:21]
  assign array_1_io_f_i = F_1; // @[SWChisel.scala 198:21]
  assign array_1_io_ve_i = V1_2; // @[SWChisel.scala 197:22]
  assign array_1_io_vf_i = V1_1; // @[SWChisel.scala 199:22]
  assign array_1_io_vv_i = V2_1; // @[SWChisel.scala 200:22]
  assign array_2_io_q = io_q_2_b; // @[SWChisel.scala 220:19]
  assign array_2_io_r = 8'hc7 == r_count_2_io_out ? io_r_199_b : _GEN_898; // @[SWChisel.scala 221:{19,19}]
  assign array_2_io_e_i = E_2; // @[SWChisel.scala 196:21]
  assign array_2_io_f_i = F_2; // @[SWChisel.scala 198:21]
  assign array_2_io_ve_i = V1_3; // @[SWChisel.scala 197:22]
  assign array_2_io_vf_i = V1_2; // @[SWChisel.scala 199:22]
  assign array_2_io_vv_i = V2_2; // @[SWChisel.scala 200:22]
  assign array_3_io_q = io_q_3_b; // @[SWChisel.scala 220:19]
  assign array_3_io_r = 8'hc7 == r_count_3_io_out ? io_r_199_b : _GEN_1098; // @[SWChisel.scala 221:{19,19}]
  assign array_3_io_e_i = E_3; // @[SWChisel.scala 196:21]
  assign array_3_io_f_i = F_3; // @[SWChisel.scala 198:21]
  assign array_3_io_ve_i = V1_4; // @[SWChisel.scala 197:22]
  assign array_3_io_vf_i = V1_3; // @[SWChisel.scala 199:22]
  assign array_3_io_vv_i = V2_3; // @[SWChisel.scala 200:22]
  assign array_4_io_q = io_q_4_b; // @[SWChisel.scala 220:19]
  assign array_4_io_r = 8'hc7 == r_count_4_io_out ? io_r_199_b : _GEN_1298; // @[SWChisel.scala 221:{19,19}]
  assign array_4_io_e_i = E_4; // @[SWChisel.scala 196:21]
  assign array_4_io_f_i = F_4; // @[SWChisel.scala 198:21]
  assign array_4_io_ve_i = V1_5; // @[SWChisel.scala 197:22]
  assign array_4_io_vf_i = V1_4; // @[SWChisel.scala 199:22]
  assign array_4_io_vv_i = V2_4; // @[SWChisel.scala 200:22]
  assign array_5_io_q = io_q_5_b; // @[SWChisel.scala 220:19]
  assign array_5_io_r = 8'hc7 == r_count_5_io_out ? io_r_199_b : _GEN_1498; // @[SWChisel.scala 221:{19,19}]
  assign array_5_io_e_i = E_5; // @[SWChisel.scala 196:21]
  assign array_5_io_f_i = F_5; // @[SWChisel.scala 198:21]
  assign array_5_io_ve_i = V1_6; // @[SWChisel.scala 197:22]
  assign array_5_io_vf_i = V1_5; // @[SWChisel.scala 199:22]
  assign array_5_io_vv_i = V2_5; // @[SWChisel.scala 200:22]
  assign array_6_io_q = io_q_6_b; // @[SWChisel.scala 220:19]
  assign array_6_io_r = 8'hc7 == r_count_6_io_out ? io_r_199_b : _GEN_1698; // @[SWChisel.scala 221:{19,19}]
  assign array_6_io_e_i = E_6; // @[SWChisel.scala 196:21]
  assign array_6_io_f_i = F_6; // @[SWChisel.scala 198:21]
  assign array_6_io_ve_i = V1_7; // @[SWChisel.scala 197:22]
  assign array_6_io_vf_i = V1_6; // @[SWChisel.scala 199:22]
  assign array_6_io_vv_i = V2_6; // @[SWChisel.scala 200:22]
  assign array_7_io_q = io_q_7_b; // @[SWChisel.scala 220:19]
  assign array_7_io_r = 8'hc7 == r_count_7_io_out ? io_r_199_b : _GEN_1898; // @[SWChisel.scala 221:{19,19}]
  assign array_7_io_e_i = E_7; // @[SWChisel.scala 196:21]
  assign array_7_io_f_i = F_7; // @[SWChisel.scala 198:21]
  assign array_7_io_ve_i = V1_8; // @[SWChisel.scala 197:22]
  assign array_7_io_vf_i = V1_7; // @[SWChisel.scala 199:22]
  assign array_7_io_vv_i = V2_7; // @[SWChisel.scala 200:22]
  assign array_8_io_q = io_q_8_b; // @[SWChisel.scala 220:19]
  assign array_8_io_r = 8'hc7 == r_count_8_io_out ? io_r_199_b : _GEN_2098; // @[SWChisel.scala 221:{19,19}]
  assign array_8_io_e_i = E_8; // @[SWChisel.scala 196:21]
  assign array_8_io_f_i = F_8; // @[SWChisel.scala 198:21]
  assign array_8_io_ve_i = V1_9; // @[SWChisel.scala 197:22]
  assign array_8_io_vf_i = V1_8; // @[SWChisel.scala 199:22]
  assign array_8_io_vv_i = V2_8; // @[SWChisel.scala 200:22]
  assign array_9_io_q = io_q_9_b; // @[SWChisel.scala 220:19]
  assign array_9_io_r = 8'hc7 == r_count_9_io_out ? io_r_199_b : _GEN_2298; // @[SWChisel.scala 221:{19,19}]
  assign array_9_io_e_i = E_9; // @[SWChisel.scala 196:21]
  assign array_9_io_f_i = F_9; // @[SWChisel.scala 198:21]
  assign array_9_io_ve_i = V1_10; // @[SWChisel.scala 197:22]
  assign array_9_io_vf_i = V1_9; // @[SWChisel.scala 199:22]
  assign array_9_io_vv_i = V2_9; // @[SWChisel.scala 200:22]
  assign array_10_io_q = io_q_10_b; // @[SWChisel.scala 220:19]
  assign array_10_io_r = 8'hc7 == r_count_10_io_out ? io_r_199_b : _GEN_2498; // @[SWChisel.scala 221:{19,19}]
  assign array_10_io_e_i = E_10; // @[SWChisel.scala 196:21]
  assign array_10_io_f_i = F_10; // @[SWChisel.scala 198:21]
  assign array_10_io_ve_i = V1_11; // @[SWChisel.scala 197:22]
  assign array_10_io_vf_i = V1_10; // @[SWChisel.scala 199:22]
  assign array_10_io_vv_i = V2_10; // @[SWChisel.scala 200:22]
  assign array_11_io_q = io_q_11_b; // @[SWChisel.scala 220:19]
  assign array_11_io_r = 8'hc7 == r_count_11_io_out ? io_r_199_b : _GEN_2698; // @[SWChisel.scala 221:{19,19}]
  assign array_11_io_e_i = E_11; // @[SWChisel.scala 196:21]
  assign array_11_io_f_i = F_11; // @[SWChisel.scala 198:21]
  assign array_11_io_ve_i = V1_12; // @[SWChisel.scala 197:22]
  assign array_11_io_vf_i = V1_11; // @[SWChisel.scala 199:22]
  assign array_11_io_vv_i = V2_11; // @[SWChisel.scala 200:22]
  assign array_12_io_q = io_q_12_b; // @[SWChisel.scala 220:19]
  assign array_12_io_r = 8'hc7 == r_count_12_io_out ? io_r_199_b : _GEN_2898; // @[SWChisel.scala 221:{19,19}]
  assign array_12_io_e_i = E_12; // @[SWChisel.scala 196:21]
  assign array_12_io_f_i = F_12; // @[SWChisel.scala 198:21]
  assign array_12_io_ve_i = V1_13; // @[SWChisel.scala 197:22]
  assign array_12_io_vf_i = V1_12; // @[SWChisel.scala 199:22]
  assign array_12_io_vv_i = V2_12; // @[SWChisel.scala 200:22]
  assign array_13_io_q = io_q_13_b; // @[SWChisel.scala 220:19]
  assign array_13_io_r = 8'hc7 == r_count_13_io_out ? io_r_199_b : _GEN_3098; // @[SWChisel.scala 221:{19,19}]
  assign array_13_io_e_i = E_13; // @[SWChisel.scala 196:21]
  assign array_13_io_f_i = F_13; // @[SWChisel.scala 198:21]
  assign array_13_io_ve_i = V1_14; // @[SWChisel.scala 197:22]
  assign array_13_io_vf_i = V1_13; // @[SWChisel.scala 199:22]
  assign array_13_io_vv_i = V2_13; // @[SWChisel.scala 200:22]
  assign array_14_io_q = io_q_14_b; // @[SWChisel.scala 220:19]
  assign array_14_io_r = 8'hc7 == r_count_14_io_out ? io_r_199_b : _GEN_3298; // @[SWChisel.scala 221:{19,19}]
  assign array_14_io_e_i = E_14; // @[SWChisel.scala 196:21]
  assign array_14_io_f_i = F_14; // @[SWChisel.scala 198:21]
  assign array_14_io_ve_i = V1_15; // @[SWChisel.scala 197:22]
  assign array_14_io_vf_i = V1_14; // @[SWChisel.scala 199:22]
  assign array_14_io_vv_i = V2_14; // @[SWChisel.scala 200:22]
  assign array_15_io_q = io_q_15_b; // @[SWChisel.scala 220:19]
  assign array_15_io_r = 8'hc7 == r_count_15_io_out ? io_r_199_b : _GEN_3498; // @[SWChisel.scala 221:{19,19}]
  assign array_15_io_e_i = E_15; // @[SWChisel.scala 196:21]
  assign array_15_io_f_i = F_15; // @[SWChisel.scala 198:21]
  assign array_15_io_ve_i = V1_16; // @[SWChisel.scala 197:22]
  assign array_15_io_vf_i = V1_15; // @[SWChisel.scala 199:22]
  assign array_15_io_vv_i = V2_15; // @[SWChisel.scala 200:22]
  assign array_16_io_q = io_q_16_b; // @[SWChisel.scala 220:19]
  assign array_16_io_r = 8'hc7 == r_count_16_io_out ? io_r_199_b : _GEN_3698; // @[SWChisel.scala 221:{19,19}]
  assign array_16_io_e_i = E_16; // @[SWChisel.scala 196:21]
  assign array_16_io_f_i = F_16; // @[SWChisel.scala 198:21]
  assign array_16_io_ve_i = V1_17; // @[SWChisel.scala 197:22]
  assign array_16_io_vf_i = V1_16; // @[SWChisel.scala 199:22]
  assign array_16_io_vv_i = V2_16; // @[SWChisel.scala 200:22]
  assign array_17_io_q = io_q_17_b; // @[SWChisel.scala 220:19]
  assign array_17_io_r = 8'hc7 == r_count_17_io_out ? io_r_199_b : _GEN_3898; // @[SWChisel.scala 221:{19,19}]
  assign array_17_io_e_i = E_17; // @[SWChisel.scala 196:21]
  assign array_17_io_f_i = F_17; // @[SWChisel.scala 198:21]
  assign array_17_io_ve_i = V1_18; // @[SWChisel.scala 197:22]
  assign array_17_io_vf_i = V1_17; // @[SWChisel.scala 199:22]
  assign array_17_io_vv_i = V2_17; // @[SWChisel.scala 200:22]
  assign array_18_io_q = io_q_18_b; // @[SWChisel.scala 220:19]
  assign array_18_io_r = 8'hc7 == r_count_18_io_out ? io_r_199_b : _GEN_4098; // @[SWChisel.scala 221:{19,19}]
  assign array_18_io_e_i = E_18; // @[SWChisel.scala 196:21]
  assign array_18_io_f_i = F_18; // @[SWChisel.scala 198:21]
  assign array_18_io_ve_i = V1_19; // @[SWChisel.scala 197:22]
  assign array_18_io_vf_i = V1_18; // @[SWChisel.scala 199:22]
  assign array_18_io_vv_i = V2_18; // @[SWChisel.scala 200:22]
  assign array_19_io_q = io_q_19_b; // @[SWChisel.scala 220:19]
  assign array_19_io_r = 8'hc7 == r_count_19_io_out ? io_r_199_b : _GEN_4298; // @[SWChisel.scala 221:{19,19}]
  assign array_19_io_e_i = E_19; // @[SWChisel.scala 196:21]
  assign array_19_io_f_i = F_19; // @[SWChisel.scala 198:21]
  assign array_19_io_ve_i = V1_20; // @[SWChisel.scala 197:22]
  assign array_19_io_vf_i = V1_19; // @[SWChisel.scala 199:22]
  assign array_19_io_vv_i = V2_19; // @[SWChisel.scala 200:22]
  assign array_20_io_q = io_q_20_b; // @[SWChisel.scala 220:19]
  assign array_20_io_r = 8'hc7 == r_count_20_io_out ? io_r_199_b : _GEN_4498; // @[SWChisel.scala 221:{19,19}]
  assign array_20_io_e_i = E_20; // @[SWChisel.scala 196:21]
  assign array_20_io_f_i = F_20; // @[SWChisel.scala 198:21]
  assign array_20_io_ve_i = V1_21; // @[SWChisel.scala 197:22]
  assign array_20_io_vf_i = V1_20; // @[SWChisel.scala 199:22]
  assign array_20_io_vv_i = V2_20; // @[SWChisel.scala 200:22]
  assign array_21_io_q = io_q_21_b; // @[SWChisel.scala 220:19]
  assign array_21_io_r = 8'hc7 == r_count_21_io_out ? io_r_199_b : _GEN_4698; // @[SWChisel.scala 221:{19,19}]
  assign array_21_io_e_i = E_21; // @[SWChisel.scala 196:21]
  assign array_21_io_f_i = F_21; // @[SWChisel.scala 198:21]
  assign array_21_io_ve_i = V1_22; // @[SWChisel.scala 197:22]
  assign array_21_io_vf_i = V1_21; // @[SWChisel.scala 199:22]
  assign array_21_io_vv_i = V2_21; // @[SWChisel.scala 200:22]
  assign array_22_io_q = io_q_22_b; // @[SWChisel.scala 220:19]
  assign array_22_io_r = 8'hc7 == r_count_22_io_out ? io_r_199_b : _GEN_4898; // @[SWChisel.scala 221:{19,19}]
  assign array_22_io_e_i = E_22; // @[SWChisel.scala 196:21]
  assign array_22_io_f_i = F_22; // @[SWChisel.scala 198:21]
  assign array_22_io_ve_i = V1_23; // @[SWChisel.scala 197:22]
  assign array_22_io_vf_i = V1_22; // @[SWChisel.scala 199:22]
  assign array_22_io_vv_i = V2_22; // @[SWChisel.scala 200:22]
  assign array_23_io_q = io_q_23_b; // @[SWChisel.scala 220:19]
  assign array_23_io_r = 8'hc7 == r_count_23_io_out ? io_r_199_b : _GEN_5098; // @[SWChisel.scala 221:{19,19}]
  assign array_23_io_e_i = E_23; // @[SWChisel.scala 196:21]
  assign array_23_io_f_i = F_23; // @[SWChisel.scala 198:21]
  assign array_23_io_ve_i = V1_24; // @[SWChisel.scala 197:22]
  assign array_23_io_vf_i = V1_23; // @[SWChisel.scala 199:22]
  assign array_23_io_vv_i = V2_23; // @[SWChisel.scala 200:22]
  assign array_24_io_q = io_q_24_b; // @[SWChisel.scala 220:19]
  assign array_24_io_r = 8'hc7 == r_count_24_io_out ? io_r_199_b : _GEN_5298; // @[SWChisel.scala 221:{19,19}]
  assign array_24_io_e_i = E_24; // @[SWChisel.scala 196:21]
  assign array_24_io_f_i = F_24; // @[SWChisel.scala 198:21]
  assign array_24_io_ve_i = V1_25; // @[SWChisel.scala 197:22]
  assign array_24_io_vf_i = V1_24; // @[SWChisel.scala 199:22]
  assign array_24_io_vv_i = V2_24; // @[SWChisel.scala 200:22]
  assign array_25_io_q = io_q_25_b; // @[SWChisel.scala 220:19]
  assign array_25_io_r = 8'hc7 == r_count_25_io_out ? io_r_199_b : _GEN_5498; // @[SWChisel.scala 221:{19,19}]
  assign array_25_io_e_i = E_25; // @[SWChisel.scala 196:21]
  assign array_25_io_f_i = F_25; // @[SWChisel.scala 198:21]
  assign array_25_io_ve_i = V1_26; // @[SWChisel.scala 197:22]
  assign array_25_io_vf_i = V1_25; // @[SWChisel.scala 199:22]
  assign array_25_io_vv_i = V2_25; // @[SWChisel.scala 200:22]
  assign array_26_io_q = io_q_26_b; // @[SWChisel.scala 220:19]
  assign array_26_io_r = 8'hc7 == r_count_26_io_out ? io_r_199_b : _GEN_5698; // @[SWChisel.scala 221:{19,19}]
  assign array_26_io_e_i = E_26; // @[SWChisel.scala 196:21]
  assign array_26_io_f_i = F_26; // @[SWChisel.scala 198:21]
  assign array_26_io_ve_i = V1_27; // @[SWChisel.scala 197:22]
  assign array_26_io_vf_i = V1_26; // @[SWChisel.scala 199:22]
  assign array_26_io_vv_i = V2_26; // @[SWChisel.scala 200:22]
  assign array_27_io_q = io_q_27_b; // @[SWChisel.scala 220:19]
  assign array_27_io_r = 8'hc7 == r_count_27_io_out ? io_r_199_b : _GEN_5898; // @[SWChisel.scala 221:{19,19}]
  assign array_27_io_e_i = E_27; // @[SWChisel.scala 196:21]
  assign array_27_io_f_i = F_27; // @[SWChisel.scala 198:21]
  assign array_27_io_ve_i = V1_28; // @[SWChisel.scala 197:22]
  assign array_27_io_vf_i = V1_27; // @[SWChisel.scala 199:22]
  assign array_27_io_vv_i = V2_27; // @[SWChisel.scala 200:22]
  assign array_28_io_q = io_q_28_b; // @[SWChisel.scala 220:19]
  assign array_28_io_r = 8'hc7 == r_count_28_io_out ? io_r_199_b : _GEN_6098; // @[SWChisel.scala 221:{19,19}]
  assign array_28_io_e_i = E_28; // @[SWChisel.scala 196:21]
  assign array_28_io_f_i = F_28; // @[SWChisel.scala 198:21]
  assign array_28_io_ve_i = V1_29; // @[SWChisel.scala 197:22]
  assign array_28_io_vf_i = V1_28; // @[SWChisel.scala 199:22]
  assign array_28_io_vv_i = V2_28; // @[SWChisel.scala 200:22]
  assign array_29_io_q = io_q_29_b; // @[SWChisel.scala 220:19]
  assign array_29_io_r = 8'hc7 == r_count_29_io_out ? io_r_199_b : _GEN_6298; // @[SWChisel.scala 221:{19,19}]
  assign array_29_io_e_i = E_29; // @[SWChisel.scala 196:21]
  assign array_29_io_f_i = F_29; // @[SWChisel.scala 198:21]
  assign array_29_io_ve_i = V1_30; // @[SWChisel.scala 197:22]
  assign array_29_io_vf_i = V1_29; // @[SWChisel.scala 199:22]
  assign array_29_io_vv_i = V2_29; // @[SWChisel.scala 200:22]
  assign array_30_io_q = io_q_30_b; // @[SWChisel.scala 220:19]
  assign array_30_io_r = 8'hc7 == r_count_30_io_out ? io_r_199_b : _GEN_6498; // @[SWChisel.scala 221:{19,19}]
  assign array_30_io_e_i = E_30; // @[SWChisel.scala 196:21]
  assign array_30_io_f_i = F_30; // @[SWChisel.scala 198:21]
  assign array_30_io_ve_i = V1_31; // @[SWChisel.scala 197:22]
  assign array_30_io_vf_i = V1_30; // @[SWChisel.scala 199:22]
  assign array_30_io_vv_i = V2_30; // @[SWChisel.scala 200:22]
  assign array_31_io_q = io_q_31_b; // @[SWChisel.scala 220:19]
  assign array_31_io_r = 8'hc7 == r_count_31_io_out ? io_r_199_b : _GEN_6698; // @[SWChisel.scala 221:{19,19}]
  assign array_31_io_e_i = E_31; // @[SWChisel.scala 196:21]
  assign array_31_io_f_i = F_31; // @[SWChisel.scala 198:21]
  assign array_31_io_ve_i = V1_32; // @[SWChisel.scala 197:22]
  assign array_31_io_vf_i = V1_31; // @[SWChisel.scala 199:22]
  assign array_31_io_vv_i = V2_31; // @[SWChisel.scala 200:22]
  assign array_32_io_q = io_q_32_b; // @[SWChisel.scala 220:19]
  assign array_32_io_r = 8'hc7 == r_count_32_io_out ? io_r_199_b : _GEN_6898; // @[SWChisel.scala 221:{19,19}]
  assign array_32_io_e_i = E_32; // @[SWChisel.scala 196:21]
  assign array_32_io_f_i = F_32; // @[SWChisel.scala 198:21]
  assign array_32_io_ve_i = V1_33; // @[SWChisel.scala 197:22]
  assign array_32_io_vf_i = V1_32; // @[SWChisel.scala 199:22]
  assign array_32_io_vv_i = V2_32; // @[SWChisel.scala 200:22]
  assign array_33_io_q = io_q_33_b; // @[SWChisel.scala 220:19]
  assign array_33_io_r = 8'hc7 == r_count_33_io_out ? io_r_199_b : _GEN_7098; // @[SWChisel.scala 221:{19,19}]
  assign array_33_io_e_i = E_33; // @[SWChisel.scala 196:21]
  assign array_33_io_f_i = F_33; // @[SWChisel.scala 198:21]
  assign array_33_io_ve_i = V1_34; // @[SWChisel.scala 197:22]
  assign array_33_io_vf_i = V1_33; // @[SWChisel.scala 199:22]
  assign array_33_io_vv_i = V2_33; // @[SWChisel.scala 200:22]
  assign array_34_io_q = io_q_34_b; // @[SWChisel.scala 220:19]
  assign array_34_io_r = 8'hc7 == r_count_34_io_out ? io_r_199_b : _GEN_7298; // @[SWChisel.scala 221:{19,19}]
  assign array_34_io_e_i = E_34; // @[SWChisel.scala 196:21]
  assign array_34_io_f_i = F_34; // @[SWChisel.scala 198:21]
  assign array_34_io_ve_i = V1_35; // @[SWChisel.scala 197:22]
  assign array_34_io_vf_i = V1_34; // @[SWChisel.scala 199:22]
  assign array_34_io_vv_i = V2_34; // @[SWChisel.scala 200:22]
  assign array_35_io_q = io_q_35_b; // @[SWChisel.scala 220:19]
  assign array_35_io_r = 8'hc7 == r_count_35_io_out ? io_r_199_b : _GEN_7498; // @[SWChisel.scala 221:{19,19}]
  assign array_35_io_e_i = E_35; // @[SWChisel.scala 196:21]
  assign array_35_io_f_i = F_35; // @[SWChisel.scala 198:21]
  assign array_35_io_ve_i = V1_36; // @[SWChisel.scala 197:22]
  assign array_35_io_vf_i = V1_35; // @[SWChisel.scala 199:22]
  assign array_35_io_vv_i = V2_35; // @[SWChisel.scala 200:22]
  assign array_36_io_q = io_q_36_b; // @[SWChisel.scala 220:19]
  assign array_36_io_r = 8'hc7 == r_count_36_io_out ? io_r_199_b : _GEN_7698; // @[SWChisel.scala 221:{19,19}]
  assign array_36_io_e_i = E_36; // @[SWChisel.scala 196:21]
  assign array_36_io_f_i = F_36; // @[SWChisel.scala 198:21]
  assign array_36_io_ve_i = V1_37; // @[SWChisel.scala 197:22]
  assign array_36_io_vf_i = V1_36; // @[SWChisel.scala 199:22]
  assign array_36_io_vv_i = V2_36; // @[SWChisel.scala 200:22]
  assign array_37_io_q = io_q_37_b; // @[SWChisel.scala 220:19]
  assign array_37_io_r = 8'hc7 == r_count_37_io_out ? io_r_199_b : _GEN_7898; // @[SWChisel.scala 221:{19,19}]
  assign array_37_io_e_i = E_37; // @[SWChisel.scala 196:21]
  assign array_37_io_f_i = F_37; // @[SWChisel.scala 198:21]
  assign array_37_io_ve_i = V1_38; // @[SWChisel.scala 197:22]
  assign array_37_io_vf_i = V1_37; // @[SWChisel.scala 199:22]
  assign array_37_io_vv_i = V2_37; // @[SWChisel.scala 200:22]
  assign array_38_io_q = io_q_38_b; // @[SWChisel.scala 220:19]
  assign array_38_io_r = 8'hc7 == r_count_38_io_out ? io_r_199_b : _GEN_8098; // @[SWChisel.scala 221:{19,19}]
  assign array_38_io_e_i = E_38; // @[SWChisel.scala 196:21]
  assign array_38_io_f_i = F_38; // @[SWChisel.scala 198:21]
  assign array_38_io_ve_i = V1_39; // @[SWChisel.scala 197:22]
  assign array_38_io_vf_i = V1_38; // @[SWChisel.scala 199:22]
  assign array_38_io_vv_i = V2_38; // @[SWChisel.scala 200:22]
  assign array_39_io_q = io_q_39_b; // @[SWChisel.scala 220:19]
  assign array_39_io_r = 8'hc7 == r_count_39_io_out ? io_r_199_b : _GEN_8298; // @[SWChisel.scala 221:{19,19}]
  assign array_39_io_e_i = E_39; // @[SWChisel.scala 196:21]
  assign array_39_io_f_i = F_39; // @[SWChisel.scala 198:21]
  assign array_39_io_ve_i = V1_40; // @[SWChisel.scala 197:22]
  assign array_39_io_vf_i = V1_39; // @[SWChisel.scala 199:22]
  assign array_39_io_vv_i = V2_39; // @[SWChisel.scala 200:22]
  assign array_40_io_q = io_q_40_b; // @[SWChisel.scala 220:19]
  assign array_40_io_r = 8'hc7 == r_count_40_io_out ? io_r_199_b : _GEN_8498; // @[SWChisel.scala 221:{19,19}]
  assign array_40_io_e_i = E_40; // @[SWChisel.scala 196:21]
  assign array_40_io_f_i = F_40; // @[SWChisel.scala 198:21]
  assign array_40_io_ve_i = V1_41; // @[SWChisel.scala 197:22]
  assign array_40_io_vf_i = V1_40; // @[SWChisel.scala 199:22]
  assign array_40_io_vv_i = V2_40; // @[SWChisel.scala 200:22]
  assign array_41_io_q = io_q_41_b; // @[SWChisel.scala 220:19]
  assign array_41_io_r = 8'hc7 == r_count_41_io_out ? io_r_199_b : _GEN_8698; // @[SWChisel.scala 221:{19,19}]
  assign array_41_io_e_i = E_41; // @[SWChisel.scala 196:21]
  assign array_41_io_f_i = F_41; // @[SWChisel.scala 198:21]
  assign array_41_io_ve_i = V1_42; // @[SWChisel.scala 197:22]
  assign array_41_io_vf_i = V1_41; // @[SWChisel.scala 199:22]
  assign array_41_io_vv_i = V2_41; // @[SWChisel.scala 200:22]
  assign array_42_io_q = io_q_42_b; // @[SWChisel.scala 220:19]
  assign array_42_io_r = 8'hc7 == r_count_42_io_out ? io_r_199_b : _GEN_8898; // @[SWChisel.scala 221:{19,19}]
  assign array_42_io_e_i = E_42; // @[SWChisel.scala 196:21]
  assign array_42_io_f_i = F_42; // @[SWChisel.scala 198:21]
  assign array_42_io_ve_i = V1_43; // @[SWChisel.scala 197:22]
  assign array_42_io_vf_i = V1_42; // @[SWChisel.scala 199:22]
  assign array_42_io_vv_i = V2_42; // @[SWChisel.scala 200:22]
  assign array_43_io_q = io_q_43_b; // @[SWChisel.scala 220:19]
  assign array_43_io_r = 8'hc7 == r_count_43_io_out ? io_r_199_b : _GEN_9098; // @[SWChisel.scala 221:{19,19}]
  assign array_43_io_e_i = E_43; // @[SWChisel.scala 196:21]
  assign array_43_io_f_i = F_43; // @[SWChisel.scala 198:21]
  assign array_43_io_ve_i = V1_44; // @[SWChisel.scala 197:22]
  assign array_43_io_vf_i = V1_43; // @[SWChisel.scala 199:22]
  assign array_43_io_vv_i = V2_43; // @[SWChisel.scala 200:22]
  assign array_44_io_q = io_q_44_b; // @[SWChisel.scala 220:19]
  assign array_44_io_r = 8'hc7 == r_count_44_io_out ? io_r_199_b : _GEN_9298; // @[SWChisel.scala 221:{19,19}]
  assign array_44_io_e_i = E_44; // @[SWChisel.scala 196:21]
  assign array_44_io_f_i = F_44; // @[SWChisel.scala 198:21]
  assign array_44_io_ve_i = V1_45; // @[SWChisel.scala 197:22]
  assign array_44_io_vf_i = V1_44; // @[SWChisel.scala 199:22]
  assign array_44_io_vv_i = V2_44; // @[SWChisel.scala 200:22]
  assign array_45_io_q = io_q_45_b; // @[SWChisel.scala 220:19]
  assign array_45_io_r = 8'hc7 == r_count_45_io_out ? io_r_199_b : _GEN_9498; // @[SWChisel.scala 221:{19,19}]
  assign array_45_io_e_i = E_45; // @[SWChisel.scala 196:21]
  assign array_45_io_f_i = F_45; // @[SWChisel.scala 198:21]
  assign array_45_io_ve_i = V1_46; // @[SWChisel.scala 197:22]
  assign array_45_io_vf_i = V1_45; // @[SWChisel.scala 199:22]
  assign array_45_io_vv_i = V2_45; // @[SWChisel.scala 200:22]
  assign array_46_io_q = io_q_46_b; // @[SWChisel.scala 220:19]
  assign array_46_io_r = 8'hc7 == r_count_46_io_out ? io_r_199_b : _GEN_9698; // @[SWChisel.scala 221:{19,19}]
  assign array_46_io_e_i = E_46; // @[SWChisel.scala 196:21]
  assign array_46_io_f_i = F_46; // @[SWChisel.scala 198:21]
  assign array_46_io_ve_i = V1_47; // @[SWChisel.scala 197:22]
  assign array_46_io_vf_i = V1_46; // @[SWChisel.scala 199:22]
  assign array_46_io_vv_i = V2_46; // @[SWChisel.scala 200:22]
  assign array_47_io_q = io_q_47_b; // @[SWChisel.scala 220:19]
  assign array_47_io_r = 8'hc7 == r_count_47_io_out ? io_r_199_b : _GEN_9898; // @[SWChisel.scala 221:{19,19}]
  assign array_47_io_e_i = E_47; // @[SWChisel.scala 196:21]
  assign array_47_io_f_i = F_47; // @[SWChisel.scala 198:21]
  assign array_47_io_ve_i = V1_48; // @[SWChisel.scala 197:22]
  assign array_47_io_vf_i = V1_47; // @[SWChisel.scala 199:22]
  assign array_47_io_vv_i = V2_47; // @[SWChisel.scala 200:22]
  assign array_48_io_q = io_q_48_b; // @[SWChisel.scala 220:19]
  assign array_48_io_r = 8'hc7 == r_count_48_io_out ? io_r_199_b : _GEN_10098; // @[SWChisel.scala 221:{19,19}]
  assign array_48_io_e_i = E_48; // @[SWChisel.scala 196:21]
  assign array_48_io_f_i = F_48; // @[SWChisel.scala 198:21]
  assign array_48_io_ve_i = V1_49; // @[SWChisel.scala 197:22]
  assign array_48_io_vf_i = V1_48; // @[SWChisel.scala 199:22]
  assign array_48_io_vv_i = V2_48; // @[SWChisel.scala 200:22]
  assign array_49_io_q = io_q_49_b; // @[SWChisel.scala 220:19]
  assign array_49_io_r = 8'hc7 == r_count_49_io_out ? io_r_199_b : _GEN_10298; // @[SWChisel.scala 221:{19,19}]
  assign array_49_io_e_i = E_49; // @[SWChisel.scala 196:21]
  assign array_49_io_f_i = F_49; // @[SWChisel.scala 198:21]
  assign array_49_io_ve_i = V1_50; // @[SWChisel.scala 197:22]
  assign array_49_io_vf_i = V1_49; // @[SWChisel.scala 199:22]
  assign array_49_io_vv_i = V2_49; // @[SWChisel.scala 200:22]
  assign array_50_io_q = io_q_50_b; // @[SWChisel.scala 220:19]
  assign array_50_io_r = 8'hc7 == r_count_50_io_out ? io_r_199_b : _GEN_10498; // @[SWChisel.scala 221:{19,19}]
  assign array_50_io_e_i = E_50; // @[SWChisel.scala 196:21]
  assign array_50_io_f_i = F_50; // @[SWChisel.scala 198:21]
  assign array_50_io_ve_i = V1_51; // @[SWChisel.scala 197:22]
  assign array_50_io_vf_i = V1_50; // @[SWChisel.scala 199:22]
  assign array_50_io_vv_i = V2_50; // @[SWChisel.scala 200:22]
  assign array_51_io_q = io_q_51_b; // @[SWChisel.scala 220:19]
  assign array_51_io_r = 8'hc7 == r_count_51_io_out ? io_r_199_b : _GEN_10698; // @[SWChisel.scala 221:{19,19}]
  assign array_51_io_e_i = E_51; // @[SWChisel.scala 196:21]
  assign array_51_io_f_i = F_51; // @[SWChisel.scala 198:21]
  assign array_51_io_ve_i = V1_52; // @[SWChisel.scala 197:22]
  assign array_51_io_vf_i = V1_51; // @[SWChisel.scala 199:22]
  assign array_51_io_vv_i = V2_51; // @[SWChisel.scala 200:22]
  assign array_52_io_q = io_q_52_b; // @[SWChisel.scala 220:19]
  assign array_52_io_r = 8'hc7 == r_count_52_io_out ? io_r_199_b : _GEN_10898; // @[SWChisel.scala 221:{19,19}]
  assign array_52_io_e_i = E_52; // @[SWChisel.scala 196:21]
  assign array_52_io_f_i = F_52; // @[SWChisel.scala 198:21]
  assign array_52_io_ve_i = V1_53; // @[SWChisel.scala 197:22]
  assign array_52_io_vf_i = V1_52; // @[SWChisel.scala 199:22]
  assign array_52_io_vv_i = V2_52; // @[SWChisel.scala 200:22]
  assign array_53_io_q = io_q_53_b; // @[SWChisel.scala 220:19]
  assign array_53_io_r = 8'hc7 == r_count_53_io_out ? io_r_199_b : _GEN_11098; // @[SWChisel.scala 221:{19,19}]
  assign array_53_io_e_i = E_53; // @[SWChisel.scala 196:21]
  assign array_53_io_f_i = F_53; // @[SWChisel.scala 198:21]
  assign array_53_io_ve_i = V1_54; // @[SWChisel.scala 197:22]
  assign array_53_io_vf_i = V1_53; // @[SWChisel.scala 199:22]
  assign array_53_io_vv_i = V2_53; // @[SWChisel.scala 200:22]
  assign array_54_io_q = io_q_54_b; // @[SWChisel.scala 220:19]
  assign array_54_io_r = 8'hc7 == r_count_54_io_out ? io_r_199_b : _GEN_11298; // @[SWChisel.scala 221:{19,19}]
  assign array_54_io_e_i = E_54; // @[SWChisel.scala 196:21]
  assign array_54_io_f_i = F_54; // @[SWChisel.scala 198:21]
  assign array_54_io_ve_i = V1_55; // @[SWChisel.scala 197:22]
  assign array_54_io_vf_i = V1_54; // @[SWChisel.scala 199:22]
  assign array_54_io_vv_i = V2_54; // @[SWChisel.scala 200:22]
  assign array_55_io_q = io_q_55_b; // @[SWChisel.scala 220:19]
  assign array_55_io_r = 8'hc7 == r_count_55_io_out ? io_r_199_b : _GEN_11498; // @[SWChisel.scala 221:{19,19}]
  assign array_55_io_e_i = E_55; // @[SWChisel.scala 196:21]
  assign array_55_io_f_i = F_55; // @[SWChisel.scala 198:21]
  assign array_55_io_ve_i = V1_56; // @[SWChisel.scala 197:22]
  assign array_55_io_vf_i = V1_55; // @[SWChisel.scala 199:22]
  assign array_55_io_vv_i = V2_55; // @[SWChisel.scala 200:22]
  assign array_56_io_q = io_q_56_b; // @[SWChisel.scala 220:19]
  assign array_56_io_r = 8'hc7 == r_count_56_io_out ? io_r_199_b : _GEN_11698; // @[SWChisel.scala 221:{19,19}]
  assign array_56_io_e_i = E_56; // @[SWChisel.scala 196:21]
  assign array_56_io_f_i = F_56; // @[SWChisel.scala 198:21]
  assign array_56_io_ve_i = V1_57; // @[SWChisel.scala 197:22]
  assign array_56_io_vf_i = V1_56; // @[SWChisel.scala 199:22]
  assign array_56_io_vv_i = V2_56; // @[SWChisel.scala 200:22]
  assign array_57_io_q = io_q_57_b; // @[SWChisel.scala 220:19]
  assign array_57_io_r = 8'hc7 == r_count_57_io_out ? io_r_199_b : _GEN_11898; // @[SWChisel.scala 221:{19,19}]
  assign array_57_io_e_i = E_57; // @[SWChisel.scala 196:21]
  assign array_57_io_f_i = F_57; // @[SWChisel.scala 198:21]
  assign array_57_io_ve_i = V1_58; // @[SWChisel.scala 197:22]
  assign array_57_io_vf_i = V1_57; // @[SWChisel.scala 199:22]
  assign array_57_io_vv_i = V2_57; // @[SWChisel.scala 200:22]
  assign array_58_io_q = io_q_58_b; // @[SWChisel.scala 220:19]
  assign array_58_io_r = 8'hc7 == r_count_58_io_out ? io_r_199_b : _GEN_12098; // @[SWChisel.scala 221:{19,19}]
  assign array_58_io_e_i = E_58; // @[SWChisel.scala 196:21]
  assign array_58_io_f_i = F_58; // @[SWChisel.scala 198:21]
  assign array_58_io_ve_i = V1_59; // @[SWChisel.scala 197:22]
  assign array_58_io_vf_i = V1_58; // @[SWChisel.scala 199:22]
  assign array_58_io_vv_i = V2_58; // @[SWChisel.scala 200:22]
  assign array_59_io_q = io_q_59_b; // @[SWChisel.scala 220:19]
  assign array_59_io_r = 8'hc7 == r_count_59_io_out ? io_r_199_b : _GEN_12298; // @[SWChisel.scala 221:{19,19}]
  assign array_59_io_e_i = E_59; // @[SWChisel.scala 196:21]
  assign array_59_io_f_i = F_59; // @[SWChisel.scala 198:21]
  assign array_59_io_ve_i = V1_60; // @[SWChisel.scala 197:22]
  assign array_59_io_vf_i = V1_59; // @[SWChisel.scala 199:22]
  assign array_59_io_vv_i = V2_59; // @[SWChisel.scala 200:22]
  assign array_60_io_q = io_q_60_b; // @[SWChisel.scala 220:19]
  assign array_60_io_r = 8'hc7 == r_count_60_io_out ? io_r_199_b : _GEN_12498; // @[SWChisel.scala 221:{19,19}]
  assign array_60_io_e_i = E_60; // @[SWChisel.scala 196:21]
  assign array_60_io_f_i = F_60; // @[SWChisel.scala 198:21]
  assign array_60_io_ve_i = V1_61; // @[SWChisel.scala 197:22]
  assign array_60_io_vf_i = V1_60; // @[SWChisel.scala 199:22]
  assign array_60_io_vv_i = V2_60; // @[SWChisel.scala 200:22]
  assign array_61_io_q = io_q_61_b; // @[SWChisel.scala 220:19]
  assign array_61_io_r = 8'hc7 == r_count_61_io_out ? io_r_199_b : _GEN_12698; // @[SWChisel.scala 221:{19,19}]
  assign array_61_io_e_i = E_61; // @[SWChisel.scala 196:21]
  assign array_61_io_f_i = F_61; // @[SWChisel.scala 198:21]
  assign array_61_io_ve_i = V1_62; // @[SWChisel.scala 197:22]
  assign array_61_io_vf_i = V1_61; // @[SWChisel.scala 199:22]
  assign array_61_io_vv_i = V2_61; // @[SWChisel.scala 200:22]
  assign array_62_io_q = io_q_62_b; // @[SWChisel.scala 220:19]
  assign array_62_io_r = 8'hc7 == r_count_62_io_out ? io_r_199_b : _GEN_12898; // @[SWChisel.scala 221:{19,19}]
  assign array_62_io_e_i = E_62; // @[SWChisel.scala 196:21]
  assign array_62_io_f_i = F_62; // @[SWChisel.scala 198:21]
  assign array_62_io_ve_i = V1_63; // @[SWChisel.scala 197:22]
  assign array_62_io_vf_i = V1_62; // @[SWChisel.scala 199:22]
  assign array_62_io_vv_i = V2_62; // @[SWChisel.scala 200:22]
  assign array_63_io_q = io_q_63_b; // @[SWChisel.scala 220:19]
  assign array_63_io_r = 8'hc7 == r_count_63_io_out ? io_r_199_b : _GEN_13098; // @[SWChisel.scala 221:{19,19}]
  assign array_63_io_e_i = E_63; // @[SWChisel.scala 196:21]
  assign array_63_io_f_i = F_63; // @[SWChisel.scala 198:21]
  assign array_63_io_ve_i = V1_64; // @[SWChisel.scala 197:22]
  assign array_63_io_vf_i = V1_63; // @[SWChisel.scala 199:22]
  assign array_63_io_vv_i = V2_63; // @[SWChisel.scala 200:22]
  assign array_64_io_q = io_q_64_b; // @[SWChisel.scala 220:19]
  assign array_64_io_r = 8'hc7 == r_count_64_io_out ? io_r_199_b : _GEN_13298; // @[SWChisel.scala 221:{19,19}]
  assign array_64_io_e_i = E_64; // @[SWChisel.scala 196:21]
  assign array_64_io_f_i = F_64; // @[SWChisel.scala 198:21]
  assign array_64_io_ve_i = V1_65; // @[SWChisel.scala 197:22]
  assign array_64_io_vf_i = V1_64; // @[SWChisel.scala 199:22]
  assign array_64_io_vv_i = V2_64; // @[SWChisel.scala 200:22]
  assign array_65_io_q = io_q_65_b; // @[SWChisel.scala 220:19]
  assign array_65_io_r = 8'hc7 == r_count_65_io_out ? io_r_199_b : _GEN_13498; // @[SWChisel.scala 221:{19,19}]
  assign array_65_io_e_i = E_65; // @[SWChisel.scala 196:21]
  assign array_65_io_f_i = F_65; // @[SWChisel.scala 198:21]
  assign array_65_io_ve_i = V1_66; // @[SWChisel.scala 197:22]
  assign array_65_io_vf_i = V1_65; // @[SWChisel.scala 199:22]
  assign array_65_io_vv_i = V2_65; // @[SWChisel.scala 200:22]
  assign array_66_io_q = io_q_66_b; // @[SWChisel.scala 220:19]
  assign array_66_io_r = 8'hc7 == r_count_66_io_out ? io_r_199_b : _GEN_13698; // @[SWChisel.scala 221:{19,19}]
  assign array_66_io_e_i = E_66; // @[SWChisel.scala 196:21]
  assign array_66_io_f_i = F_66; // @[SWChisel.scala 198:21]
  assign array_66_io_ve_i = V1_67; // @[SWChisel.scala 197:22]
  assign array_66_io_vf_i = V1_66; // @[SWChisel.scala 199:22]
  assign array_66_io_vv_i = V2_66; // @[SWChisel.scala 200:22]
  assign array_67_io_q = io_q_67_b; // @[SWChisel.scala 220:19]
  assign array_67_io_r = 8'hc7 == r_count_67_io_out ? io_r_199_b : _GEN_13898; // @[SWChisel.scala 221:{19,19}]
  assign array_67_io_e_i = E_67; // @[SWChisel.scala 196:21]
  assign array_67_io_f_i = F_67; // @[SWChisel.scala 198:21]
  assign array_67_io_ve_i = V1_68; // @[SWChisel.scala 197:22]
  assign array_67_io_vf_i = V1_67; // @[SWChisel.scala 199:22]
  assign array_67_io_vv_i = V2_67; // @[SWChisel.scala 200:22]
  assign array_68_io_q = io_q_68_b; // @[SWChisel.scala 220:19]
  assign array_68_io_r = 8'hc7 == r_count_68_io_out ? io_r_199_b : _GEN_14098; // @[SWChisel.scala 221:{19,19}]
  assign array_68_io_e_i = E_68; // @[SWChisel.scala 196:21]
  assign array_68_io_f_i = F_68; // @[SWChisel.scala 198:21]
  assign array_68_io_ve_i = V1_69; // @[SWChisel.scala 197:22]
  assign array_68_io_vf_i = V1_68; // @[SWChisel.scala 199:22]
  assign array_68_io_vv_i = V2_68; // @[SWChisel.scala 200:22]
  assign array_69_io_q = io_q_69_b; // @[SWChisel.scala 220:19]
  assign array_69_io_r = 8'hc7 == r_count_69_io_out ? io_r_199_b : _GEN_14298; // @[SWChisel.scala 221:{19,19}]
  assign array_69_io_e_i = E_69; // @[SWChisel.scala 196:21]
  assign array_69_io_f_i = F_69; // @[SWChisel.scala 198:21]
  assign array_69_io_ve_i = V1_70; // @[SWChisel.scala 197:22]
  assign array_69_io_vf_i = V1_69; // @[SWChisel.scala 199:22]
  assign array_69_io_vv_i = V2_69; // @[SWChisel.scala 200:22]
  assign array_70_io_q = io_q_70_b; // @[SWChisel.scala 220:19]
  assign array_70_io_r = 8'hc7 == r_count_70_io_out ? io_r_199_b : _GEN_14498; // @[SWChisel.scala 221:{19,19}]
  assign array_70_io_e_i = E_70; // @[SWChisel.scala 196:21]
  assign array_70_io_f_i = F_70; // @[SWChisel.scala 198:21]
  assign array_70_io_ve_i = V1_71; // @[SWChisel.scala 197:22]
  assign array_70_io_vf_i = V1_70; // @[SWChisel.scala 199:22]
  assign array_70_io_vv_i = V2_70; // @[SWChisel.scala 200:22]
  assign array_71_io_q = io_q_71_b; // @[SWChisel.scala 220:19]
  assign array_71_io_r = 8'hc7 == r_count_71_io_out ? io_r_199_b : _GEN_14698; // @[SWChisel.scala 221:{19,19}]
  assign array_71_io_e_i = E_71; // @[SWChisel.scala 196:21]
  assign array_71_io_f_i = F_71; // @[SWChisel.scala 198:21]
  assign array_71_io_ve_i = V1_72; // @[SWChisel.scala 197:22]
  assign array_71_io_vf_i = V1_71; // @[SWChisel.scala 199:22]
  assign array_71_io_vv_i = V2_71; // @[SWChisel.scala 200:22]
  assign array_72_io_q = io_q_72_b; // @[SWChisel.scala 220:19]
  assign array_72_io_r = 8'hc7 == r_count_72_io_out ? io_r_199_b : _GEN_14898; // @[SWChisel.scala 221:{19,19}]
  assign array_72_io_e_i = E_72; // @[SWChisel.scala 196:21]
  assign array_72_io_f_i = F_72; // @[SWChisel.scala 198:21]
  assign array_72_io_ve_i = V1_73; // @[SWChisel.scala 197:22]
  assign array_72_io_vf_i = V1_72; // @[SWChisel.scala 199:22]
  assign array_72_io_vv_i = V2_72; // @[SWChisel.scala 200:22]
  assign array_73_io_q = io_q_73_b; // @[SWChisel.scala 220:19]
  assign array_73_io_r = 8'hc7 == r_count_73_io_out ? io_r_199_b : _GEN_15098; // @[SWChisel.scala 221:{19,19}]
  assign array_73_io_e_i = E_73; // @[SWChisel.scala 196:21]
  assign array_73_io_f_i = F_73; // @[SWChisel.scala 198:21]
  assign array_73_io_ve_i = V1_74; // @[SWChisel.scala 197:22]
  assign array_73_io_vf_i = V1_73; // @[SWChisel.scala 199:22]
  assign array_73_io_vv_i = V2_73; // @[SWChisel.scala 200:22]
  assign array_74_io_q = io_q_74_b; // @[SWChisel.scala 220:19]
  assign array_74_io_r = 8'hc7 == r_count_74_io_out ? io_r_199_b : _GEN_15298; // @[SWChisel.scala 221:{19,19}]
  assign array_74_io_e_i = E_74; // @[SWChisel.scala 196:21]
  assign array_74_io_f_i = F_74; // @[SWChisel.scala 198:21]
  assign array_74_io_ve_i = V1_75; // @[SWChisel.scala 197:22]
  assign array_74_io_vf_i = V1_74; // @[SWChisel.scala 199:22]
  assign array_74_io_vv_i = V2_74; // @[SWChisel.scala 200:22]
  assign array_75_io_q = io_q_75_b; // @[SWChisel.scala 220:19]
  assign array_75_io_r = 8'hc7 == r_count_75_io_out ? io_r_199_b : _GEN_15498; // @[SWChisel.scala 221:{19,19}]
  assign array_75_io_e_i = E_75; // @[SWChisel.scala 196:21]
  assign array_75_io_f_i = F_75; // @[SWChisel.scala 198:21]
  assign array_75_io_ve_i = V1_76; // @[SWChisel.scala 197:22]
  assign array_75_io_vf_i = V1_75; // @[SWChisel.scala 199:22]
  assign array_75_io_vv_i = V2_75; // @[SWChisel.scala 200:22]
  assign array_76_io_q = io_q_76_b; // @[SWChisel.scala 220:19]
  assign array_76_io_r = 8'hc7 == r_count_76_io_out ? io_r_199_b : _GEN_15698; // @[SWChisel.scala 221:{19,19}]
  assign array_76_io_e_i = E_76; // @[SWChisel.scala 196:21]
  assign array_76_io_f_i = F_76; // @[SWChisel.scala 198:21]
  assign array_76_io_ve_i = V1_77; // @[SWChisel.scala 197:22]
  assign array_76_io_vf_i = V1_76; // @[SWChisel.scala 199:22]
  assign array_76_io_vv_i = V2_76; // @[SWChisel.scala 200:22]
  assign array_77_io_q = io_q_77_b; // @[SWChisel.scala 220:19]
  assign array_77_io_r = 8'hc7 == r_count_77_io_out ? io_r_199_b : _GEN_15898; // @[SWChisel.scala 221:{19,19}]
  assign array_77_io_e_i = E_77; // @[SWChisel.scala 196:21]
  assign array_77_io_f_i = F_77; // @[SWChisel.scala 198:21]
  assign array_77_io_ve_i = V1_78; // @[SWChisel.scala 197:22]
  assign array_77_io_vf_i = V1_77; // @[SWChisel.scala 199:22]
  assign array_77_io_vv_i = V2_77; // @[SWChisel.scala 200:22]
  assign array_78_io_q = io_q_78_b; // @[SWChisel.scala 220:19]
  assign array_78_io_r = 8'hc7 == r_count_78_io_out ? io_r_199_b : _GEN_16098; // @[SWChisel.scala 221:{19,19}]
  assign array_78_io_e_i = E_78; // @[SWChisel.scala 196:21]
  assign array_78_io_f_i = F_78; // @[SWChisel.scala 198:21]
  assign array_78_io_ve_i = V1_79; // @[SWChisel.scala 197:22]
  assign array_78_io_vf_i = V1_78; // @[SWChisel.scala 199:22]
  assign array_78_io_vv_i = V2_78; // @[SWChisel.scala 200:22]
  assign array_79_io_q = io_q_79_b; // @[SWChisel.scala 220:19]
  assign array_79_io_r = 8'hc7 == r_count_79_io_out ? io_r_199_b : _GEN_16298; // @[SWChisel.scala 221:{19,19}]
  assign array_79_io_e_i = E_79; // @[SWChisel.scala 196:21]
  assign array_79_io_f_i = F_79; // @[SWChisel.scala 198:21]
  assign array_79_io_ve_i = V1_80; // @[SWChisel.scala 197:22]
  assign array_79_io_vf_i = V1_79; // @[SWChisel.scala 199:22]
  assign array_79_io_vv_i = V2_79; // @[SWChisel.scala 200:22]
  assign array_80_io_q = io_q_80_b; // @[SWChisel.scala 220:19]
  assign array_80_io_r = 8'hc7 == r_count_80_io_out ? io_r_199_b : _GEN_16498; // @[SWChisel.scala 221:{19,19}]
  assign array_80_io_e_i = E_80; // @[SWChisel.scala 196:21]
  assign array_80_io_f_i = F_80; // @[SWChisel.scala 198:21]
  assign array_80_io_ve_i = V1_81; // @[SWChisel.scala 197:22]
  assign array_80_io_vf_i = V1_80; // @[SWChisel.scala 199:22]
  assign array_80_io_vv_i = V2_80; // @[SWChisel.scala 200:22]
  assign array_81_io_q = io_q_81_b; // @[SWChisel.scala 220:19]
  assign array_81_io_r = 8'hc7 == r_count_81_io_out ? io_r_199_b : _GEN_16698; // @[SWChisel.scala 221:{19,19}]
  assign array_81_io_e_i = E_81; // @[SWChisel.scala 196:21]
  assign array_81_io_f_i = F_81; // @[SWChisel.scala 198:21]
  assign array_81_io_ve_i = V1_82; // @[SWChisel.scala 197:22]
  assign array_81_io_vf_i = V1_81; // @[SWChisel.scala 199:22]
  assign array_81_io_vv_i = V2_81; // @[SWChisel.scala 200:22]
  assign array_82_io_q = io_q_82_b; // @[SWChisel.scala 220:19]
  assign array_82_io_r = 8'hc7 == r_count_82_io_out ? io_r_199_b : _GEN_16898; // @[SWChisel.scala 221:{19,19}]
  assign array_82_io_e_i = E_82; // @[SWChisel.scala 196:21]
  assign array_82_io_f_i = F_82; // @[SWChisel.scala 198:21]
  assign array_82_io_ve_i = V1_83; // @[SWChisel.scala 197:22]
  assign array_82_io_vf_i = V1_82; // @[SWChisel.scala 199:22]
  assign array_82_io_vv_i = V2_82; // @[SWChisel.scala 200:22]
  assign array_83_io_q = io_q_83_b; // @[SWChisel.scala 220:19]
  assign array_83_io_r = 8'hc7 == r_count_83_io_out ? io_r_199_b : _GEN_17098; // @[SWChisel.scala 221:{19,19}]
  assign array_83_io_e_i = E_83; // @[SWChisel.scala 196:21]
  assign array_83_io_f_i = F_83; // @[SWChisel.scala 198:21]
  assign array_83_io_ve_i = V1_84; // @[SWChisel.scala 197:22]
  assign array_83_io_vf_i = V1_83; // @[SWChisel.scala 199:22]
  assign array_83_io_vv_i = V2_83; // @[SWChisel.scala 200:22]
  assign array_84_io_q = io_q_84_b; // @[SWChisel.scala 220:19]
  assign array_84_io_r = 8'hc7 == r_count_84_io_out ? io_r_199_b : _GEN_17298; // @[SWChisel.scala 221:{19,19}]
  assign array_84_io_e_i = E_84; // @[SWChisel.scala 196:21]
  assign array_84_io_f_i = F_84; // @[SWChisel.scala 198:21]
  assign array_84_io_ve_i = V1_85; // @[SWChisel.scala 197:22]
  assign array_84_io_vf_i = V1_84; // @[SWChisel.scala 199:22]
  assign array_84_io_vv_i = V2_84; // @[SWChisel.scala 200:22]
  assign array_85_io_q = io_q_85_b; // @[SWChisel.scala 220:19]
  assign array_85_io_r = 8'hc7 == r_count_85_io_out ? io_r_199_b : _GEN_17498; // @[SWChisel.scala 221:{19,19}]
  assign array_85_io_e_i = E_85; // @[SWChisel.scala 196:21]
  assign array_85_io_f_i = F_85; // @[SWChisel.scala 198:21]
  assign array_85_io_ve_i = V1_86; // @[SWChisel.scala 197:22]
  assign array_85_io_vf_i = V1_85; // @[SWChisel.scala 199:22]
  assign array_85_io_vv_i = V2_85; // @[SWChisel.scala 200:22]
  assign array_86_io_q = io_q_86_b; // @[SWChisel.scala 220:19]
  assign array_86_io_r = 8'hc7 == r_count_86_io_out ? io_r_199_b : _GEN_17698; // @[SWChisel.scala 221:{19,19}]
  assign array_86_io_e_i = E_86; // @[SWChisel.scala 196:21]
  assign array_86_io_f_i = F_86; // @[SWChisel.scala 198:21]
  assign array_86_io_ve_i = V1_87; // @[SWChisel.scala 197:22]
  assign array_86_io_vf_i = V1_86; // @[SWChisel.scala 199:22]
  assign array_86_io_vv_i = V2_86; // @[SWChisel.scala 200:22]
  assign array_87_io_q = io_q_87_b; // @[SWChisel.scala 220:19]
  assign array_87_io_r = 8'hc7 == r_count_87_io_out ? io_r_199_b : _GEN_17898; // @[SWChisel.scala 221:{19,19}]
  assign array_87_io_e_i = E_87; // @[SWChisel.scala 196:21]
  assign array_87_io_f_i = F_87; // @[SWChisel.scala 198:21]
  assign array_87_io_ve_i = V1_88; // @[SWChisel.scala 197:22]
  assign array_87_io_vf_i = V1_87; // @[SWChisel.scala 199:22]
  assign array_87_io_vv_i = V2_87; // @[SWChisel.scala 200:22]
  assign array_88_io_q = io_q_88_b; // @[SWChisel.scala 220:19]
  assign array_88_io_r = 8'hc7 == r_count_88_io_out ? io_r_199_b : _GEN_18098; // @[SWChisel.scala 221:{19,19}]
  assign array_88_io_e_i = E_88; // @[SWChisel.scala 196:21]
  assign array_88_io_f_i = F_88; // @[SWChisel.scala 198:21]
  assign array_88_io_ve_i = V1_89; // @[SWChisel.scala 197:22]
  assign array_88_io_vf_i = V1_88; // @[SWChisel.scala 199:22]
  assign array_88_io_vv_i = V2_88; // @[SWChisel.scala 200:22]
  assign array_89_io_q = io_q_89_b; // @[SWChisel.scala 220:19]
  assign array_89_io_r = 8'hc7 == r_count_89_io_out ? io_r_199_b : _GEN_18298; // @[SWChisel.scala 221:{19,19}]
  assign array_89_io_e_i = E_89; // @[SWChisel.scala 196:21]
  assign array_89_io_f_i = F_89; // @[SWChisel.scala 198:21]
  assign array_89_io_ve_i = V1_90; // @[SWChisel.scala 197:22]
  assign array_89_io_vf_i = V1_89; // @[SWChisel.scala 199:22]
  assign array_89_io_vv_i = V2_89; // @[SWChisel.scala 200:22]
  assign array_90_io_q = io_q_90_b; // @[SWChisel.scala 220:19]
  assign array_90_io_r = 8'hc7 == r_count_90_io_out ? io_r_199_b : _GEN_18498; // @[SWChisel.scala 221:{19,19}]
  assign array_90_io_e_i = E_90; // @[SWChisel.scala 196:21]
  assign array_90_io_f_i = F_90; // @[SWChisel.scala 198:21]
  assign array_90_io_ve_i = V1_91; // @[SWChisel.scala 197:22]
  assign array_90_io_vf_i = V1_90; // @[SWChisel.scala 199:22]
  assign array_90_io_vv_i = V2_90; // @[SWChisel.scala 200:22]
  assign array_91_io_q = io_q_91_b; // @[SWChisel.scala 220:19]
  assign array_91_io_r = 8'hc7 == r_count_91_io_out ? io_r_199_b : _GEN_18698; // @[SWChisel.scala 221:{19,19}]
  assign array_91_io_e_i = E_91; // @[SWChisel.scala 196:21]
  assign array_91_io_f_i = F_91; // @[SWChisel.scala 198:21]
  assign array_91_io_ve_i = V1_92; // @[SWChisel.scala 197:22]
  assign array_91_io_vf_i = V1_91; // @[SWChisel.scala 199:22]
  assign array_91_io_vv_i = V2_91; // @[SWChisel.scala 200:22]
  assign array_92_io_q = io_q_92_b; // @[SWChisel.scala 220:19]
  assign array_92_io_r = 8'hc7 == r_count_92_io_out ? io_r_199_b : _GEN_18898; // @[SWChisel.scala 221:{19,19}]
  assign array_92_io_e_i = E_92; // @[SWChisel.scala 196:21]
  assign array_92_io_f_i = F_92; // @[SWChisel.scala 198:21]
  assign array_92_io_ve_i = V1_93; // @[SWChisel.scala 197:22]
  assign array_92_io_vf_i = V1_92; // @[SWChisel.scala 199:22]
  assign array_92_io_vv_i = V2_92; // @[SWChisel.scala 200:22]
  assign array_93_io_q = io_q_93_b; // @[SWChisel.scala 220:19]
  assign array_93_io_r = 8'hc7 == r_count_93_io_out ? io_r_199_b : _GEN_19098; // @[SWChisel.scala 221:{19,19}]
  assign array_93_io_e_i = E_93; // @[SWChisel.scala 196:21]
  assign array_93_io_f_i = F_93; // @[SWChisel.scala 198:21]
  assign array_93_io_ve_i = V1_94; // @[SWChisel.scala 197:22]
  assign array_93_io_vf_i = V1_93; // @[SWChisel.scala 199:22]
  assign array_93_io_vv_i = V2_93; // @[SWChisel.scala 200:22]
  assign array_94_io_q = io_q_94_b; // @[SWChisel.scala 220:19]
  assign array_94_io_r = 8'hc7 == r_count_94_io_out ? io_r_199_b : _GEN_19298; // @[SWChisel.scala 221:{19,19}]
  assign array_94_io_e_i = E_94; // @[SWChisel.scala 196:21]
  assign array_94_io_f_i = F_94; // @[SWChisel.scala 198:21]
  assign array_94_io_ve_i = V1_95; // @[SWChisel.scala 197:22]
  assign array_94_io_vf_i = V1_94; // @[SWChisel.scala 199:22]
  assign array_94_io_vv_i = V2_94; // @[SWChisel.scala 200:22]
  assign array_95_io_q = io_q_95_b; // @[SWChisel.scala 220:19]
  assign array_95_io_r = 8'hc7 == r_count_95_io_out ? io_r_199_b : _GEN_19498; // @[SWChisel.scala 221:{19,19}]
  assign array_95_io_e_i = E_95; // @[SWChisel.scala 196:21]
  assign array_95_io_f_i = F_95; // @[SWChisel.scala 198:21]
  assign array_95_io_ve_i = V1_96; // @[SWChisel.scala 197:22]
  assign array_95_io_vf_i = V1_95; // @[SWChisel.scala 199:22]
  assign array_95_io_vv_i = V2_95; // @[SWChisel.scala 200:22]
  assign array_96_io_q = io_q_96_b; // @[SWChisel.scala 220:19]
  assign array_96_io_r = 8'hc7 == r_count_96_io_out ? io_r_199_b : _GEN_19698; // @[SWChisel.scala 221:{19,19}]
  assign array_96_io_e_i = E_96; // @[SWChisel.scala 196:21]
  assign array_96_io_f_i = F_96; // @[SWChisel.scala 198:21]
  assign array_96_io_ve_i = V1_97; // @[SWChisel.scala 197:22]
  assign array_96_io_vf_i = V1_96; // @[SWChisel.scala 199:22]
  assign array_96_io_vv_i = V2_96; // @[SWChisel.scala 200:22]
  assign array_97_io_q = io_q_97_b; // @[SWChisel.scala 220:19]
  assign array_97_io_r = 8'hc7 == r_count_97_io_out ? io_r_199_b : _GEN_19898; // @[SWChisel.scala 221:{19,19}]
  assign array_97_io_e_i = E_97; // @[SWChisel.scala 196:21]
  assign array_97_io_f_i = F_97; // @[SWChisel.scala 198:21]
  assign array_97_io_ve_i = V1_98; // @[SWChisel.scala 197:22]
  assign array_97_io_vf_i = V1_97; // @[SWChisel.scala 199:22]
  assign array_97_io_vv_i = V2_97; // @[SWChisel.scala 200:22]
  assign array_98_io_q = io_q_98_b; // @[SWChisel.scala 220:19]
  assign array_98_io_r = 8'hc7 == r_count_98_io_out ? io_r_199_b : _GEN_20098; // @[SWChisel.scala 221:{19,19}]
  assign array_98_io_e_i = E_98; // @[SWChisel.scala 196:21]
  assign array_98_io_f_i = F_98; // @[SWChisel.scala 198:21]
  assign array_98_io_ve_i = V1_99; // @[SWChisel.scala 197:22]
  assign array_98_io_vf_i = V1_98; // @[SWChisel.scala 199:22]
  assign array_98_io_vv_i = V2_98; // @[SWChisel.scala 200:22]
  assign array_99_io_q = io_q_99_b; // @[SWChisel.scala 220:19]
  assign array_99_io_r = 8'hc7 == r_count_99_io_out ? io_r_199_b : _GEN_20298; // @[SWChisel.scala 221:{19,19}]
  assign array_99_io_e_i = E_99; // @[SWChisel.scala 196:21]
  assign array_99_io_f_i = F_99; // @[SWChisel.scala 198:21]
  assign array_99_io_ve_i = V1_100; // @[SWChisel.scala 197:22]
  assign array_99_io_vf_i = V1_99; // @[SWChisel.scala 199:22]
  assign array_99_io_vv_i = V2_99; // @[SWChisel.scala 200:22]
  assign r_count_0_clock = clock;
  assign r_count_0_reset = reset;
  assign r_count_0_io_en = start_reg_0; // @[SWChisel.scala 192:22]
  assign r_count_1_clock = clock;
  assign r_count_1_reset = reset;
  assign r_count_1_io_en = start_reg_1; // @[SWChisel.scala 192:22]
  assign r_count_2_clock = clock;
  assign r_count_2_reset = reset;
  assign r_count_2_io_en = start_reg_2; // @[SWChisel.scala 192:22]
  assign r_count_3_clock = clock;
  assign r_count_3_reset = reset;
  assign r_count_3_io_en = start_reg_3; // @[SWChisel.scala 192:22]
  assign r_count_4_clock = clock;
  assign r_count_4_reset = reset;
  assign r_count_4_io_en = start_reg_4; // @[SWChisel.scala 192:22]
  assign r_count_5_clock = clock;
  assign r_count_5_reset = reset;
  assign r_count_5_io_en = start_reg_5; // @[SWChisel.scala 192:22]
  assign r_count_6_clock = clock;
  assign r_count_6_reset = reset;
  assign r_count_6_io_en = start_reg_6; // @[SWChisel.scala 192:22]
  assign r_count_7_clock = clock;
  assign r_count_7_reset = reset;
  assign r_count_7_io_en = start_reg_7; // @[SWChisel.scala 192:22]
  assign r_count_8_clock = clock;
  assign r_count_8_reset = reset;
  assign r_count_8_io_en = start_reg_8; // @[SWChisel.scala 192:22]
  assign r_count_9_clock = clock;
  assign r_count_9_reset = reset;
  assign r_count_9_io_en = start_reg_9; // @[SWChisel.scala 192:22]
  assign r_count_10_clock = clock;
  assign r_count_10_reset = reset;
  assign r_count_10_io_en = start_reg_10; // @[SWChisel.scala 192:22]
  assign r_count_11_clock = clock;
  assign r_count_11_reset = reset;
  assign r_count_11_io_en = start_reg_11; // @[SWChisel.scala 192:22]
  assign r_count_12_clock = clock;
  assign r_count_12_reset = reset;
  assign r_count_12_io_en = start_reg_12; // @[SWChisel.scala 192:22]
  assign r_count_13_clock = clock;
  assign r_count_13_reset = reset;
  assign r_count_13_io_en = start_reg_13; // @[SWChisel.scala 192:22]
  assign r_count_14_clock = clock;
  assign r_count_14_reset = reset;
  assign r_count_14_io_en = start_reg_14; // @[SWChisel.scala 192:22]
  assign r_count_15_clock = clock;
  assign r_count_15_reset = reset;
  assign r_count_15_io_en = start_reg_15; // @[SWChisel.scala 192:22]
  assign r_count_16_clock = clock;
  assign r_count_16_reset = reset;
  assign r_count_16_io_en = start_reg_16; // @[SWChisel.scala 192:22]
  assign r_count_17_clock = clock;
  assign r_count_17_reset = reset;
  assign r_count_17_io_en = start_reg_17; // @[SWChisel.scala 192:22]
  assign r_count_18_clock = clock;
  assign r_count_18_reset = reset;
  assign r_count_18_io_en = start_reg_18; // @[SWChisel.scala 192:22]
  assign r_count_19_clock = clock;
  assign r_count_19_reset = reset;
  assign r_count_19_io_en = start_reg_19; // @[SWChisel.scala 192:22]
  assign r_count_20_clock = clock;
  assign r_count_20_reset = reset;
  assign r_count_20_io_en = start_reg_20; // @[SWChisel.scala 192:22]
  assign r_count_21_clock = clock;
  assign r_count_21_reset = reset;
  assign r_count_21_io_en = start_reg_21; // @[SWChisel.scala 192:22]
  assign r_count_22_clock = clock;
  assign r_count_22_reset = reset;
  assign r_count_22_io_en = start_reg_22; // @[SWChisel.scala 192:22]
  assign r_count_23_clock = clock;
  assign r_count_23_reset = reset;
  assign r_count_23_io_en = start_reg_23; // @[SWChisel.scala 192:22]
  assign r_count_24_clock = clock;
  assign r_count_24_reset = reset;
  assign r_count_24_io_en = start_reg_24; // @[SWChisel.scala 192:22]
  assign r_count_25_clock = clock;
  assign r_count_25_reset = reset;
  assign r_count_25_io_en = start_reg_25; // @[SWChisel.scala 192:22]
  assign r_count_26_clock = clock;
  assign r_count_26_reset = reset;
  assign r_count_26_io_en = start_reg_26; // @[SWChisel.scala 192:22]
  assign r_count_27_clock = clock;
  assign r_count_27_reset = reset;
  assign r_count_27_io_en = start_reg_27; // @[SWChisel.scala 192:22]
  assign r_count_28_clock = clock;
  assign r_count_28_reset = reset;
  assign r_count_28_io_en = start_reg_28; // @[SWChisel.scala 192:22]
  assign r_count_29_clock = clock;
  assign r_count_29_reset = reset;
  assign r_count_29_io_en = start_reg_29; // @[SWChisel.scala 192:22]
  assign r_count_30_clock = clock;
  assign r_count_30_reset = reset;
  assign r_count_30_io_en = start_reg_30; // @[SWChisel.scala 192:22]
  assign r_count_31_clock = clock;
  assign r_count_31_reset = reset;
  assign r_count_31_io_en = start_reg_31; // @[SWChisel.scala 192:22]
  assign r_count_32_clock = clock;
  assign r_count_32_reset = reset;
  assign r_count_32_io_en = start_reg_32; // @[SWChisel.scala 192:22]
  assign r_count_33_clock = clock;
  assign r_count_33_reset = reset;
  assign r_count_33_io_en = start_reg_33; // @[SWChisel.scala 192:22]
  assign r_count_34_clock = clock;
  assign r_count_34_reset = reset;
  assign r_count_34_io_en = start_reg_34; // @[SWChisel.scala 192:22]
  assign r_count_35_clock = clock;
  assign r_count_35_reset = reset;
  assign r_count_35_io_en = start_reg_35; // @[SWChisel.scala 192:22]
  assign r_count_36_clock = clock;
  assign r_count_36_reset = reset;
  assign r_count_36_io_en = start_reg_36; // @[SWChisel.scala 192:22]
  assign r_count_37_clock = clock;
  assign r_count_37_reset = reset;
  assign r_count_37_io_en = start_reg_37; // @[SWChisel.scala 192:22]
  assign r_count_38_clock = clock;
  assign r_count_38_reset = reset;
  assign r_count_38_io_en = start_reg_38; // @[SWChisel.scala 192:22]
  assign r_count_39_clock = clock;
  assign r_count_39_reset = reset;
  assign r_count_39_io_en = start_reg_39; // @[SWChisel.scala 192:22]
  assign r_count_40_clock = clock;
  assign r_count_40_reset = reset;
  assign r_count_40_io_en = start_reg_40; // @[SWChisel.scala 192:22]
  assign r_count_41_clock = clock;
  assign r_count_41_reset = reset;
  assign r_count_41_io_en = start_reg_41; // @[SWChisel.scala 192:22]
  assign r_count_42_clock = clock;
  assign r_count_42_reset = reset;
  assign r_count_42_io_en = start_reg_42; // @[SWChisel.scala 192:22]
  assign r_count_43_clock = clock;
  assign r_count_43_reset = reset;
  assign r_count_43_io_en = start_reg_43; // @[SWChisel.scala 192:22]
  assign r_count_44_clock = clock;
  assign r_count_44_reset = reset;
  assign r_count_44_io_en = start_reg_44; // @[SWChisel.scala 192:22]
  assign r_count_45_clock = clock;
  assign r_count_45_reset = reset;
  assign r_count_45_io_en = start_reg_45; // @[SWChisel.scala 192:22]
  assign r_count_46_clock = clock;
  assign r_count_46_reset = reset;
  assign r_count_46_io_en = start_reg_46; // @[SWChisel.scala 192:22]
  assign r_count_47_clock = clock;
  assign r_count_47_reset = reset;
  assign r_count_47_io_en = start_reg_47; // @[SWChisel.scala 192:22]
  assign r_count_48_clock = clock;
  assign r_count_48_reset = reset;
  assign r_count_48_io_en = start_reg_48; // @[SWChisel.scala 192:22]
  assign r_count_49_clock = clock;
  assign r_count_49_reset = reset;
  assign r_count_49_io_en = start_reg_49; // @[SWChisel.scala 192:22]
  assign r_count_50_clock = clock;
  assign r_count_50_reset = reset;
  assign r_count_50_io_en = start_reg_50; // @[SWChisel.scala 192:22]
  assign r_count_51_clock = clock;
  assign r_count_51_reset = reset;
  assign r_count_51_io_en = start_reg_51; // @[SWChisel.scala 192:22]
  assign r_count_52_clock = clock;
  assign r_count_52_reset = reset;
  assign r_count_52_io_en = start_reg_52; // @[SWChisel.scala 192:22]
  assign r_count_53_clock = clock;
  assign r_count_53_reset = reset;
  assign r_count_53_io_en = start_reg_53; // @[SWChisel.scala 192:22]
  assign r_count_54_clock = clock;
  assign r_count_54_reset = reset;
  assign r_count_54_io_en = start_reg_54; // @[SWChisel.scala 192:22]
  assign r_count_55_clock = clock;
  assign r_count_55_reset = reset;
  assign r_count_55_io_en = start_reg_55; // @[SWChisel.scala 192:22]
  assign r_count_56_clock = clock;
  assign r_count_56_reset = reset;
  assign r_count_56_io_en = start_reg_56; // @[SWChisel.scala 192:22]
  assign r_count_57_clock = clock;
  assign r_count_57_reset = reset;
  assign r_count_57_io_en = start_reg_57; // @[SWChisel.scala 192:22]
  assign r_count_58_clock = clock;
  assign r_count_58_reset = reset;
  assign r_count_58_io_en = start_reg_58; // @[SWChisel.scala 192:22]
  assign r_count_59_clock = clock;
  assign r_count_59_reset = reset;
  assign r_count_59_io_en = start_reg_59; // @[SWChisel.scala 192:22]
  assign r_count_60_clock = clock;
  assign r_count_60_reset = reset;
  assign r_count_60_io_en = start_reg_60; // @[SWChisel.scala 192:22]
  assign r_count_61_clock = clock;
  assign r_count_61_reset = reset;
  assign r_count_61_io_en = start_reg_61; // @[SWChisel.scala 192:22]
  assign r_count_62_clock = clock;
  assign r_count_62_reset = reset;
  assign r_count_62_io_en = start_reg_62; // @[SWChisel.scala 192:22]
  assign r_count_63_clock = clock;
  assign r_count_63_reset = reset;
  assign r_count_63_io_en = start_reg_63; // @[SWChisel.scala 192:22]
  assign r_count_64_clock = clock;
  assign r_count_64_reset = reset;
  assign r_count_64_io_en = start_reg_64; // @[SWChisel.scala 192:22]
  assign r_count_65_clock = clock;
  assign r_count_65_reset = reset;
  assign r_count_65_io_en = start_reg_65; // @[SWChisel.scala 192:22]
  assign r_count_66_clock = clock;
  assign r_count_66_reset = reset;
  assign r_count_66_io_en = start_reg_66; // @[SWChisel.scala 192:22]
  assign r_count_67_clock = clock;
  assign r_count_67_reset = reset;
  assign r_count_67_io_en = start_reg_67; // @[SWChisel.scala 192:22]
  assign r_count_68_clock = clock;
  assign r_count_68_reset = reset;
  assign r_count_68_io_en = start_reg_68; // @[SWChisel.scala 192:22]
  assign r_count_69_clock = clock;
  assign r_count_69_reset = reset;
  assign r_count_69_io_en = start_reg_69; // @[SWChisel.scala 192:22]
  assign r_count_70_clock = clock;
  assign r_count_70_reset = reset;
  assign r_count_70_io_en = start_reg_70; // @[SWChisel.scala 192:22]
  assign r_count_71_clock = clock;
  assign r_count_71_reset = reset;
  assign r_count_71_io_en = start_reg_71; // @[SWChisel.scala 192:22]
  assign r_count_72_clock = clock;
  assign r_count_72_reset = reset;
  assign r_count_72_io_en = start_reg_72; // @[SWChisel.scala 192:22]
  assign r_count_73_clock = clock;
  assign r_count_73_reset = reset;
  assign r_count_73_io_en = start_reg_73; // @[SWChisel.scala 192:22]
  assign r_count_74_clock = clock;
  assign r_count_74_reset = reset;
  assign r_count_74_io_en = start_reg_74; // @[SWChisel.scala 192:22]
  assign r_count_75_clock = clock;
  assign r_count_75_reset = reset;
  assign r_count_75_io_en = start_reg_75; // @[SWChisel.scala 192:22]
  assign r_count_76_clock = clock;
  assign r_count_76_reset = reset;
  assign r_count_76_io_en = start_reg_76; // @[SWChisel.scala 192:22]
  assign r_count_77_clock = clock;
  assign r_count_77_reset = reset;
  assign r_count_77_io_en = start_reg_77; // @[SWChisel.scala 192:22]
  assign r_count_78_clock = clock;
  assign r_count_78_reset = reset;
  assign r_count_78_io_en = start_reg_78; // @[SWChisel.scala 192:22]
  assign r_count_79_clock = clock;
  assign r_count_79_reset = reset;
  assign r_count_79_io_en = start_reg_79; // @[SWChisel.scala 192:22]
  assign r_count_80_clock = clock;
  assign r_count_80_reset = reset;
  assign r_count_80_io_en = start_reg_80; // @[SWChisel.scala 192:22]
  assign r_count_81_clock = clock;
  assign r_count_81_reset = reset;
  assign r_count_81_io_en = start_reg_81; // @[SWChisel.scala 192:22]
  assign r_count_82_clock = clock;
  assign r_count_82_reset = reset;
  assign r_count_82_io_en = start_reg_82; // @[SWChisel.scala 192:22]
  assign r_count_83_clock = clock;
  assign r_count_83_reset = reset;
  assign r_count_83_io_en = start_reg_83; // @[SWChisel.scala 192:22]
  assign r_count_84_clock = clock;
  assign r_count_84_reset = reset;
  assign r_count_84_io_en = start_reg_84; // @[SWChisel.scala 192:22]
  assign r_count_85_clock = clock;
  assign r_count_85_reset = reset;
  assign r_count_85_io_en = start_reg_85; // @[SWChisel.scala 192:22]
  assign r_count_86_clock = clock;
  assign r_count_86_reset = reset;
  assign r_count_86_io_en = start_reg_86; // @[SWChisel.scala 192:22]
  assign r_count_87_clock = clock;
  assign r_count_87_reset = reset;
  assign r_count_87_io_en = start_reg_87; // @[SWChisel.scala 192:22]
  assign r_count_88_clock = clock;
  assign r_count_88_reset = reset;
  assign r_count_88_io_en = start_reg_88; // @[SWChisel.scala 192:22]
  assign r_count_89_clock = clock;
  assign r_count_89_reset = reset;
  assign r_count_89_io_en = start_reg_89; // @[SWChisel.scala 192:22]
  assign r_count_90_clock = clock;
  assign r_count_90_reset = reset;
  assign r_count_90_io_en = start_reg_90; // @[SWChisel.scala 192:22]
  assign r_count_91_clock = clock;
  assign r_count_91_reset = reset;
  assign r_count_91_io_en = start_reg_91; // @[SWChisel.scala 192:22]
  assign r_count_92_clock = clock;
  assign r_count_92_reset = reset;
  assign r_count_92_io_en = start_reg_92; // @[SWChisel.scala 192:22]
  assign r_count_93_clock = clock;
  assign r_count_93_reset = reset;
  assign r_count_93_io_en = start_reg_93; // @[SWChisel.scala 192:22]
  assign r_count_94_clock = clock;
  assign r_count_94_reset = reset;
  assign r_count_94_io_en = start_reg_94; // @[SWChisel.scala 192:22]
  assign r_count_95_clock = clock;
  assign r_count_95_reset = reset;
  assign r_count_95_io_en = start_reg_95; // @[SWChisel.scala 192:22]
  assign r_count_96_clock = clock;
  assign r_count_96_reset = reset;
  assign r_count_96_io_en = start_reg_96; // @[SWChisel.scala 192:22]
  assign r_count_97_clock = clock;
  assign r_count_97_reset = reset;
  assign r_count_97_io_en = start_reg_97; // @[SWChisel.scala 192:22]
  assign r_count_98_clock = clock;
  assign r_count_98_reset = reset;
  assign r_count_98_io_en = start_reg_98; // @[SWChisel.scala 192:22]
  assign r_count_99_clock = clock;
  assign r_count_99_reset = reset;
  assign r_count_99_io_en = start_reg_99; // @[SWChisel.scala 192:22]
  assign max_clock = clock;
  assign max_reset = reset;
  assign max_io_start = start_reg_99; // @[SWChisel.scala 178:16]
  assign max_io_in = V1_100; // @[SWChisel.scala 177:13]
  always @(posedge clock) begin
    if (reset) begin // @[SWChisel.scala 162:18]
      E_0 <= -16'sh2; // @[SWChisel.scala 162:18]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      E_0 <= array_0_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_1 <= -16'sh3; // @[SWChisel.scala 162:18]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      E_1 <= array_1_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_2 <= -16'sh4; // @[SWChisel.scala 162:18]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      E_2 <= array_2_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_3 <= -16'sh5; // @[SWChisel.scala 162:18]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      E_3 <= array_3_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_4 <= -16'sh6; // @[SWChisel.scala 162:18]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      E_4 <= array_4_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_5 <= -16'sh7; // @[SWChisel.scala 162:18]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      E_5 <= array_5_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_6 <= -16'sh8; // @[SWChisel.scala 162:18]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      E_6 <= array_6_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_7 <= -16'sh9; // @[SWChisel.scala 162:18]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      E_7 <= array_7_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_8 <= -16'sha; // @[SWChisel.scala 162:18]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      E_8 <= array_8_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_9 <= -16'shb; // @[SWChisel.scala 162:18]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      E_9 <= array_9_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_10 <= -16'shc; // @[SWChisel.scala 162:18]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      E_10 <= array_10_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_11 <= -16'shd; // @[SWChisel.scala 162:18]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      E_11 <= array_11_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_12 <= -16'she; // @[SWChisel.scala 162:18]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      E_12 <= array_12_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_13 <= -16'shf; // @[SWChisel.scala 162:18]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      E_13 <= array_13_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_14 <= -16'sh10; // @[SWChisel.scala 162:18]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      E_14 <= array_14_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_15 <= -16'sh11; // @[SWChisel.scala 162:18]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      E_15 <= array_15_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_16 <= -16'sh12; // @[SWChisel.scala 162:18]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      E_16 <= array_16_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_17 <= -16'sh13; // @[SWChisel.scala 162:18]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      E_17 <= array_17_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_18 <= -16'sh14; // @[SWChisel.scala 162:18]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      E_18 <= array_18_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_19 <= -16'sh15; // @[SWChisel.scala 162:18]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      E_19 <= array_19_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_20 <= -16'sh16; // @[SWChisel.scala 162:18]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      E_20 <= array_20_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_21 <= -16'sh17; // @[SWChisel.scala 162:18]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      E_21 <= array_21_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_22 <= -16'sh18; // @[SWChisel.scala 162:18]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      E_22 <= array_22_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_23 <= -16'sh19; // @[SWChisel.scala 162:18]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      E_23 <= array_23_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_24 <= -16'sh1a; // @[SWChisel.scala 162:18]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      E_24 <= array_24_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_25 <= -16'sh1b; // @[SWChisel.scala 162:18]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      E_25 <= array_25_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_26 <= -16'sh1c; // @[SWChisel.scala 162:18]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      E_26 <= array_26_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_27 <= -16'sh1d; // @[SWChisel.scala 162:18]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      E_27 <= array_27_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_28 <= -16'sh1e; // @[SWChisel.scala 162:18]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      E_28 <= array_28_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_29 <= -16'sh1f; // @[SWChisel.scala 162:18]
    end else if (start_reg_29) begin // @[SWChisel.scala 207:25]
      E_29 <= array_29_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_30 <= -16'sh20; // @[SWChisel.scala 162:18]
    end else if (start_reg_30) begin // @[SWChisel.scala 207:25]
      E_30 <= array_30_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_31 <= -16'sh21; // @[SWChisel.scala 162:18]
    end else if (start_reg_31) begin // @[SWChisel.scala 207:25]
      E_31 <= array_31_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_32 <= -16'sh22; // @[SWChisel.scala 162:18]
    end else if (start_reg_32) begin // @[SWChisel.scala 207:25]
      E_32 <= array_32_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_33 <= -16'sh23; // @[SWChisel.scala 162:18]
    end else if (start_reg_33) begin // @[SWChisel.scala 207:25]
      E_33 <= array_33_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_34 <= -16'sh24; // @[SWChisel.scala 162:18]
    end else if (start_reg_34) begin // @[SWChisel.scala 207:25]
      E_34 <= array_34_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_35 <= -16'sh25; // @[SWChisel.scala 162:18]
    end else if (start_reg_35) begin // @[SWChisel.scala 207:25]
      E_35 <= array_35_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_36 <= -16'sh26; // @[SWChisel.scala 162:18]
    end else if (start_reg_36) begin // @[SWChisel.scala 207:25]
      E_36 <= array_36_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_37 <= -16'sh27; // @[SWChisel.scala 162:18]
    end else if (start_reg_37) begin // @[SWChisel.scala 207:25]
      E_37 <= array_37_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_38 <= -16'sh28; // @[SWChisel.scala 162:18]
    end else if (start_reg_38) begin // @[SWChisel.scala 207:25]
      E_38 <= array_38_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_39 <= -16'sh29; // @[SWChisel.scala 162:18]
    end else if (start_reg_39) begin // @[SWChisel.scala 207:25]
      E_39 <= array_39_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_40 <= -16'sh2a; // @[SWChisel.scala 162:18]
    end else if (start_reg_40) begin // @[SWChisel.scala 207:25]
      E_40 <= array_40_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_41 <= -16'sh2b; // @[SWChisel.scala 162:18]
    end else if (start_reg_41) begin // @[SWChisel.scala 207:25]
      E_41 <= array_41_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_42 <= -16'sh2c; // @[SWChisel.scala 162:18]
    end else if (start_reg_42) begin // @[SWChisel.scala 207:25]
      E_42 <= array_42_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_43 <= -16'sh2d; // @[SWChisel.scala 162:18]
    end else if (start_reg_43) begin // @[SWChisel.scala 207:25]
      E_43 <= array_43_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_44 <= -16'sh2e; // @[SWChisel.scala 162:18]
    end else if (start_reg_44) begin // @[SWChisel.scala 207:25]
      E_44 <= array_44_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_45 <= -16'sh2f; // @[SWChisel.scala 162:18]
    end else if (start_reg_45) begin // @[SWChisel.scala 207:25]
      E_45 <= array_45_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_46 <= -16'sh30; // @[SWChisel.scala 162:18]
    end else if (start_reg_46) begin // @[SWChisel.scala 207:25]
      E_46 <= array_46_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_47 <= -16'sh31; // @[SWChisel.scala 162:18]
    end else if (start_reg_47) begin // @[SWChisel.scala 207:25]
      E_47 <= array_47_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_48 <= -16'sh32; // @[SWChisel.scala 162:18]
    end else if (start_reg_48) begin // @[SWChisel.scala 207:25]
      E_48 <= array_48_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_49 <= -16'sh33; // @[SWChisel.scala 162:18]
    end else if (start_reg_49) begin // @[SWChisel.scala 207:25]
      E_49 <= array_49_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_50 <= -16'sh34; // @[SWChisel.scala 162:18]
    end else if (start_reg_50) begin // @[SWChisel.scala 207:25]
      E_50 <= array_50_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_51 <= -16'sh35; // @[SWChisel.scala 162:18]
    end else if (start_reg_51) begin // @[SWChisel.scala 207:25]
      E_51 <= array_51_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_52 <= -16'sh36; // @[SWChisel.scala 162:18]
    end else if (start_reg_52) begin // @[SWChisel.scala 207:25]
      E_52 <= array_52_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_53 <= -16'sh37; // @[SWChisel.scala 162:18]
    end else if (start_reg_53) begin // @[SWChisel.scala 207:25]
      E_53 <= array_53_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_54 <= -16'sh38; // @[SWChisel.scala 162:18]
    end else if (start_reg_54) begin // @[SWChisel.scala 207:25]
      E_54 <= array_54_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_55 <= -16'sh39; // @[SWChisel.scala 162:18]
    end else if (start_reg_55) begin // @[SWChisel.scala 207:25]
      E_55 <= array_55_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_56 <= -16'sh3a; // @[SWChisel.scala 162:18]
    end else if (start_reg_56) begin // @[SWChisel.scala 207:25]
      E_56 <= array_56_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_57 <= -16'sh3b; // @[SWChisel.scala 162:18]
    end else if (start_reg_57) begin // @[SWChisel.scala 207:25]
      E_57 <= array_57_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_58 <= -16'sh3c; // @[SWChisel.scala 162:18]
    end else if (start_reg_58) begin // @[SWChisel.scala 207:25]
      E_58 <= array_58_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_59 <= -16'sh3d; // @[SWChisel.scala 162:18]
    end else if (start_reg_59) begin // @[SWChisel.scala 207:25]
      E_59 <= array_59_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_60 <= -16'sh3e; // @[SWChisel.scala 162:18]
    end else if (start_reg_60) begin // @[SWChisel.scala 207:25]
      E_60 <= array_60_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_61 <= -16'sh3f; // @[SWChisel.scala 162:18]
    end else if (start_reg_61) begin // @[SWChisel.scala 207:25]
      E_61 <= array_61_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_62 <= -16'sh40; // @[SWChisel.scala 162:18]
    end else if (start_reg_62) begin // @[SWChisel.scala 207:25]
      E_62 <= array_62_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_63 <= -16'sh41; // @[SWChisel.scala 162:18]
    end else if (start_reg_63) begin // @[SWChisel.scala 207:25]
      E_63 <= array_63_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_64 <= -16'sh42; // @[SWChisel.scala 162:18]
    end else if (start_reg_64) begin // @[SWChisel.scala 207:25]
      E_64 <= array_64_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_65 <= -16'sh43; // @[SWChisel.scala 162:18]
    end else if (start_reg_65) begin // @[SWChisel.scala 207:25]
      E_65 <= array_65_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_66 <= -16'sh44; // @[SWChisel.scala 162:18]
    end else if (start_reg_66) begin // @[SWChisel.scala 207:25]
      E_66 <= array_66_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_67 <= -16'sh45; // @[SWChisel.scala 162:18]
    end else if (start_reg_67) begin // @[SWChisel.scala 207:25]
      E_67 <= array_67_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_68 <= -16'sh46; // @[SWChisel.scala 162:18]
    end else if (start_reg_68) begin // @[SWChisel.scala 207:25]
      E_68 <= array_68_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_69 <= -16'sh47; // @[SWChisel.scala 162:18]
    end else if (start_reg_69) begin // @[SWChisel.scala 207:25]
      E_69 <= array_69_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_70 <= -16'sh48; // @[SWChisel.scala 162:18]
    end else if (start_reg_70) begin // @[SWChisel.scala 207:25]
      E_70 <= array_70_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_71 <= -16'sh49; // @[SWChisel.scala 162:18]
    end else if (start_reg_71) begin // @[SWChisel.scala 207:25]
      E_71 <= array_71_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_72 <= -16'sh4a; // @[SWChisel.scala 162:18]
    end else if (start_reg_72) begin // @[SWChisel.scala 207:25]
      E_72 <= array_72_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_73 <= -16'sh4b; // @[SWChisel.scala 162:18]
    end else if (start_reg_73) begin // @[SWChisel.scala 207:25]
      E_73 <= array_73_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_74 <= -16'sh4c; // @[SWChisel.scala 162:18]
    end else if (start_reg_74) begin // @[SWChisel.scala 207:25]
      E_74 <= array_74_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_75 <= -16'sh4d; // @[SWChisel.scala 162:18]
    end else if (start_reg_75) begin // @[SWChisel.scala 207:25]
      E_75 <= array_75_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_76 <= -16'sh4e; // @[SWChisel.scala 162:18]
    end else if (start_reg_76) begin // @[SWChisel.scala 207:25]
      E_76 <= array_76_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_77 <= -16'sh4f; // @[SWChisel.scala 162:18]
    end else if (start_reg_77) begin // @[SWChisel.scala 207:25]
      E_77 <= array_77_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_78 <= -16'sh50; // @[SWChisel.scala 162:18]
    end else if (start_reg_78) begin // @[SWChisel.scala 207:25]
      E_78 <= array_78_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_79 <= -16'sh51; // @[SWChisel.scala 162:18]
    end else if (start_reg_79) begin // @[SWChisel.scala 207:25]
      E_79 <= array_79_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_80 <= -16'sh52; // @[SWChisel.scala 162:18]
    end else if (start_reg_80) begin // @[SWChisel.scala 207:25]
      E_80 <= array_80_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_81 <= -16'sh53; // @[SWChisel.scala 162:18]
    end else if (start_reg_81) begin // @[SWChisel.scala 207:25]
      E_81 <= array_81_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_82 <= -16'sh54; // @[SWChisel.scala 162:18]
    end else if (start_reg_82) begin // @[SWChisel.scala 207:25]
      E_82 <= array_82_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_83 <= -16'sh55; // @[SWChisel.scala 162:18]
    end else if (start_reg_83) begin // @[SWChisel.scala 207:25]
      E_83 <= array_83_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_84 <= -16'sh56; // @[SWChisel.scala 162:18]
    end else if (start_reg_84) begin // @[SWChisel.scala 207:25]
      E_84 <= array_84_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_85 <= -16'sh57; // @[SWChisel.scala 162:18]
    end else if (start_reg_85) begin // @[SWChisel.scala 207:25]
      E_85 <= array_85_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_86 <= -16'sh58; // @[SWChisel.scala 162:18]
    end else if (start_reg_86) begin // @[SWChisel.scala 207:25]
      E_86 <= array_86_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_87 <= -16'sh59; // @[SWChisel.scala 162:18]
    end else if (start_reg_87) begin // @[SWChisel.scala 207:25]
      E_87 <= array_87_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_88 <= -16'sh5a; // @[SWChisel.scala 162:18]
    end else if (start_reg_88) begin // @[SWChisel.scala 207:25]
      E_88 <= array_88_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_89 <= -16'sh5b; // @[SWChisel.scala 162:18]
    end else if (start_reg_89) begin // @[SWChisel.scala 207:25]
      E_89 <= array_89_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_90 <= -16'sh5c; // @[SWChisel.scala 162:18]
    end else if (start_reg_90) begin // @[SWChisel.scala 207:25]
      E_90 <= array_90_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_91 <= -16'sh5d; // @[SWChisel.scala 162:18]
    end else if (start_reg_91) begin // @[SWChisel.scala 207:25]
      E_91 <= array_91_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_92 <= -16'sh5e; // @[SWChisel.scala 162:18]
    end else if (start_reg_92) begin // @[SWChisel.scala 207:25]
      E_92 <= array_92_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_93 <= -16'sh5f; // @[SWChisel.scala 162:18]
    end else if (start_reg_93) begin // @[SWChisel.scala 207:25]
      E_93 <= array_93_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_94 <= -16'sh60; // @[SWChisel.scala 162:18]
    end else if (start_reg_94) begin // @[SWChisel.scala 207:25]
      E_94 <= array_94_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_95 <= -16'sh61; // @[SWChisel.scala 162:18]
    end else if (start_reg_95) begin // @[SWChisel.scala 207:25]
      E_95 <= array_95_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_96 <= -16'sh62; // @[SWChisel.scala 162:18]
    end else if (start_reg_96) begin // @[SWChisel.scala 207:25]
      E_96 <= array_96_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_97 <= -16'sh63; // @[SWChisel.scala 162:18]
    end else if (start_reg_97) begin // @[SWChisel.scala 207:25]
      E_97 <= array_97_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_98 <= -16'sh64; // @[SWChisel.scala 162:18]
    end else if (start_reg_98) begin // @[SWChisel.scala 207:25]
      E_98 <= array_98_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_99 <= -16'sh65; // @[SWChisel.scala 162:18]
    end else if (start_reg_99) begin // @[SWChisel.scala 207:25]
      E_99 <= array_99_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_1 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      F_1 <= array_0_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_2 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      F_2 <= array_1_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_3 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      F_3 <= array_2_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_4 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      F_4 <= array_3_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_5 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      F_5 <= array_4_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_6 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      F_6 <= array_5_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_7 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      F_7 <= array_6_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_8 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      F_8 <= array_7_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_9 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      F_9 <= array_8_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_10 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      F_10 <= array_9_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_11 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      F_11 <= array_10_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_12 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      F_12 <= array_11_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_13 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      F_13 <= array_12_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_14 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      F_14 <= array_13_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_15 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      F_15 <= array_14_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_16 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      F_16 <= array_15_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_17 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      F_17 <= array_16_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_18 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      F_18 <= array_17_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_19 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      F_19 <= array_18_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_20 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      F_20 <= array_19_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_21 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      F_21 <= array_20_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_22 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      F_22 <= array_21_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_23 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      F_23 <= array_22_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_24 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      F_24 <= array_23_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_25 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      F_25 <= array_24_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_26 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      F_26 <= array_25_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_27 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      F_27 <= array_26_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_28 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      F_28 <= array_27_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_29 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      F_29 <= array_28_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_30 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_29) begin // @[SWChisel.scala 207:25]
      F_30 <= array_29_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_31 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_30) begin // @[SWChisel.scala 207:25]
      F_31 <= array_30_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_32 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_31) begin // @[SWChisel.scala 207:25]
      F_32 <= array_31_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_33 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_32) begin // @[SWChisel.scala 207:25]
      F_33 <= array_32_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_34 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_33) begin // @[SWChisel.scala 207:25]
      F_34 <= array_33_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_35 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_34) begin // @[SWChisel.scala 207:25]
      F_35 <= array_34_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_36 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_35) begin // @[SWChisel.scala 207:25]
      F_36 <= array_35_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_37 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_36) begin // @[SWChisel.scala 207:25]
      F_37 <= array_36_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_38 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_37) begin // @[SWChisel.scala 207:25]
      F_38 <= array_37_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_39 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_38) begin // @[SWChisel.scala 207:25]
      F_39 <= array_38_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_40 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_39) begin // @[SWChisel.scala 207:25]
      F_40 <= array_39_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_41 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_40) begin // @[SWChisel.scala 207:25]
      F_41 <= array_40_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_42 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_41) begin // @[SWChisel.scala 207:25]
      F_42 <= array_41_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_43 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_42) begin // @[SWChisel.scala 207:25]
      F_43 <= array_42_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_44 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_43) begin // @[SWChisel.scala 207:25]
      F_44 <= array_43_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_45 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_44) begin // @[SWChisel.scala 207:25]
      F_45 <= array_44_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_46 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_45) begin // @[SWChisel.scala 207:25]
      F_46 <= array_45_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_47 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_46) begin // @[SWChisel.scala 207:25]
      F_47 <= array_46_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_48 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_47) begin // @[SWChisel.scala 207:25]
      F_48 <= array_47_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_49 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_48) begin // @[SWChisel.scala 207:25]
      F_49 <= array_48_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_50 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_49) begin // @[SWChisel.scala 207:25]
      F_50 <= array_49_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_51 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_50) begin // @[SWChisel.scala 207:25]
      F_51 <= array_50_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_52 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_51) begin // @[SWChisel.scala 207:25]
      F_52 <= array_51_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_53 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_52) begin // @[SWChisel.scala 207:25]
      F_53 <= array_52_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_54 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_53) begin // @[SWChisel.scala 207:25]
      F_54 <= array_53_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_55 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_54) begin // @[SWChisel.scala 207:25]
      F_55 <= array_54_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_56 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_55) begin // @[SWChisel.scala 207:25]
      F_56 <= array_55_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_57 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_56) begin // @[SWChisel.scala 207:25]
      F_57 <= array_56_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_58 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_57) begin // @[SWChisel.scala 207:25]
      F_58 <= array_57_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_59 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_58) begin // @[SWChisel.scala 207:25]
      F_59 <= array_58_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_60 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_59) begin // @[SWChisel.scala 207:25]
      F_60 <= array_59_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_61 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_60) begin // @[SWChisel.scala 207:25]
      F_61 <= array_60_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_62 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_61) begin // @[SWChisel.scala 207:25]
      F_62 <= array_61_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_63 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_62) begin // @[SWChisel.scala 207:25]
      F_63 <= array_62_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_64 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_63) begin // @[SWChisel.scala 207:25]
      F_64 <= array_63_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_65 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_64) begin // @[SWChisel.scala 207:25]
      F_65 <= array_64_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_66 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_65) begin // @[SWChisel.scala 207:25]
      F_66 <= array_65_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_67 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_66) begin // @[SWChisel.scala 207:25]
      F_67 <= array_66_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_68 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_67) begin // @[SWChisel.scala 207:25]
      F_68 <= array_67_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_69 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_68) begin // @[SWChisel.scala 207:25]
      F_69 <= array_68_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_70 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_69) begin // @[SWChisel.scala 207:25]
      F_70 <= array_69_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_71 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_70) begin // @[SWChisel.scala 207:25]
      F_71 <= array_70_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_72 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_71) begin // @[SWChisel.scala 207:25]
      F_72 <= array_71_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_73 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_72) begin // @[SWChisel.scala 207:25]
      F_73 <= array_72_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_74 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_73) begin // @[SWChisel.scala 207:25]
      F_74 <= array_73_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_75 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_74) begin // @[SWChisel.scala 207:25]
      F_75 <= array_74_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_76 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_75) begin // @[SWChisel.scala 207:25]
      F_76 <= array_75_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_77 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_76) begin // @[SWChisel.scala 207:25]
      F_77 <= array_76_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_78 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_77) begin // @[SWChisel.scala 207:25]
      F_78 <= array_77_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_79 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_78) begin // @[SWChisel.scala 207:25]
      F_79 <= array_78_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_80 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_79) begin // @[SWChisel.scala 207:25]
      F_80 <= array_79_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_81 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_80) begin // @[SWChisel.scala 207:25]
      F_81 <= array_80_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_82 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_81) begin // @[SWChisel.scala 207:25]
      F_82 <= array_81_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_83 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_82) begin // @[SWChisel.scala 207:25]
      F_83 <= array_82_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_84 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_83) begin // @[SWChisel.scala 207:25]
      F_84 <= array_83_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_85 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_84) begin // @[SWChisel.scala 207:25]
      F_85 <= array_84_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_86 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_85) begin // @[SWChisel.scala 207:25]
      F_86 <= array_85_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_87 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_86) begin // @[SWChisel.scala 207:25]
      F_87 <= array_86_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_88 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_87) begin // @[SWChisel.scala 207:25]
      F_88 <= array_87_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_89 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_88) begin // @[SWChisel.scala 207:25]
      F_89 <= array_88_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_90 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_89) begin // @[SWChisel.scala 207:25]
      F_90 <= array_89_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_91 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_90) begin // @[SWChisel.scala 207:25]
      F_91 <= array_90_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_92 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_91) begin // @[SWChisel.scala 207:25]
      F_92 <= array_91_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_93 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_92) begin // @[SWChisel.scala 207:25]
      F_93 <= array_92_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_94 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_93) begin // @[SWChisel.scala 207:25]
      F_94 <= array_93_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_95 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_94) begin // @[SWChisel.scala 207:25]
      F_95 <= array_94_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_96 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_95) begin // @[SWChisel.scala 207:25]
      F_96 <= array_95_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_97 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_96) begin // @[SWChisel.scala 207:25]
      F_97 <= array_96_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_98 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_97) begin // @[SWChisel.scala 207:25]
      F_98 <= array_97_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_99 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_98) begin // @[SWChisel.scala 207:25]
      F_99 <= array_98_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_0 <= -16'sh1; // @[SWChisel.scala 164:19]
    end else begin
      V1_0 <= 16'sh0; // @[SWChisel.scala 165:9]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_1 <= -16'sh2; // @[SWChisel.scala 164:19]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      V1_1 <= array_0_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_2 <= -16'sh3; // @[SWChisel.scala 164:19]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      V1_2 <= array_1_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_3 <= -16'sh4; // @[SWChisel.scala 164:19]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      V1_3 <= array_2_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_4 <= -16'sh5; // @[SWChisel.scala 164:19]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      V1_4 <= array_3_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_5 <= -16'sh6; // @[SWChisel.scala 164:19]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      V1_5 <= array_4_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_6 <= -16'sh7; // @[SWChisel.scala 164:19]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      V1_6 <= array_5_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_7 <= -16'sh8; // @[SWChisel.scala 164:19]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      V1_7 <= array_6_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_8 <= -16'sh9; // @[SWChisel.scala 164:19]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      V1_8 <= array_7_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_9 <= -16'sha; // @[SWChisel.scala 164:19]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      V1_9 <= array_8_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_10 <= -16'shb; // @[SWChisel.scala 164:19]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      V1_10 <= array_9_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_11 <= -16'shc; // @[SWChisel.scala 164:19]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      V1_11 <= array_10_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_12 <= -16'shd; // @[SWChisel.scala 164:19]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      V1_12 <= array_11_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_13 <= -16'she; // @[SWChisel.scala 164:19]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      V1_13 <= array_12_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_14 <= -16'shf; // @[SWChisel.scala 164:19]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      V1_14 <= array_13_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_15 <= -16'sh10; // @[SWChisel.scala 164:19]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      V1_15 <= array_14_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_16 <= -16'sh11; // @[SWChisel.scala 164:19]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      V1_16 <= array_15_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_17 <= -16'sh12; // @[SWChisel.scala 164:19]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      V1_17 <= array_16_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_18 <= -16'sh13; // @[SWChisel.scala 164:19]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      V1_18 <= array_17_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_19 <= -16'sh14; // @[SWChisel.scala 164:19]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      V1_19 <= array_18_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_20 <= -16'sh15; // @[SWChisel.scala 164:19]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      V1_20 <= array_19_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_21 <= -16'sh16; // @[SWChisel.scala 164:19]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      V1_21 <= array_20_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_22 <= -16'sh17; // @[SWChisel.scala 164:19]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      V1_22 <= array_21_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_23 <= -16'sh18; // @[SWChisel.scala 164:19]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      V1_23 <= array_22_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_24 <= -16'sh19; // @[SWChisel.scala 164:19]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      V1_24 <= array_23_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_25 <= -16'sh1a; // @[SWChisel.scala 164:19]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      V1_25 <= array_24_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_26 <= -16'sh1b; // @[SWChisel.scala 164:19]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      V1_26 <= array_25_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_27 <= -16'sh1c; // @[SWChisel.scala 164:19]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      V1_27 <= array_26_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_28 <= -16'sh1d; // @[SWChisel.scala 164:19]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      V1_28 <= array_27_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_29 <= -16'sh1e; // @[SWChisel.scala 164:19]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      V1_29 <= array_28_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_30 <= -16'sh1f; // @[SWChisel.scala 164:19]
    end else if (start_reg_29) begin // @[SWChisel.scala 207:25]
      V1_30 <= array_29_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_31 <= -16'sh20; // @[SWChisel.scala 164:19]
    end else if (start_reg_30) begin // @[SWChisel.scala 207:25]
      V1_31 <= array_30_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_32 <= -16'sh21; // @[SWChisel.scala 164:19]
    end else if (start_reg_31) begin // @[SWChisel.scala 207:25]
      V1_32 <= array_31_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_33 <= -16'sh22; // @[SWChisel.scala 164:19]
    end else if (start_reg_32) begin // @[SWChisel.scala 207:25]
      V1_33 <= array_32_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_34 <= -16'sh23; // @[SWChisel.scala 164:19]
    end else if (start_reg_33) begin // @[SWChisel.scala 207:25]
      V1_34 <= array_33_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_35 <= -16'sh24; // @[SWChisel.scala 164:19]
    end else if (start_reg_34) begin // @[SWChisel.scala 207:25]
      V1_35 <= array_34_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_36 <= -16'sh25; // @[SWChisel.scala 164:19]
    end else if (start_reg_35) begin // @[SWChisel.scala 207:25]
      V1_36 <= array_35_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_37 <= -16'sh26; // @[SWChisel.scala 164:19]
    end else if (start_reg_36) begin // @[SWChisel.scala 207:25]
      V1_37 <= array_36_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_38 <= -16'sh27; // @[SWChisel.scala 164:19]
    end else if (start_reg_37) begin // @[SWChisel.scala 207:25]
      V1_38 <= array_37_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_39 <= -16'sh28; // @[SWChisel.scala 164:19]
    end else if (start_reg_38) begin // @[SWChisel.scala 207:25]
      V1_39 <= array_38_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_40 <= -16'sh29; // @[SWChisel.scala 164:19]
    end else if (start_reg_39) begin // @[SWChisel.scala 207:25]
      V1_40 <= array_39_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_41 <= -16'sh2a; // @[SWChisel.scala 164:19]
    end else if (start_reg_40) begin // @[SWChisel.scala 207:25]
      V1_41 <= array_40_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_42 <= -16'sh2b; // @[SWChisel.scala 164:19]
    end else if (start_reg_41) begin // @[SWChisel.scala 207:25]
      V1_42 <= array_41_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_43 <= -16'sh2c; // @[SWChisel.scala 164:19]
    end else if (start_reg_42) begin // @[SWChisel.scala 207:25]
      V1_43 <= array_42_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_44 <= -16'sh2d; // @[SWChisel.scala 164:19]
    end else if (start_reg_43) begin // @[SWChisel.scala 207:25]
      V1_44 <= array_43_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_45 <= -16'sh2e; // @[SWChisel.scala 164:19]
    end else if (start_reg_44) begin // @[SWChisel.scala 207:25]
      V1_45 <= array_44_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_46 <= -16'sh2f; // @[SWChisel.scala 164:19]
    end else if (start_reg_45) begin // @[SWChisel.scala 207:25]
      V1_46 <= array_45_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_47 <= -16'sh30; // @[SWChisel.scala 164:19]
    end else if (start_reg_46) begin // @[SWChisel.scala 207:25]
      V1_47 <= array_46_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_48 <= -16'sh31; // @[SWChisel.scala 164:19]
    end else if (start_reg_47) begin // @[SWChisel.scala 207:25]
      V1_48 <= array_47_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_49 <= -16'sh32; // @[SWChisel.scala 164:19]
    end else if (start_reg_48) begin // @[SWChisel.scala 207:25]
      V1_49 <= array_48_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_50 <= -16'sh33; // @[SWChisel.scala 164:19]
    end else if (start_reg_49) begin // @[SWChisel.scala 207:25]
      V1_50 <= array_49_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_51 <= -16'sh34; // @[SWChisel.scala 164:19]
    end else if (start_reg_50) begin // @[SWChisel.scala 207:25]
      V1_51 <= array_50_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_52 <= -16'sh35; // @[SWChisel.scala 164:19]
    end else if (start_reg_51) begin // @[SWChisel.scala 207:25]
      V1_52 <= array_51_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_53 <= -16'sh36; // @[SWChisel.scala 164:19]
    end else if (start_reg_52) begin // @[SWChisel.scala 207:25]
      V1_53 <= array_52_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_54 <= -16'sh37; // @[SWChisel.scala 164:19]
    end else if (start_reg_53) begin // @[SWChisel.scala 207:25]
      V1_54 <= array_53_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_55 <= -16'sh38; // @[SWChisel.scala 164:19]
    end else if (start_reg_54) begin // @[SWChisel.scala 207:25]
      V1_55 <= array_54_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_56 <= -16'sh39; // @[SWChisel.scala 164:19]
    end else if (start_reg_55) begin // @[SWChisel.scala 207:25]
      V1_56 <= array_55_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_57 <= -16'sh3a; // @[SWChisel.scala 164:19]
    end else if (start_reg_56) begin // @[SWChisel.scala 207:25]
      V1_57 <= array_56_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_58 <= -16'sh3b; // @[SWChisel.scala 164:19]
    end else if (start_reg_57) begin // @[SWChisel.scala 207:25]
      V1_58 <= array_57_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_59 <= -16'sh3c; // @[SWChisel.scala 164:19]
    end else if (start_reg_58) begin // @[SWChisel.scala 207:25]
      V1_59 <= array_58_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_60 <= -16'sh3d; // @[SWChisel.scala 164:19]
    end else if (start_reg_59) begin // @[SWChisel.scala 207:25]
      V1_60 <= array_59_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_61 <= -16'sh3e; // @[SWChisel.scala 164:19]
    end else if (start_reg_60) begin // @[SWChisel.scala 207:25]
      V1_61 <= array_60_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_62 <= -16'sh3f; // @[SWChisel.scala 164:19]
    end else if (start_reg_61) begin // @[SWChisel.scala 207:25]
      V1_62 <= array_61_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_63 <= -16'sh40; // @[SWChisel.scala 164:19]
    end else if (start_reg_62) begin // @[SWChisel.scala 207:25]
      V1_63 <= array_62_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_64 <= -16'sh41; // @[SWChisel.scala 164:19]
    end else if (start_reg_63) begin // @[SWChisel.scala 207:25]
      V1_64 <= array_63_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_65 <= -16'sh42; // @[SWChisel.scala 164:19]
    end else if (start_reg_64) begin // @[SWChisel.scala 207:25]
      V1_65 <= array_64_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_66 <= -16'sh43; // @[SWChisel.scala 164:19]
    end else if (start_reg_65) begin // @[SWChisel.scala 207:25]
      V1_66 <= array_65_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_67 <= -16'sh44; // @[SWChisel.scala 164:19]
    end else if (start_reg_66) begin // @[SWChisel.scala 207:25]
      V1_67 <= array_66_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_68 <= -16'sh45; // @[SWChisel.scala 164:19]
    end else if (start_reg_67) begin // @[SWChisel.scala 207:25]
      V1_68 <= array_67_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_69 <= -16'sh46; // @[SWChisel.scala 164:19]
    end else if (start_reg_68) begin // @[SWChisel.scala 207:25]
      V1_69 <= array_68_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_70 <= -16'sh47; // @[SWChisel.scala 164:19]
    end else if (start_reg_69) begin // @[SWChisel.scala 207:25]
      V1_70 <= array_69_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_71 <= -16'sh48; // @[SWChisel.scala 164:19]
    end else if (start_reg_70) begin // @[SWChisel.scala 207:25]
      V1_71 <= array_70_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_72 <= -16'sh49; // @[SWChisel.scala 164:19]
    end else if (start_reg_71) begin // @[SWChisel.scala 207:25]
      V1_72 <= array_71_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_73 <= -16'sh4a; // @[SWChisel.scala 164:19]
    end else if (start_reg_72) begin // @[SWChisel.scala 207:25]
      V1_73 <= array_72_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_74 <= -16'sh4b; // @[SWChisel.scala 164:19]
    end else if (start_reg_73) begin // @[SWChisel.scala 207:25]
      V1_74 <= array_73_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_75 <= -16'sh4c; // @[SWChisel.scala 164:19]
    end else if (start_reg_74) begin // @[SWChisel.scala 207:25]
      V1_75 <= array_74_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_76 <= -16'sh4d; // @[SWChisel.scala 164:19]
    end else if (start_reg_75) begin // @[SWChisel.scala 207:25]
      V1_76 <= array_75_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_77 <= -16'sh4e; // @[SWChisel.scala 164:19]
    end else if (start_reg_76) begin // @[SWChisel.scala 207:25]
      V1_77 <= array_76_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_78 <= -16'sh4f; // @[SWChisel.scala 164:19]
    end else if (start_reg_77) begin // @[SWChisel.scala 207:25]
      V1_78 <= array_77_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_79 <= -16'sh50; // @[SWChisel.scala 164:19]
    end else if (start_reg_78) begin // @[SWChisel.scala 207:25]
      V1_79 <= array_78_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_80 <= -16'sh51; // @[SWChisel.scala 164:19]
    end else if (start_reg_79) begin // @[SWChisel.scala 207:25]
      V1_80 <= array_79_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_81 <= -16'sh52; // @[SWChisel.scala 164:19]
    end else if (start_reg_80) begin // @[SWChisel.scala 207:25]
      V1_81 <= array_80_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_82 <= -16'sh53; // @[SWChisel.scala 164:19]
    end else if (start_reg_81) begin // @[SWChisel.scala 207:25]
      V1_82 <= array_81_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_83 <= -16'sh54; // @[SWChisel.scala 164:19]
    end else if (start_reg_82) begin // @[SWChisel.scala 207:25]
      V1_83 <= array_82_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_84 <= -16'sh55; // @[SWChisel.scala 164:19]
    end else if (start_reg_83) begin // @[SWChisel.scala 207:25]
      V1_84 <= array_83_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_85 <= -16'sh56; // @[SWChisel.scala 164:19]
    end else if (start_reg_84) begin // @[SWChisel.scala 207:25]
      V1_85 <= array_84_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_86 <= -16'sh57; // @[SWChisel.scala 164:19]
    end else if (start_reg_85) begin // @[SWChisel.scala 207:25]
      V1_86 <= array_85_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_87 <= -16'sh58; // @[SWChisel.scala 164:19]
    end else if (start_reg_86) begin // @[SWChisel.scala 207:25]
      V1_87 <= array_86_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_88 <= -16'sh59; // @[SWChisel.scala 164:19]
    end else if (start_reg_87) begin // @[SWChisel.scala 207:25]
      V1_88 <= array_87_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_89 <= -16'sh5a; // @[SWChisel.scala 164:19]
    end else if (start_reg_88) begin // @[SWChisel.scala 207:25]
      V1_89 <= array_88_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_90 <= -16'sh5b; // @[SWChisel.scala 164:19]
    end else if (start_reg_89) begin // @[SWChisel.scala 207:25]
      V1_90 <= array_89_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_91 <= -16'sh5c; // @[SWChisel.scala 164:19]
    end else if (start_reg_90) begin // @[SWChisel.scala 207:25]
      V1_91 <= array_90_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_92 <= -16'sh5d; // @[SWChisel.scala 164:19]
    end else if (start_reg_91) begin // @[SWChisel.scala 207:25]
      V1_92 <= array_91_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_93 <= -16'sh5e; // @[SWChisel.scala 164:19]
    end else if (start_reg_92) begin // @[SWChisel.scala 207:25]
      V1_93 <= array_92_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_94 <= -16'sh5f; // @[SWChisel.scala 164:19]
    end else if (start_reg_93) begin // @[SWChisel.scala 207:25]
      V1_94 <= array_93_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_95 <= -16'sh60; // @[SWChisel.scala 164:19]
    end else if (start_reg_94) begin // @[SWChisel.scala 207:25]
      V1_95 <= array_94_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_96 <= -16'sh61; // @[SWChisel.scala 164:19]
    end else if (start_reg_95) begin // @[SWChisel.scala 207:25]
      V1_96 <= array_95_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_97 <= -16'sh62; // @[SWChisel.scala 164:19]
    end else if (start_reg_96) begin // @[SWChisel.scala 207:25]
      V1_97 <= array_96_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_98 <= -16'sh63; // @[SWChisel.scala 164:19]
    end else if (start_reg_97) begin // @[SWChisel.scala 207:25]
      V1_98 <= array_97_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_99 <= -16'sh64; // @[SWChisel.scala 164:19]
    end else if (start_reg_98) begin // @[SWChisel.scala 207:25]
      V1_99 <= array_98_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_100 <= -16'sh65; // @[SWChisel.scala 164:19]
    end else if (start_reg_99) begin // @[SWChisel.scala 207:25]
      V1_100 <= array_99_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_0 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_0 <= V1_0; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_1 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_1 <= V1_1; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_2 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_2 <= V1_2; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_3 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_3 <= V1_3; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_4 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_4 <= V1_4; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_5 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_5 <= V1_5; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_6 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_6 <= V1_6; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_7 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_7 <= V1_7; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_8 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_8 <= V1_8; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_9 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_9 <= V1_9; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_10 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_10 <= V1_10; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_11 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_11 <= V1_11; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_12 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_12 <= V1_12; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_13 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_13 <= V1_13; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_14 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_14 <= V1_14; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_15 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_15 <= V1_15; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_16 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_16 <= V1_16; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_17 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_17 <= V1_17; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_18 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_18 <= V1_18; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_19 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_19 <= V1_19; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_20 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_20 <= V1_20; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_21 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_21 <= V1_21; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_22 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_22 <= V1_22; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_23 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_23 <= V1_23; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_24 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_24 <= V1_24; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_25 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_25 <= V1_25; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_26 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_26 <= V1_26; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_27 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_27 <= V1_27; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_28 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_28 <= V1_28; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_29 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_29 <= V1_29; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_30 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_30 <= V1_30; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_31 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_31 <= V1_31; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_32 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_32 <= V1_32; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_33 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_33 <= V1_33; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_34 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_34 <= V1_34; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_35 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_35 <= V1_35; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_36 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_36 <= V1_36; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_37 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_37 <= V1_37; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_38 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_38 <= V1_38; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_39 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_39 <= V1_39; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_40 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_40 <= V1_40; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_41 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_41 <= V1_41; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_42 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_42 <= V1_42; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_43 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_43 <= V1_43; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_44 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_44 <= V1_44; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_45 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_45 <= V1_45; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_46 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_46 <= V1_46; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_47 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_47 <= V1_47; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_48 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_48 <= V1_48; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_49 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_49 <= V1_49; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_50 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_50 <= V1_50; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_51 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_51 <= V1_51; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_52 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_52 <= V1_52; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_53 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_53 <= V1_53; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_54 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_54 <= V1_54; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_55 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_55 <= V1_55; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_56 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_56 <= V1_56; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_57 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_57 <= V1_57; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_58 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_58 <= V1_58; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_59 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_59 <= V1_59; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_60 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_60 <= V1_60; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_61 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_61 <= V1_61; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_62 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_62 <= V1_62; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_63 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_63 <= V1_63; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_64 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_64 <= V1_64; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_65 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_65 <= V1_65; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_66 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_66 <= V1_66; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_67 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_67 <= V1_67; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_68 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_68 <= V1_68; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_69 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_69 <= V1_69; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_70 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_70 <= V1_70; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_71 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_71 <= V1_71; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_72 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_72 <= V1_72; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_73 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_73 <= V1_73; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_74 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_74 <= V1_74; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_75 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_75 <= V1_75; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_76 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_76 <= V1_76; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_77 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_77 <= V1_77; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_78 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_78 <= V1_78; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_79 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_79 <= V1_79; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_80 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_80 <= V1_80; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_81 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_81 <= V1_81; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_82 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_82 <= V1_82; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_83 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_83 <= V1_83; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_84 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_84 <= V1_84; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_85 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_85 <= V1_85; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_86 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_86 <= V1_86; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_87 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_87 <= V1_87; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_88 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_88 <= V1_88; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_89 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_89 <= V1_89; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_90 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_90 <= V1_90; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_91 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_91 <= V1_91; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_92 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_92 <= V1_92; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_93 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_93 <= V1_93; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_94 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_94 <= V1_94; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_95 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_95 <= V1_95; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_96 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_96 <= V1_96; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_97 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_97 <= V1_97; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_98 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_98 <= V1_98; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_99 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_99 <= V1_99; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_0 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_0 <= io_start; // @[SWChisel.scala 185:16]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_1 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_1 <= start_reg_0; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_2 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_2 <= start_reg_1; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_3 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_3 <= start_reg_2; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_4 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_4 <= start_reg_3; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_5 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_5 <= start_reg_4; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_6 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_6 <= start_reg_5; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_7 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_7 <= start_reg_6; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_8 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_8 <= start_reg_7; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_9 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_9 <= start_reg_8; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_10 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_10 <= start_reg_9; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_11 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_11 <= start_reg_10; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_12 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_12 <= start_reg_11; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_13 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_13 <= start_reg_12; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_14 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_14 <= start_reg_13; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_15 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_15 <= start_reg_14; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_16 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_16 <= start_reg_15; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_17 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_17 <= start_reg_16; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_18 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_18 <= start_reg_17; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_19 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_19 <= start_reg_18; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_20 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_20 <= start_reg_19; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_21 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_21 <= start_reg_20; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_22 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_22 <= start_reg_21; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_23 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_23 <= start_reg_22; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_24 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_24 <= start_reg_23; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_25 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_25 <= start_reg_24; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_26 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_26 <= start_reg_25; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_27 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_27 <= start_reg_26; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_28 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_28 <= start_reg_27; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_29 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_29 <= start_reg_28; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_30 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_30 <= start_reg_29; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_31 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_31 <= start_reg_30; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_32 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_32 <= start_reg_31; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_33 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_33 <= start_reg_32; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_34 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_34 <= start_reg_33; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_35 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_35 <= start_reg_34; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_36 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_36 <= start_reg_35; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_37 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_37 <= start_reg_36; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_38 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_38 <= start_reg_37; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_39 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_39 <= start_reg_38; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_40 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_40 <= start_reg_39; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_41 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_41 <= start_reg_40; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_42 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_42 <= start_reg_41; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_43 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_43 <= start_reg_42; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_44 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_44 <= start_reg_43; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_45 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_45 <= start_reg_44; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_46 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_46 <= start_reg_45; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_47 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_47 <= start_reg_46; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_48 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_48 <= start_reg_47; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_49 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_49 <= start_reg_48; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_50 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_50 <= start_reg_49; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_51 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_51 <= start_reg_50; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_52 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_52 <= start_reg_51; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_53 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_53 <= start_reg_52; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_54 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_54 <= start_reg_53; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_55 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_55 <= start_reg_54; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_56 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_56 <= start_reg_55; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_57 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_57 <= start_reg_56; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_58 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_58 <= start_reg_57; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_59 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_59 <= start_reg_58; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_60 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_60 <= start_reg_59; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_61 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_61 <= start_reg_60; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_62 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_62 <= start_reg_61; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_63 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_63 <= start_reg_62; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_64 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_64 <= start_reg_63; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_65 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_65 <= start_reg_64; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_66 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_66 <= start_reg_65; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_67 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_67 <= start_reg_66; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_68 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_68 <= start_reg_67; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_69 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_69 <= start_reg_68; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_70 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_70 <= start_reg_69; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_71 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_71 <= start_reg_70; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_72 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_72 <= start_reg_71; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_73 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_73 <= start_reg_72; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_74 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_74 <= start_reg_73; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_75 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_75 <= start_reg_74; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_76 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_76 <= start_reg_75; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_77 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_77 <= start_reg_76; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_78 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_78 <= start_reg_77; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_79 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_79 <= start_reg_78; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_80 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_80 <= start_reg_79; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_81 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_81 <= start_reg_80; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_82 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_82 <= start_reg_81; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_83 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_83 <= start_reg_82; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_84 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_84 <= start_reg_83; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_85 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_85 <= start_reg_84; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_86 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_86 <= start_reg_85; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_87 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_87 <= start_reg_86; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_88 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_88 <= start_reg_87; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_89 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_89 <= start_reg_88; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_90 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_90 <= start_reg_89; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_91 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_91 <= start_reg_90; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_92 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_92 <= start_reg_91; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_93 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_93 <= start_reg_92; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_94 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_94 <= start_reg_93; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_95 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_95 <= start_reg_94; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_96 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_96 <= start_reg_95; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_97 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_97 <= start_reg_96; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_98 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_98 <= start_reg_97; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_99 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_99 <= start_reg_98; // @[SWChisel.scala 187:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  E_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  E_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  E_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  E_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  E_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  E_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  E_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  E_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  E_8 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  E_9 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  E_10 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  E_11 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  E_12 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  E_13 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  E_14 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  E_15 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  E_16 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  E_17 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  E_18 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  E_19 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  E_20 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  E_21 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  E_22 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  E_23 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  E_24 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  E_25 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  E_26 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  E_27 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  E_28 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  E_29 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  E_30 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  E_31 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  E_32 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  E_33 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  E_34 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  E_35 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  E_36 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  E_37 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  E_38 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  E_39 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  E_40 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  E_41 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  E_42 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  E_43 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  E_44 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  E_45 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  E_46 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  E_47 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  E_48 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  E_49 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  E_50 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  E_51 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  E_52 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  E_53 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  E_54 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  E_55 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  E_56 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  E_57 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  E_58 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  E_59 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  E_60 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  E_61 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  E_62 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  E_63 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  E_64 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  E_65 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  E_66 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  E_67 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  E_68 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  E_69 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  E_70 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  E_71 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  E_72 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  E_73 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  E_74 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  E_75 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  E_76 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  E_77 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  E_78 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  E_79 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  E_80 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  E_81 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  E_82 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  E_83 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  E_84 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  E_85 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  E_86 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  E_87 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  E_88 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  E_89 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  E_90 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  E_91 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  E_92 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  E_93 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  E_94 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  E_95 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  E_96 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  E_97 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  E_98 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  E_99 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  F_1 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  F_2 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  F_3 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  F_4 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  F_5 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  F_6 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  F_7 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  F_8 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  F_9 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  F_10 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  F_11 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  F_12 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  F_13 = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  F_14 = _RAND_113[15:0];
  _RAND_114 = {1{`RANDOM}};
  F_15 = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  F_16 = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  F_17 = _RAND_116[15:0];
  _RAND_117 = {1{`RANDOM}};
  F_18 = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  F_19 = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  F_20 = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  F_21 = _RAND_120[15:0];
  _RAND_121 = {1{`RANDOM}};
  F_22 = _RAND_121[15:0];
  _RAND_122 = {1{`RANDOM}};
  F_23 = _RAND_122[15:0];
  _RAND_123 = {1{`RANDOM}};
  F_24 = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  F_25 = _RAND_124[15:0];
  _RAND_125 = {1{`RANDOM}};
  F_26 = _RAND_125[15:0];
  _RAND_126 = {1{`RANDOM}};
  F_27 = _RAND_126[15:0];
  _RAND_127 = {1{`RANDOM}};
  F_28 = _RAND_127[15:0];
  _RAND_128 = {1{`RANDOM}};
  F_29 = _RAND_128[15:0];
  _RAND_129 = {1{`RANDOM}};
  F_30 = _RAND_129[15:0];
  _RAND_130 = {1{`RANDOM}};
  F_31 = _RAND_130[15:0];
  _RAND_131 = {1{`RANDOM}};
  F_32 = _RAND_131[15:0];
  _RAND_132 = {1{`RANDOM}};
  F_33 = _RAND_132[15:0];
  _RAND_133 = {1{`RANDOM}};
  F_34 = _RAND_133[15:0];
  _RAND_134 = {1{`RANDOM}};
  F_35 = _RAND_134[15:0];
  _RAND_135 = {1{`RANDOM}};
  F_36 = _RAND_135[15:0];
  _RAND_136 = {1{`RANDOM}};
  F_37 = _RAND_136[15:0];
  _RAND_137 = {1{`RANDOM}};
  F_38 = _RAND_137[15:0];
  _RAND_138 = {1{`RANDOM}};
  F_39 = _RAND_138[15:0];
  _RAND_139 = {1{`RANDOM}};
  F_40 = _RAND_139[15:0];
  _RAND_140 = {1{`RANDOM}};
  F_41 = _RAND_140[15:0];
  _RAND_141 = {1{`RANDOM}};
  F_42 = _RAND_141[15:0];
  _RAND_142 = {1{`RANDOM}};
  F_43 = _RAND_142[15:0];
  _RAND_143 = {1{`RANDOM}};
  F_44 = _RAND_143[15:0];
  _RAND_144 = {1{`RANDOM}};
  F_45 = _RAND_144[15:0];
  _RAND_145 = {1{`RANDOM}};
  F_46 = _RAND_145[15:0];
  _RAND_146 = {1{`RANDOM}};
  F_47 = _RAND_146[15:0];
  _RAND_147 = {1{`RANDOM}};
  F_48 = _RAND_147[15:0];
  _RAND_148 = {1{`RANDOM}};
  F_49 = _RAND_148[15:0];
  _RAND_149 = {1{`RANDOM}};
  F_50 = _RAND_149[15:0];
  _RAND_150 = {1{`RANDOM}};
  F_51 = _RAND_150[15:0];
  _RAND_151 = {1{`RANDOM}};
  F_52 = _RAND_151[15:0];
  _RAND_152 = {1{`RANDOM}};
  F_53 = _RAND_152[15:0];
  _RAND_153 = {1{`RANDOM}};
  F_54 = _RAND_153[15:0];
  _RAND_154 = {1{`RANDOM}};
  F_55 = _RAND_154[15:0];
  _RAND_155 = {1{`RANDOM}};
  F_56 = _RAND_155[15:0];
  _RAND_156 = {1{`RANDOM}};
  F_57 = _RAND_156[15:0];
  _RAND_157 = {1{`RANDOM}};
  F_58 = _RAND_157[15:0];
  _RAND_158 = {1{`RANDOM}};
  F_59 = _RAND_158[15:0];
  _RAND_159 = {1{`RANDOM}};
  F_60 = _RAND_159[15:0];
  _RAND_160 = {1{`RANDOM}};
  F_61 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  F_62 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  F_63 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  F_64 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  F_65 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  F_66 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  F_67 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  F_68 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  F_69 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  F_70 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  F_71 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  F_72 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  F_73 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  F_74 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  F_75 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  F_76 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  F_77 = _RAND_176[15:0];
  _RAND_177 = {1{`RANDOM}};
  F_78 = _RAND_177[15:0];
  _RAND_178 = {1{`RANDOM}};
  F_79 = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  F_80 = _RAND_179[15:0];
  _RAND_180 = {1{`RANDOM}};
  F_81 = _RAND_180[15:0];
  _RAND_181 = {1{`RANDOM}};
  F_82 = _RAND_181[15:0];
  _RAND_182 = {1{`RANDOM}};
  F_83 = _RAND_182[15:0];
  _RAND_183 = {1{`RANDOM}};
  F_84 = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  F_85 = _RAND_184[15:0];
  _RAND_185 = {1{`RANDOM}};
  F_86 = _RAND_185[15:0];
  _RAND_186 = {1{`RANDOM}};
  F_87 = _RAND_186[15:0];
  _RAND_187 = {1{`RANDOM}};
  F_88 = _RAND_187[15:0];
  _RAND_188 = {1{`RANDOM}};
  F_89 = _RAND_188[15:0];
  _RAND_189 = {1{`RANDOM}};
  F_90 = _RAND_189[15:0];
  _RAND_190 = {1{`RANDOM}};
  F_91 = _RAND_190[15:0];
  _RAND_191 = {1{`RANDOM}};
  F_92 = _RAND_191[15:0];
  _RAND_192 = {1{`RANDOM}};
  F_93 = _RAND_192[15:0];
  _RAND_193 = {1{`RANDOM}};
  F_94 = _RAND_193[15:0];
  _RAND_194 = {1{`RANDOM}};
  F_95 = _RAND_194[15:0];
  _RAND_195 = {1{`RANDOM}};
  F_96 = _RAND_195[15:0];
  _RAND_196 = {1{`RANDOM}};
  F_97 = _RAND_196[15:0];
  _RAND_197 = {1{`RANDOM}};
  F_98 = _RAND_197[15:0];
  _RAND_198 = {1{`RANDOM}};
  F_99 = _RAND_198[15:0];
  _RAND_199 = {1{`RANDOM}};
  V1_0 = _RAND_199[15:0];
  _RAND_200 = {1{`RANDOM}};
  V1_1 = _RAND_200[15:0];
  _RAND_201 = {1{`RANDOM}};
  V1_2 = _RAND_201[15:0];
  _RAND_202 = {1{`RANDOM}};
  V1_3 = _RAND_202[15:0];
  _RAND_203 = {1{`RANDOM}};
  V1_4 = _RAND_203[15:0];
  _RAND_204 = {1{`RANDOM}};
  V1_5 = _RAND_204[15:0];
  _RAND_205 = {1{`RANDOM}};
  V1_6 = _RAND_205[15:0];
  _RAND_206 = {1{`RANDOM}};
  V1_7 = _RAND_206[15:0];
  _RAND_207 = {1{`RANDOM}};
  V1_8 = _RAND_207[15:0];
  _RAND_208 = {1{`RANDOM}};
  V1_9 = _RAND_208[15:0];
  _RAND_209 = {1{`RANDOM}};
  V1_10 = _RAND_209[15:0];
  _RAND_210 = {1{`RANDOM}};
  V1_11 = _RAND_210[15:0];
  _RAND_211 = {1{`RANDOM}};
  V1_12 = _RAND_211[15:0];
  _RAND_212 = {1{`RANDOM}};
  V1_13 = _RAND_212[15:0];
  _RAND_213 = {1{`RANDOM}};
  V1_14 = _RAND_213[15:0];
  _RAND_214 = {1{`RANDOM}};
  V1_15 = _RAND_214[15:0];
  _RAND_215 = {1{`RANDOM}};
  V1_16 = _RAND_215[15:0];
  _RAND_216 = {1{`RANDOM}};
  V1_17 = _RAND_216[15:0];
  _RAND_217 = {1{`RANDOM}};
  V1_18 = _RAND_217[15:0];
  _RAND_218 = {1{`RANDOM}};
  V1_19 = _RAND_218[15:0];
  _RAND_219 = {1{`RANDOM}};
  V1_20 = _RAND_219[15:0];
  _RAND_220 = {1{`RANDOM}};
  V1_21 = _RAND_220[15:0];
  _RAND_221 = {1{`RANDOM}};
  V1_22 = _RAND_221[15:0];
  _RAND_222 = {1{`RANDOM}};
  V1_23 = _RAND_222[15:0];
  _RAND_223 = {1{`RANDOM}};
  V1_24 = _RAND_223[15:0];
  _RAND_224 = {1{`RANDOM}};
  V1_25 = _RAND_224[15:0];
  _RAND_225 = {1{`RANDOM}};
  V1_26 = _RAND_225[15:0];
  _RAND_226 = {1{`RANDOM}};
  V1_27 = _RAND_226[15:0];
  _RAND_227 = {1{`RANDOM}};
  V1_28 = _RAND_227[15:0];
  _RAND_228 = {1{`RANDOM}};
  V1_29 = _RAND_228[15:0];
  _RAND_229 = {1{`RANDOM}};
  V1_30 = _RAND_229[15:0];
  _RAND_230 = {1{`RANDOM}};
  V1_31 = _RAND_230[15:0];
  _RAND_231 = {1{`RANDOM}};
  V1_32 = _RAND_231[15:0];
  _RAND_232 = {1{`RANDOM}};
  V1_33 = _RAND_232[15:0];
  _RAND_233 = {1{`RANDOM}};
  V1_34 = _RAND_233[15:0];
  _RAND_234 = {1{`RANDOM}};
  V1_35 = _RAND_234[15:0];
  _RAND_235 = {1{`RANDOM}};
  V1_36 = _RAND_235[15:0];
  _RAND_236 = {1{`RANDOM}};
  V1_37 = _RAND_236[15:0];
  _RAND_237 = {1{`RANDOM}};
  V1_38 = _RAND_237[15:0];
  _RAND_238 = {1{`RANDOM}};
  V1_39 = _RAND_238[15:0];
  _RAND_239 = {1{`RANDOM}};
  V1_40 = _RAND_239[15:0];
  _RAND_240 = {1{`RANDOM}};
  V1_41 = _RAND_240[15:0];
  _RAND_241 = {1{`RANDOM}};
  V1_42 = _RAND_241[15:0];
  _RAND_242 = {1{`RANDOM}};
  V1_43 = _RAND_242[15:0];
  _RAND_243 = {1{`RANDOM}};
  V1_44 = _RAND_243[15:0];
  _RAND_244 = {1{`RANDOM}};
  V1_45 = _RAND_244[15:0];
  _RAND_245 = {1{`RANDOM}};
  V1_46 = _RAND_245[15:0];
  _RAND_246 = {1{`RANDOM}};
  V1_47 = _RAND_246[15:0];
  _RAND_247 = {1{`RANDOM}};
  V1_48 = _RAND_247[15:0];
  _RAND_248 = {1{`RANDOM}};
  V1_49 = _RAND_248[15:0];
  _RAND_249 = {1{`RANDOM}};
  V1_50 = _RAND_249[15:0];
  _RAND_250 = {1{`RANDOM}};
  V1_51 = _RAND_250[15:0];
  _RAND_251 = {1{`RANDOM}};
  V1_52 = _RAND_251[15:0];
  _RAND_252 = {1{`RANDOM}};
  V1_53 = _RAND_252[15:0];
  _RAND_253 = {1{`RANDOM}};
  V1_54 = _RAND_253[15:0];
  _RAND_254 = {1{`RANDOM}};
  V1_55 = _RAND_254[15:0];
  _RAND_255 = {1{`RANDOM}};
  V1_56 = _RAND_255[15:0];
  _RAND_256 = {1{`RANDOM}};
  V1_57 = _RAND_256[15:0];
  _RAND_257 = {1{`RANDOM}};
  V1_58 = _RAND_257[15:0];
  _RAND_258 = {1{`RANDOM}};
  V1_59 = _RAND_258[15:0];
  _RAND_259 = {1{`RANDOM}};
  V1_60 = _RAND_259[15:0];
  _RAND_260 = {1{`RANDOM}};
  V1_61 = _RAND_260[15:0];
  _RAND_261 = {1{`RANDOM}};
  V1_62 = _RAND_261[15:0];
  _RAND_262 = {1{`RANDOM}};
  V1_63 = _RAND_262[15:0];
  _RAND_263 = {1{`RANDOM}};
  V1_64 = _RAND_263[15:0];
  _RAND_264 = {1{`RANDOM}};
  V1_65 = _RAND_264[15:0];
  _RAND_265 = {1{`RANDOM}};
  V1_66 = _RAND_265[15:0];
  _RAND_266 = {1{`RANDOM}};
  V1_67 = _RAND_266[15:0];
  _RAND_267 = {1{`RANDOM}};
  V1_68 = _RAND_267[15:0];
  _RAND_268 = {1{`RANDOM}};
  V1_69 = _RAND_268[15:0];
  _RAND_269 = {1{`RANDOM}};
  V1_70 = _RAND_269[15:0];
  _RAND_270 = {1{`RANDOM}};
  V1_71 = _RAND_270[15:0];
  _RAND_271 = {1{`RANDOM}};
  V1_72 = _RAND_271[15:0];
  _RAND_272 = {1{`RANDOM}};
  V1_73 = _RAND_272[15:0];
  _RAND_273 = {1{`RANDOM}};
  V1_74 = _RAND_273[15:0];
  _RAND_274 = {1{`RANDOM}};
  V1_75 = _RAND_274[15:0];
  _RAND_275 = {1{`RANDOM}};
  V1_76 = _RAND_275[15:0];
  _RAND_276 = {1{`RANDOM}};
  V1_77 = _RAND_276[15:0];
  _RAND_277 = {1{`RANDOM}};
  V1_78 = _RAND_277[15:0];
  _RAND_278 = {1{`RANDOM}};
  V1_79 = _RAND_278[15:0];
  _RAND_279 = {1{`RANDOM}};
  V1_80 = _RAND_279[15:0];
  _RAND_280 = {1{`RANDOM}};
  V1_81 = _RAND_280[15:0];
  _RAND_281 = {1{`RANDOM}};
  V1_82 = _RAND_281[15:0];
  _RAND_282 = {1{`RANDOM}};
  V1_83 = _RAND_282[15:0];
  _RAND_283 = {1{`RANDOM}};
  V1_84 = _RAND_283[15:0];
  _RAND_284 = {1{`RANDOM}};
  V1_85 = _RAND_284[15:0];
  _RAND_285 = {1{`RANDOM}};
  V1_86 = _RAND_285[15:0];
  _RAND_286 = {1{`RANDOM}};
  V1_87 = _RAND_286[15:0];
  _RAND_287 = {1{`RANDOM}};
  V1_88 = _RAND_287[15:0];
  _RAND_288 = {1{`RANDOM}};
  V1_89 = _RAND_288[15:0];
  _RAND_289 = {1{`RANDOM}};
  V1_90 = _RAND_289[15:0];
  _RAND_290 = {1{`RANDOM}};
  V1_91 = _RAND_290[15:0];
  _RAND_291 = {1{`RANDOM}};
  V1_92 = _RAND_291[15:0];
  _RAND_292 = {1{`RANDOM}};
  V1_93 = _RAND_292[15:0];
  _RAND_293 = {1{`RANDOM}};
  V1_94 = _RAND_293[15:0];
  _RAND_294 = {1{`RANDOM}};
  V1_95 = _RAND_294[15:0];
  _RAND_295 = {1{`RANDOM}};
  V1_96 = _RAND_295[15:0];
  _RAND_296 = {1{`RANDOM}};
  V1_97 = _RAND_296[15:0];
  _RAND_297 = {1{`RANDOM}};
  V1_98 = _RAND_297[15:0];
  _RAND_298 = {1{`RANDOM}};
  V1_99 = _RAND_298[15:0];
  _RAND_299 = {1{`RANDOM}};
  V1_100 = _RAND_299[15:0];
  _RAND_300 = {1{`RANDOM}};
  V2_0 = _RAND_300[15:0];
  _RAND_301 = {1{`RANDOM}};
  V2_1 = _RAND_301[15:0];
  _RAND_302 = {1{`RANDOM}};
  V2_2 = _RAND_302[15:0];
  _RAND_303 = {1{`RANDOM}};
  V2_3 = _RAND_303[15:0];
  _RAND_304 = {1{`RANDOM}};
  V2_4 = _RAND_304[15:0];
  _RAND_305 = {1{`RANDOM}};
  V2_5 = _RAND_305[15:0];
  _RAND_306 = {1{`RANDOM}};
  V2_6 = _RAND_306[15:0];
  _RAND_307 = {1{`RANDOM}};
  V2_7 = _RAND_307[15:0];
  _RAND_308 = {1{`RANDOM}};
  V2_8 = _RAND_308[15:0];
  _RAND_309 = {1{`RANDOM}};
  V2_9 = _RAND_309[15:0];
  _RAND_310 = {1{`RANDOM}};
  V2_10 = _RAND_310[15:0];
  _RAND_311 = {1{`RANDOM}};
  V2_11 = _RAND_311[15:0];
  _RAND_312 = {1{`RANDOM}};
  V2_12 = _RAND_312[15:0];
  _RAND_313 = {1{`RANDOM}};
  V2_13 = _RAND_313[15:0];
  _RAND_314 = {1{`RANDOM}};
  V2_14 = _RAND_314[15:0];
  _RAND_315 = {1{`RANDOM}};
  V2_15 = _RAND_315[15:0];
  _RAND_316 = {1{`RANDOM}};
  V2_16 = _RAND_316[15:0];
  _RAND_317 = {1{`RANDOM}};
  V2_17 = _RAND_317[15:0];
  _RAND_318 = {1{`RANDOM}};
  V2_18 = _RAND_318[15:0];
  _RAND_319 = {1{`RANDOM}};
  V2_19 = _RAND_319[15:0];
  _RAND_320 = {1{`RANDOM}};
  V2_20 = _RAND_320[15:0];
  _RAND_321 = {1{`RANDOM}};
  V2_21 = _RAND_321[15:0];
  _RAND_322 = {1{`RANDOM}};
  V2_22 = _RAND_322[15:0];
  _RAND_323 = {1{`RANDOM}};
  V2_23 = _RAND_323[15:0];
  _RAND_324 = {1{`RANDOM}};
  V2_24 = _RAND_324[15:0];
  _RAND_325 = {1{`RANDOM}};
  V2_25 = _RAND_325[15:0];
  _RAND_326 = {1{`RANDOM}};
  V2_26 = _RAND_326[15:0];
  _RAND_327 = {1{`RANDOM}};
  V2_27 = _RAND_327[15:0];
  _RAND_328 = {1{`RANDOM}};
  V2_28 = _RAND_328[15:0];
  _RAND_329 = {1{`RANDOM}};
  V2_29 = _RAND_329[15:0];
  _RAND_330 = {1{`RANDOM}};
  V2_30 = _RAND_330[15:0];
  _RAND_331 = {1{`RANDOM}};
  V2_31 = _RAND_331[15:0];
  _RAND_332 = {1{`RANDOM}};
  V2_32 = _RAND_332[15:0];
  _RAND_333 = {1{`RANDOM}};
  V2_33 = _RAND_333[15:0];
  _RAND_334 = {1{`RANDOM}};
  V2_34 = _RAND_334[15:0];
  _RAND_335 = {1{`RANDOM}};
  V2_35 = _RAND_335[15:0];
  _RAND_336 = {1{`RANDOM}};
  V2_36 = _RAND_336[15:0];
  _RAND_337 = {1{`RANDOM}};
  V2_37 = _RAND_337[15:0];
  _RAND_338 = {1{`RANDOM}};
  V2_38 = _RAND_338[15:0];
  _RAND_339 = {1{`RANDOM}};
  V2_39 = _RAND_339[15:0];
  _RAND_340 = {1{`RANDOM}};
  V2_40 = _RAND_340[15:0];
  _RAND_341 = {1{`RANDOM}};
  V2_41 = _RAND_341[15:0];
  _RAND_342 = {1{`RANDOM}};
  V2_42 = _RAND_342[15:0];
  _RAND_343 = {1{`RANDOM}};
  V2_43 = _RAND_343[15:0];
  _RAND_344 = {1{`RANDOM}};
  V2_44 = _RAND_344[15:0];
  _RAND_345 = {1{`RANDOM}};
  V2_45 = _RAND_345[15:0];
  _RAND_346 = {1{`RANDOM}};
  V2_46 = _RAND_346[15:0];
  _RAND_347 = {1{`RANDOM}};
  V2_47 = _RAND_347[15:0];
  _RAND_348 = {1{`RANDOM}};
  V2_48 = _RAND_348[15:0];
  _RAND_349 = {1{`RANDOM}};
  V2_49 = _RAND_349[15:0];
  _RAND_350 = {1{`RANDOM}};
  V2_50 = _RAND_350[15:0];
  _RAND_351 = {1{`RANDOM}};
  V2_51 = _RAND_351[15:0];
  _RAND_352 = {1{`RANDOM}};
  V2_52 = _RAND_352[15:0];
  _RAND_353 = {1{`RANDOM}};
  V2_53 = _RAND_353[15:0];
  _RAND_354 = {1{`RANDOM}};
  V2_54 = _RAND_354[15:0];
  _RAND_355 = {1{`RANDOM}};
  V2_55 = _RAND_355[15:0];
  _RAND_356 = {1{`RANDOM}};
  V2_56 = _RAND_356[15:0];
  _RAND_357 = {1{`RANDOM}};
  V2_57 = _RAND_357[15:0];
  _RAND_358 = {1{`RANDOM}};
  V2_58 = _RAND_358[15:0];
  _RAND_359 = {1{`RANDOM}};
  V2_59 = _RAND_359[15:0];
  _RAND_360 = {1{`RANDOM}};
  V2_60 = _RAND_360[15:0];
  _RAND_361 = {1{`RANDOM}};
  V2_61 = _RAND_361[15:0];
  _RAND_362 = {1{`RANDOM}};
  V2_62 = _RAND_362[15:0];
  _RAND_363 = {1{`RANDOM}};
  V2_63 = _RAND_363[15:0];
  _RAND_364 = {1{`RANDOM}};
  V2_64 = _RAND_364[15:0];
  _RAND_365 = {1{`RANDOM}};
  V2_65 = _RAND_365[15:0];
  _RAND_366 = {1{`RANDOM}};
  V2_66 = _RAND_366[15:0];
  _RAND_367 = {1{`RANDOM}};
  V2_67 = _RAND_367[15:0];
  _RAND_368 = {1{`RANDOM}};
  V2_68 = _RAND_368[15:0];
  _RAND_369 = {1{`RANDOM}};
  V2_69 = _RAND_369[15:0];
  _RAND_370 = {1{`RANDOM}};
  V2_70 = _RAND_370[15:0];
  _RAND_371 = {1{`RANDOM}};
  V2_71 = _RAND_371[15:0];
  _RAND_372 = {1{`RANDOM}};
  V2_72 = _RAND_372[15:0];
  _RAND_373 = {1{`RANDOM}};
  V2_73 = _RAND_373[15:0];
  _RAND_374 = {1{`RANDOM}};
  V2_74 = _RAND_374[15:0];
  _RAND_375 = {1{`RANDOM}};
  V2_75 = _RAND_375[15:0];
  _RAND_376 = {1{`RANDOM}};
  V2_76 = _RAND_376[15:0];
  _RAND_377 = {1{`RANDOM}};
  V2_77 = _RAND_377[15:0];
  _RAND_378 = {1{`RANDOM}};
  V2_78 = _RAND_378[15:0];
  _RAND_379 = {1{`RANDOM}};
  V2_79 = _RAND_379[15:0];
  _RAND_380 = {1{`RANDOM}};
  V2_80 = _RAND_380[15:0];
  _RAND_381 = {1{`RANDOM}};
  V2_81 = _RAND_381[15:0];
  _RAND_382 = {1{`RANDOM}};
  V2_82 = _RAND_382[15:0];
  _RAND_383 = {1{`RANDOM}};
  V2_83 = _RAND_383[15:0];
  _RAND_384 = {1{`RANDOM}};
  V2_84 = _RAND_384[15:0];
  _RAND_385 = {1{`RANDOM}};
  V2_85 = _RAND_385[15:0];
  _RAND_386 = {1{`RANDOM}};
  V2_86 = _RAND_386[15:0];
  _RAND_387 = {1{`RANDOM}};
  V2_87 = _RAND_387[15:0];
  _RAND_388 = {1{`RANDOM}};
  V2_88 = _RAND_388[15:0];
  _RAND_389 = {1{`RANDOM}};
  V2_89 = _RAND_389[15:0];
  _RAND_390 = {1{`RANDOM}};
  V2_90 = _RAND_390[15:0];
  _RAND_391 = {1{`RANDOM}};
  V2_91 = _RAND_391[15:0];
  _RAND_392 = {1{`RANDOM}};
  V2_92 = _RAND_392[15:0];
  _RAND_393 = {1{`RANDOM}};
  V2_93 = _RAND_393[15:0];
  _RAND_394 = {1{`RANDOM}};
  V2_94 = _RAND_394[15:0];
  _RAND_395 = {1{`RANDOM}};
  V2_95 = _RAND_395[15:0];
  _RAND_396 = {1{`RANDOM}};
  V2_96 = _RAND_396[15:0];
  _RAND_397 = {1{`RANDOM}};
  V2_97 = _RAND_397[15:0];
  _RAND_398 = {1{`RANDOM}};
  V2_98 = _RAND_398[15:0];
  _RAND_399 = {1{`RANDOM}};
  V2_99 = _RAND_399[15:0];
  _RAND_400 = {1{`RANDOM}};
  start_reg_0 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  start_reg_1 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  start_reg_2 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  start_reg_3 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  start_reg_4 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  start_reg_5 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  start_reg_6 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  start_reg_7 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  start_reg_8 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  start_reg_9 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  start_reg_10 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  start_reg_11 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  start_reg_12 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  start_reg_13 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  start_reg_14 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  start_reg_15 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  start_reg_16 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  start_reg_17 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  start_reg_18 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  start_reg_19 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  start_reg_20 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  start_reg_21 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  start_reg_22 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  start_reg_23 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  start_reg_24 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  start_reg_25 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  start_reg_26 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  start_reg_27 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  start_reg_28 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  start_reg_29 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  start_reg_30 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  start_reg_31 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  start_reg_32 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  start_reg_33 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  start_reg_34 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  start_reg_35 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  start_reg_36 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  start_reg_37 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  start_reg_38 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  start_reg_39 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  start_reg_40 = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  start_reg_41 = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  start_reg_42 = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  start_reg_43 = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  start_reg_44 = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  start_reg_45 = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  start_reg_46 = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  start_reg_47 = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  start_reg_48 = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  start_reg_49 = _RAND_449[0:0];
  _RAND_450 = {1{`RANDOM}};
  start_reg_50 = _RAND_450[0:0];
  _RAND_451 = {1{`RANDOM}};
  start_reg_51 = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  start_reg_52 = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  start_reg_53 = _RAND_453[0:0];
  _RAND_454 = {1{`RANDOM}};
  start_reg_54 = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  start_reg_55 = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  start_reg_56 = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  start_reg_57 = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  start_reg_58 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  start_reg_59 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  start_reg_60 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  start_reg_61 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  start_reg_62 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  start_reg_63 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  start_reg_64 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  start_reg_65 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  start_reg_66 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  start_reg_67 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  start_reg_68 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  start_reg_69 = _RAND_469[0:0];
  _RAND_470 = {1{`RANDOM}};
  start_reg_70 = _RAND_470[0:0];
  _RAND_471 = {1{`RANDOM}};
  start_reg_71 = _RAND_471[0:0];
  _RAND_472 = {1{`RANDOM}};
  start_reg_72 = _RAND_472[0:0];
  _RAND_473 = {1{`RANDOM}};
  start_reg_73 = _RAND_473[0:0];
  _RAND_474 = {1{`RANDOM}};
  start_reg_74 = _RAND_474[0:0];
  _RAND_475 = {1{`RANDOM}};
  start_reg_75 = _RAND_475[0:0];
  _RAND_476 = {1{`RANDOM}};
  start_reg_76 = _RAND_476[0:0];
  _RAND_477 = {1{`RANDOM}};
  start_reg_77 = _RAND_477[0:0];
  _RAND_478 = {1{`RANDOM}};
  start_reg_78 = _RAND_478[0:0];
  _RAND_479 = {1{`RANDOM}};
  start_reg_79 = _RAND_479[0:0];
  _RAND_480 = {1{`RANDOM}};
  start_reg_80 = _RAND_480[0:0];
  _RAND_481 = {1{`RANDOM}};
  start_reg_81 = _RAND_481[0:0];
  _RAND_482 = {1{`RANDOM}};
  start_reg_82 = _RAND_482[0:0];
  _RAND_483 = {1{`RANDOM}};
  start_reg_83 = _RAND_483[0:0];
  _RAND_484 = {1{`RANDOM}};
  start_reg_84 = _RAND_484[0:0];
  _RAND_485 = {1{`RANDOM}};
  start_reg_85 = _RAND_485[0:0];
  _RAND_486 = {1{`RANDOM}};
  start_reg_86 = _RAND_486[0:0];
  _RAND_487 = {1{`RANDOM}};
  start_reg_87 = _RAND_487[0:0];
  _RAND_488 = {1{`RANDOM}};
  start_reg_88 = _RAND_488[0:0];
  _RAND_489 = {1{`RANDOM}};
  start_reg_89 = _RAND_489[0:0];
  _RAND_490 = {1{`RANDOM}};
  start_reg_90 = _RAND_490[0:0];
  _RAND_491 = {1{`RANDOM}};
  start_reg_91 = _RAND_491[0:0];
  _RAND_492 = {1{`RANDOM}};
  start_reg_92 = _RAND_492[0:0];
  _RAND_493 = {1{`RANDOM}};
  start_reg_93 = _RAND_493[0:0];
  _RAND_494 = {1{`RANDOM}};
  start_reg_94 = _RAND_494[0:0];
  _RAND_495 = {1{`RANDOM}};
  start_reg_95 = _RAND_495[0:0];
  _RAND_496 = {1{`RANDOM}};
  start_reg_96 = _RAND_496[0:0];
  _RAND_497 = {1{`RANDOM}};
  start_reg_97 = _RAND_497[0:0];
  _RAND_498 = {1{`RANDOM}};
  start_reg_98 = _RAND_498[0:0];
  _RAND_499 = {1{`RANDOM}};
  start_reg_99 = _RAND_499[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
