module SWCell(
  input  [1:0]  io_q,
  input  [1:0]  io_r,
  input  [15:0] io_e_i,
  input  [15:0] io_f_i,
  input  [15:0] io_ve_i,
  input  [15:0] io_vf_i,
  input  [15:0] io_vv_i,
  output [15:0] io_e_o,
  output [15:0] io_f_o,
  output [15:0] io_v_o
);
  wire [15:0] _T_2 = $signed(io_ve_i) - 16'sh2; // @[SWChisel.scala 78:17]
  wire [15:0] _T_5 = $signed(io_e_i) - 16'sh1; // @[SWChisel.scala 78:39]
  wire [15:0] e_max = $signed(_T_2) >= $signed(_T_5) ? $signed(_T_2) : $signed(_T_5); // @[SWChisel.scala 78:51 79:11 81:11]
  wire [15:0] _T_9 = $signed(io_vf_i) - 16'sh2; // @[SWChisel.scala 85:17]
  wire [15:0] _T_12 = $signed(io_f_i) - 16'sh1; // @[SWChisel.scala 85:38]
  wire [15:0] f_max = $signed(_T_9) > $signed(_T_12) ? $signed(_T_9) : $signed(_T_12); // @[SWChisel.scala 85:50 86:11 88:11]
  wire [15:0] ef_temp = $signed(e_max) > $signed(f_max) ? $signed(e_max) : $signed(f_max); // @[SWChisel.scala 92:24 93:13 95:13]
  wire [15:0] _v_temp_T_2 = $signed(io_vv_i) + 16'sh2; // @[SWChisel.scala 100:23]
  wire [15:0] _v_temp_T_5 = $signed(io_vv_i) - 16'sh2; // @[SWChisel.scala 102:23]
  wire [15:0] v_temp = io_q == io_r ? $signed(_v_temp_T_2) : $signed(_v_temp_T_5); // @[SWChisel.scala 100:12 102:12 99:24]
  assign io_e_o = $signed(_T_2) >= $signed(_T_5) ? $signed(_T_2) : $signed(_T_5); // @[SWChisel.scala 78:51 79:11 81:11]
  assign io_f_o = $signed(_T_9) > $signed(_T_12) ? $signed(_T_9) : $signed(_T_12); // @[SWChisel.scala 85:50 86:11 88:11]
  assign io_v_o = $signed(v_temp) > $signed(ef_temp) ? $signed(v_temp) : $signed(ef_temp); // @[SWChisel.scala 106:27 107:11 109:11]
endmodule
module MyCounter(
  input        clock,
  input        reset,
  input        io_en,
  output [7:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] _io_out_T_2 = io_out + 8'h1; // @[SWChisel.scala 155:55]
  reg [7:0] io_out_r; // @[Reg.scala 35:20]
  assign io_out = io_out_r; // @[SWChisel.scala 155:12]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      io_out_r <= 8'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_out < 8'hc8) begin // @[SWChisel.scala 155:28]
        io_out_r <= _io_out_T_2;
      end else begin
        io_out_r <= 8'h0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_out_r = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MAX(
  input         clock,
  input         reset,
  input         io_start,
  input  [15:0] io_in,
  output        io_done,
  output [15:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] max; // @[SWChisel.scala 122:20]
  reg [7:0] counter; // @[SWChisel.scala 133:24]
  wire [7:0] _counter_T_1 = counter - 8'h1; // @[SWChisel.scala 135:24]
  assign io_done = counter == 8'h0; // @[SWChisel.scala 141:17]
  assign io_out = max; // @[SWChisel.scala 123:10]
  always @(posedge clock) begin
    if (reset) begin // @[SWChisel.scala 122:20]
      max <= 16'sh8000; // @[SWChisel.scala 122:20]
    end else if ($signed(io_in) > $signed(max)) begin // @[SWChisel.scala 126:22]
      max <= io_in; // @[SWChisel.scala 127:9]
    end
    if (reset) begin // @[SWChisel.scala 133:24]
      counter <= 8'hc9; // @[SWChisel.scala 133:24]
    end else if (counter == 8'h0) begin // @[SWChisel.scala 141:26]
      counter <= 8'h0; // @[SWChisel.scala 143:13]
    end else if (io_start) begin // @[SWChisel.scala 134:19]
      counter <= _counter_T_1; // @[SWChisel.scala 135:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  max = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  counter = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SW(
  input         clock,
  input         reset,
  input  [1:0]  io_q_0_b,
  input  [1:0]  io_q_1_b,
  input  [1:0]  io_q_2_b,
  input  [1:0]  io_q_3_b,
  input  [1:0]  io_q_4_b,
  input  [1:0]  io_q_5_b,
  input  [1:0]  io_q_6_b,
  input  [1:0]  io_q_7_b,
  input  [1:0]  io_q_8_b,
  input  [1:0]  io_q_9_b,
  input  [1:0]  io_q_10_b,
  input  [1:0]  io_q_11_b,
  input  [1:0]  io_q_12_b,
  input  [1:0]  io_q_13_b,
  input  [1:0]  io_q_14_b,
  input  [1:0]  io_q_15_b,
  input  [1:0]  io_q_16_b,
  input  [1:0]  io_q_17_b,
  input  [1:0]  io_q_18_b,
  input  [1:0]  io_q_19_b,
  input  [1:0]  io_q_20_b,
  input  [1:0]  io_q_21_b,
  input  [1:0]  io_q_22_b,
  input  [1:0]  io_q_23_b,
  input  [1:0]  io_q_24_b,
  input  [1:0]  io_q_25_b,
  input  [1:0]  io_q_26_b,
  input  [1:0]  io_q_27_b,
  input  [1:0]  io_q_28_b,
  input  [1:0]  io_q_29_b,
  input  [1:0]  io_q_30_b,
  input  [1:0]  io_q_31_b,
  input  [1:0]  io_q_32_b,
  input  [1:0]  io_q_33_b,
  input  [1:0]  io_q_34_b,
  input  [1:0]  io_q_35_b,
  input  [1:0]  io_q_36_b,
  input  [1:0]  io_q_37_b,
  input  [1:0]  io_q_38_b,
  input  [1:0]  io_q_39_b,
  input  [1:0]  io_r_0_b,
  input  [1:0]  io_r_1_b,
  input  [1:0]  io_r_2_b,
  input  [1:0]  io_r_3_b,
  input  [1:0]  io_r_4_b,
  input  [1:0]  io_r_5_b,
  input  [1:0]  io_r_6_b,
  input  [1:0]  io_r_7_b,
  input  [1:0]  io_r_8_b,
  input  [1:0]  io_r_9_b,
  input  [1:0]  io_r_10_b,
  input  [1:0]  io_r_11_b,
  input  [1:0]  io_r_12_b,
  input  [1:0]  io_r_13_b,
  input  [1:0]  io_r_14_b,
  input  [1:0]  io_r_15_b,
  input  [1:0]  io_r_16_b,
  input  [1:0]  io_r_17_b,
  input  [1:0]  io_r_18_b,
  input  [1:0]  io_r_19_b,
  input  [1:0]  io_r_20_b,
  input  [1:0]  io_r_21_b,
  input  [1:0]  io_r_22_b,
  input  [1:0]  io_r_23_b,
  input  [1:0]  io_r_24_b,
  input  [1:0]  io_r_25_b,
  input  [1:0]  io_r_26_b,
  input  [1:0]  io_r_27_b,
  input  [1:0]  io_r_28_b,
  input  [1:0]  io_r_29_b,
  input  [1:0]  io_r_30_b,
  input  [1:0]  io_r_31_b,
  input  [1:0]  io_r_32_b,
  input  [1:0]  io_r_33_b,
  input  [1:0]  io_r_34_b,
  input  [1:0]  io_r_35_b,
  input  [1:0]  io_r_36_b,
  input  [1:0]  io_r_37_b,
  input  [1:0]  io_r_38_b,
  input  [1:0]  io_r_39_b,
  input  [1:0]  io_r_40_b,
  input  [1:0]  io_r_41_b,
  input  [1:0]  io_r_42_b,
  input  [1:0]  io_r_43_b,
  input  [1:0]  io_r_44_b,
  input  [1:0]  io_r_45_b,
  input  [1:0]  io_r_46_b,
  input  [1:0]  io_r_47_b,
  input  [1:0]  io_r_48_b,
  input  [1:0]  io_r_49_b,
  input  [1:0]  io_r_50_b,
  input  [1:0]  io_r_51_b,
  input  [1:0]  io_r_52_b,
  input  [1:0]  io_r_53_b,
  input  [1:0]  io_r_54_b,
  input  [1:0]  io_r_55_b,
  input  [1:0]  io_r_56_b,
  input  [1:0]  io_r_57_b,
  input  [1:0]  io_r_58_b,
  input  [1:0]  io_r_59_b,
  input  [1:0]  io_r_60_b,
  input  [1:0]  io_r_61_b,
  input  [1:0]  io_r_62_b,
  input  [1:0]  io_r_63_b,
  input  [1:0]  io_r_64_b,
  input  [1:0]  io_r_65_b,
  input  [1:0]  io_r_66_b,
  input  [1:0]  io_r_67_b,
  input  [1:0]  io_r_68_b,
  input  [1:0]  io_r_69_b,
  input  [1:0]  io_r_70_b,
  input  [1:0]  io_r_71_b,
  input  [1:0]  io_r_72_b,
  input  [1:0]  io_r_73_b,
  input  [1:0]  io_r_74_b,
  input  [1:0]  io_r_75_b,
  input  [1:0]  io_r_76_b,
  input  [1:0]  io_r_77_b,
  input  [1:0]  io_r_78_b,
  input  [1:0]  io_r_79_b,
  input  [1:0]  io_r_80_b,
  input  [1:0]  io_r_81_b,
  input  [1:0]  io_r_82_b,
  input  [1:0]  io_r_83_b,
  input  [1:0]  io_r_84_b,
  input  [1:0]  io_r_85_b,
  input  [1:0]  io_r_86_b,
  input  [1:0]  io_r_87_b,
  input  [1:0]  io_r_88_b,
  input  [1:0]  io_r_89_b,
  input  [1:0]  io_r_90_b,
  input  [1:0]  io_r_91_b,
  input  [1:0]  io_r_92_b,
  input  [1:0]  io_r_93_b,
  input  [1:0]  io_r_94_b,
  input  [1:0]  io_r_95_b,
  input  [1:0]  io_r_96_b,
  input  [1:0]  io_r_97_b,
  input  [1:0]  io_r_98_b,
  input  [1:0]  io_r_99_b,
  input  [1:0]  io_r_100_b,
  input  [1:0]  io_r_101_b,
  input  [1:0]  io_r_102_b,
  input  [1:0]  io_r_103_b,
  input  [1:0]  io_r_104_b,
  input  [1:0]  io_r_105_b,
  input  [1:0]  io_r_106_b,
  input  [1:0]  io_r_107_b,
  input  [1:0]  io_r_108_b,
  input  [1:0]  io_r_109_b,
  input  [1:0]  io_r_110_b,
  input  [1:0]  io_r_111_b,
  input  [1:0]  io_r_112_b,
  input  [1:0]  io_r_113_b,
  input  [1:0]  io_r_114_b,
  input  [1:0]  io_r_115_b,
  input  [1:0]  io_r_116_b,
  input  [1:0]  io_r_117_b,
  input  [1:0]  io_r_118_b,
  input  [1:0]  io_r_119_b,
  input  [1:0]  io_r_120_b,
  input  [1:0]  io_r_121_b,
  input  [1:0]  io_r_122_b,
  input  [1:0]  io_r_123_b,
  input  [1:0]  io_r_124_b,
  input  [1:0]  io_r_125_b,
  input  [1:0]  io_r_126_b,
  input  [1:0]  io_r_127_b,
  input  [1:0]  io_r_128_b,
  input  [1:0]  io_r_129_b,
  input  [1:0]  io_r_130_b,
  input  [1:0]  io_r_131_b,
  input  [1:0]  io_r_132_b,
  input  [1:0]  io_r_133_b,
  input  [1:0]  io_r_134_b,
  input  [1:0]  io_r_135_b,
  input  [1:0]  io_r_136_b,
  input  [1:0]  io_r_137_b,
  input  [1:0]  io_r_138_b,
  input  [1:0]  io_r_139_b,
  input  [1:0]  io_r_140_b,
  input  [1:0]  io_r_141_b,
  input  [1:0]  io_r_142_b,
  input  [1:0]  io_r_143_b,
  input  [1:0]  io_r_144_b,
  input  [1:0]  io_r_145_b,
  input  [1:0]  io_r_146_b,
  input  [1:0]  io_r_147_b,
  input  [1:0]  io_r_148_b,
  input  [1:0]  io_r_149_b,
  input  [1:0]  io_r_150_b,
  input  [1:0]  io_r_151_b,
  input  [1:0]  io_r_152_b,
  input  [1:0]  io_r_153_b,
  input  [1:0]  io_r_154_b,
  input  [1:0]  io_r_155_b,
  input  [1:0]  io_r_156_b,
  input  [1:0]  io_r_157_b,
  input  [1:0]  io_r_158_b,
  input  [1:0]  io_r_159_b,
  input  [1:0]  io_r_160_b,
  input  [1:0]  io_r_161_b,
  input  [1:0]  io_r_162_b,
  input  [1:0]  io_r_163_b,
  input  [1:0]  io_r_164_b,
  input  [1:0]  io_r_165_b,
  input  [1:0]  io_r_166_b,
  input  [1:0]  io_r_167_b,
  input  [1:0]  io_r_168_b,
  input  [1:0]  io_r_169_b,
  input  [1:0]  io_r_170_b,
  input  [1:0]  io_r_171_b,
  input  [1:0]  io_r_172_b,
  input  [1:0]  io_r_173_b,
  input  [1:0]  io_r_174_b,
  input  [1:0]  io_r_175_b,
  input  [1:0]  io_r_176_b,
  input  [1:0]  io_r_177_b,
  input  [1:0]  io_r_178_b,
  input  [1:0]  io_r_179_b,
  input  [1:0]  io_r_180_b,
  input  [1:0]  io_r_181_b,
  input  [1:0]  io_r_182_b,
  input  [1:0]  io_r_183_b,
  input  [1:0]  io_r_184_b,
  input  [1:0]  io_r_185_b,
  input  [1:0]  io_r_186_b,
  input  [1:0]  io_r_187_b,
  input  [1:0]  io_r_188_b,
  input  [1:0]  io_r_189_b,
  input  [1:0]  io_r_190_b,
  input  [1:0]  io_r_191_b,
  input  [1:0]  io_r_192_b,
  input  [1:0]  io_r_193_b,
  input  [1:0]  io_r_194_b,
  input  [1:0]  io_r_195_b,
  input  [1:0]  io_r_196_b,
  input  [1:0]  io_r_197_b,
  input  [1:0]  io_r_198_b,
  input  [1:0]  io_r_199_b,
  input         io_start,
  output [15:0] io_result,
  output        io_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
`endif // RANDOMIZE_REG_INIT
  wire [1:0] array_0_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_0_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_1_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_1_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_2_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_2_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_3_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_3_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_4_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_4_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_5_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_5_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_6_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_6_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_7_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_7_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_8_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_8_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_9_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_9_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_10_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_10_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_11_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_11_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_12_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_12_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_13_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_13_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_14_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_14_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_15_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_15_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_16_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_16_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_17_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_17_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_18_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_18_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_19_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_19_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_20_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_20_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_21_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_21_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_22_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_22_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_23_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_23_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_24_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_24_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_25_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_25_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_26_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_26_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_27_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_27_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_28_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_28_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_29_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_29_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_30_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_30_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_31_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_31_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_32_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_32_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_33_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_33_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_34_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_34_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_35_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_35_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_36_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_36_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_37_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_37_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_38_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_38_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_39_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_39_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_v_o; // @[SWChisel.scala 170:39]
  wire  r_count_0_clock; // @[SWChisel.scala 171:41]
  wire  r_count_0_reset; // @[SWChisel.scala 171:41]
  wire  r_count_0_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_0_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_1_clock; // @[SWChisel.scala 171:41]
  wire  r_count_1_reset; // @[SWChisel.scala 171:41]
  wire  r_count_1_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_1_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_2_clock; // @[SWChisel.scala 171:41]
  wire  r_count_2_reset; // @[SWChisel.scala 171:41]
  wire  r_count_2_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_2_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_3_clock; // @[SWChisel.scala 171:41]
  wire  r_count_3_reset; // @[SWChisel.scala 171:41]
  wire  r_count_3_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_3_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_4_clock; // @[SWChisel.scala 171:41]
  wire  r_count_4_reset; // @[SWChisel.scala 171:41]
  wire  r_count_4_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_4_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_5_clock; // @[SWChisel.scala 171:41]
  wire  r_count_5_reset; // @[SWChisel.scala 171:41]
  wire  r_count_5_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_5_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_6_clock; // @[SWChisel.scala 171:41]
  wire  r_count_6_reset; // @[SWChisel.scala 171:41]
  wire  r_count_6_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_6_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_7_clock; // @[SWChisel.scala 171:41]
  wire  r_count_7_reset; // @[SWChisel.scala 171:41]
  wire  r_count_7_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_7_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_8_clock; // @[SWChisel.scala 171:41]
  wire  r_count_8_reset; // @[SWChisel.scala 171:41]
  wire  r_count_8_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_8_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_9_clock; // @[SWChisel.scala 171:41]
  wire  r_count_9_reset; // @[SWChisel.scala 171:41]
  wire  r_count_9_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_9_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_10_clock; // @[SWChisel.scala 171:41]
  wire  r_count_10_reset; // @[SWChisel.scala 171:41]
  wire  r_count_10_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_10_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_11_clock; // @[SWChisel.scala 171:41]
  wire  r_count_11_reset; // @[SWChisel.scala 171:41]
  wire  r_count_11_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_11_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_12_clock; // @[SWChisel.scala 171:41]
  wire  r_count_12_reset; // @[SWChisel.scala 171:41]
  wire  r_count_12_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_12_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_13_clock; // @[SWChisel.scala 171:41]
  wire  r_count_13_reset; // @[SWChisel.scala 171:41]
  wire  r_count_13_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_13_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_14_clock; // @[SWChisel.scala 171:41]
  wire  r_count_14_reset; // @[SWChisel.scala 171:41]
  wire  r_count_14_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_14_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_15_clock; // @[SWChisel.scala 171:41]
  wire  r_count_15_reset; // @[SWChisel.scala 171:41]
  wire  r_count_15_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_15_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_16_clock; // @[SWChisel.scala 171:41]
  wire  r_count_16_reset; // @[SWChisel.scala 171:41]
  wire  r_count_16_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_16_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_17_clock; // @[SWChisel.scala 171:41]
  wire  r_count_17_reset; // @[SWChisel.scala 171:41]
  wire  r_count_17_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_17_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_18_clock; // @[SWChisel.scala 171:41]
  wire  r_count_18_reset; // @[SWChisel.scala 171:41]
  wire  r_count_18_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_18_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_19_clock; // @[SWChisel.scala 171:41]
  wire  r_count_19_reset; // @[SWChisel.scala 171:41]
  wire  r_count_19_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_19_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_20_clock; // @[SWChisel.scala 171:41]
  wire  r_count_20_reset; // @[SWChisel.scala 171:41]
  wire  r_count_20_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_20_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_21_clock; // @[SWChisel.scala 171:41]
  wire  r_count_21_reset; // @[SWChisel.scala 171:41]
  wire  r_count_21_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_21_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_22_clock; // @[SWChisel.scala 171:41]
  wire  r_count_22_reset; // @[SWChisel.scala 171:41]
  wire  r_count_22_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_22_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_23_clock; // @[SWChisel.scala 171:41]
  wire  r_count_23_reset; // @[SWChisel.scala 171:41]
  wire  r_count_23_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_23_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_24_clock; // @[SWChisel.scala 171:41]
  wire  r_count_24_reset; // @[SWChisel.scala 171:41]
  wire  r_count_24_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_24_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_25_clock; // @[SWChisel.scala 171:41]
  wire  r_count_25_reset; // @[SWChisel.scala 171:41]
  wire  r_count_25_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_25_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_26_clock; // @[SWChisel.scala 171:41]
  wire  r_count_26_reset; // @[SWChisel.scala 171:41]
  wire  r_count_26_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_26_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_27_clock; // @[SWChisel.scala 171:41]
  wire  r_count_27_reset; // @[SWChisel.scala 171:41]
  wire  r_count_27_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_27_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_28_clock; // @[SWChisel.scala 171:41]
  wire  r_count_28_reset; // @[SWChisel.scala 171:41]
  wire  r_count_28_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_28_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_29_clock; // @[SWChisel.scala 171:41]
  wire  r_count_29_reset; // @[SWChisel.scala 171:41]
  wire  r_count_29_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_29_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_30_clock; // @[SWChisel.scala 171:41]
  wire  r_count_30_reset; // @[SWChisel.scala 171:41]
  wire  r_count_30_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_30_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_31_clock; // @[SWChisel.scala 171:41]
  wire  r_count_31_reset; // @[SWChisel.scala 171:41]
  wire  r_count_31_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_31_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_32_clock; // @[SWChisel.scala 171:41]
  wire  r_count_32_reset; // @[SWChisel.scala 171:41]
  wire  r_count_32_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_32_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_33_clock; // @[SWChisel.scala 171:41]
  wire  r_count_33_reset; // @[SWChisel.scala 171:41]
  wire  r_count_33_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_33_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_34_clock; // @[SWChisel.scala 171:41]
  wire  r_count_34_reset; // @[SWChisel.scala 171:41]
  wire  r_count_34_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_34_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_35_clock; // @[SWChisel.scala 171:41]
  wire  r_count_35_reset; // @[SWChisel.scala 171:41]
  wire  r_count_35_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_35_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_36_clock; // @[SWChisel.scala 171:41]
  wire  r_count_36_reset; // @[SWChisel.scala 171:41]
  wire  r_count_36_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_36_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_37_clock; // @[SWChisel.scala 171:41]
  wire  r_count_37_reset; // @[SWChisel.scala 171:41]
  wire  r_count_37_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_37_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_38_clock; // @[SWChisel.scala 171:41]
  wire  r_count_38_reset; // @[SWChisel.scala 171:41]
  wire  r_count_38_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_38_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_39_clock; // @[SWChisel.scala 171:41]
  wire  r_count_39_reset; // @[SWChisel.scala 171:41]
  wire  r_count_39_io_en; // @[SWChisel.scala 171:41]
  wire [7:0] r_count_39_io_out; // @[SWChisel.scala 171:41]
  wire  max_clock; // @[SWChisel.scala 174:19]
  wire  max_reset; // @[SWChisel.scala 174:19]
  wire  max_io_start; // @[SWChisel.scala 174:19]
  wire [15:0] max_io_in; // @[SWChisel.scala 174:19]
  wire  max_io_done; // @[SWChisel.scala 174:19]
  wire [15:0] max_io_out; // @[SWChisel.scala 174:19]
  reg [15:0] E_0; // @[SWChisel.scala 162:18]
  reg [15:0] E_1; // @[SWChisel.scala 162:18]
  reg [15:0] E_2; // @[SWChisel.scala 162:18]
  reg [15:0] E_3; // @[SWChisel.scala 162:18]
  reg [15:0] E_4; // @[SWChisel.scala 162:18]
  reg [15:0] E_5; // @[SWChisel.scala 162:18]
  reg [15:0] E_6; // @[SWChisel.scala 162:18]
  reg [15:0] E_7; // @[SWChisel.scala 162:18]
  reg [15:0] E_8; // @[SWChisel.scala 162:18]
  reg [15:0] E_9; // @[SWChisel.scala 162:18]
  reg [15:0] E_10; // @[SWChisel.scala 162:18]
  reg [15:0] E_11; // @[SWChisel.scala 162:18]
  reg [15:0] E_12; // @[SWChisel.scala 162:18]
  reg [15:0] E_13; // @[SWChisel.scala 162:18]
  reg [15:0] E_14; // @[SWChisel.scala 162:18]
  reg [15:0] E_15; // @[SWChisel.scala 162:18]
  reg [15:0] E_16; // @[SWChisel.scala 162:18]
  reg [15:0] E_17; // @[SWChisel.scala 162:18]
  reg [15:0] E_18; // @[SWChisel.scala 162:18]
  reg [15:0] E_19; // @[SWChisel.scala 162:18]
  reg [15:0] E_20; // @[SWChisel.scala 162:18]
  reg [15:0] E_21; // @[SWChisel.scala 162:18]
  reg [15:0] E_22; // @[SWChisel.scala 162:18]
  reg [15:0] E_23; // @[SWChisel.scala 162:18]
  reg [15:0] E_24; // @[SWChisel.scala 162:18]
  reg [15:0] E_25; // @[SWChisel.scala 162:18]
  reg [15:0] E_26; // @[SWChisel.scala 162:18]
  reg [15:0] E_27; // @[SWChisel.scala 162:18]
  reg [15:0] E_28; // @[SWChisel.scala 162:18]
  reg [15:0] E_29; // @[SWChisel.scala 162:18]
  reg [15:0] E_30; // @[SWChisel.scala 162:18]
  reg [15:0] E_31; // @[SWChisel.scala 162:18]
  reg [15:0] E_32; // @[SWChisel.scala 162:18]
  reg [15:0] E_33; // @[SWChisel.scala 162:18]
  reg [15:0] E_34; // @[SWChisel.scala 162:18]
  reg [15:0] E_35; // @[SWChisel.scala 162:18]
  reg [15:0] E_36; // @[SWChisel.scala 162:18]
  reg [15:0] E_37; // @[SWChisel.scala 162:18]
  reg [15:0] E_38; // @[SWChisel.scala 162:18]
  reg [15:0] E_39; // @[SWChisel.scala 162:18]
  reg [15:0] F_1; // @[SWChisel.scala 163:18]
  reg [15:0] F_2; // @[SWChisel.scala 163:18]
  reg [15:0] F_3; // @[SWChisel.scala 163:18]
  reg [15:0] F_4; // @[SWChisel.scala 163:18]
  reg [15:0] F_5; // @[SWChisel.scala 163:18]
  reg [15:0] F_6; // @[SWChisel.scala 163:18]
  reg [15:0] F_7; // @[SWChisel.scala 163:18]
  reg [15:0] F_8; // @[SWChisel.scala 163:18]
  reg [15:0] F_9; // @[SWChisel.scala 163:18]
  reg [15:0] F_10; // @[SWChisel.scala 163:18]
  reg [15:0] F_11; // @[SWChisel.scala 163:18]
  reg [15:0] F_12; // @[SWChisel.scala 163:18]
  reg [15:0] F_13; // @[SWChisel.scala 163:18]
  reg [15:0] F_14; // @[SWChisel.scala 163:18]
  reg [15:0] F_15; // @[SWChisel.scala 163:18]
  reg [15:0] F_16; // @[SWChisel.scala 163:18]
  reg [15:0] F_17; // @[SWChisel.scala 163:18]
  reg [15:0] F_18; // @[SWChisel.scala 163:18]
  reg [15:0] F_19; // @[SWChisel.scala 163:18]
  reg [15:0] F_20; // @[SWChisel.scala 163:18]
  reg [15:0] F_21; // @[SWChisel.scala 163:18]
  reg [15:0] F_22; // @[SWChisel.scala 163:18]
  reg [15:0] F_23; // @[SWChisel.scala 163:18]
  reg [15:0] F_24; // @[SWChisel.scala 163:18]
  reg [15:0] F_25; // @[SWChisel.scala 163:18]
  reg [15:0] F_26; // @[SWChisel.scala 163:18]
  reg [15:0] F_27; // @[SWChisel.scala 163:18]
  reg [15:0] F_28; // @[SWChisel.scala 163:18]
  reg [15:0] F_29; // @[SWChisel.scala 163:18]
  reg [15:0] F_30; // @[SWChisel.scala 163:18]
  reg [15:0] F_31; // @[SWChisel.scala 163:18]
  reg [15:0] F_32; // @[SWChisel.scala 163:18]
  reg [15:0] F_33; // @[SWChisel.scala 163:18]
  reg [15:0] F_34; // @[SWChisel.scala 163:18]
  reg [15:0] F_35; // @[SWChisel.scala 163:18]
  reg [15:0] F_36; // @[SWChisel.scala 163:18]
  reg [15:0] F_37; // @[SWChisel.scala 163:18]
  reg [15:0] F_38; // @[SWChisel.scala 163:18]
  reg [15:0] F_39; // @[SWChisel.scala 163:18]
  reg [15:0] V1_0; // @[SWChisel.scala 164:19]
  reg [15:0] V1_1; // @[SWChisel.scala 164:19]
  reg [15:0] V1_2; // @[SWChisel.scala 164:19]
  reg [15:0] V1_3; // @[SWChisel.scala 164:19]
  reg [15:0] V1_4; // @[SWChisel.scala 164:19]
  reg [15:0] V1_5; // @[SWChisel.scala 164:19]
  reg [15:0] V1_6; // @[SWChisel.scala 164:19]
  reg [15:0] V1_7; // @[SWChisel.scala 164:19]
  reg [15:0] V1_8; // @[SWChisel.scala 164:19]
  reg [15:0] V1_9; // @[SWChisel.scala 164:19]
  reg [15:0] V1_10; // @[SWChisel.scala 164:19]
  reg [15:0] V1_11; // @[SWChisel.scala 164:19]
  reg [15:0] V1_12; // @[SWChisel.scala 164:19]
  reg [15:0] V1_13; // @[SWChisel.scala 164:19]
  reg [15:0] V1_14; // @[SWChisel.scala 164:19]
  reg [15:0] V1_15; // @[SWChisel.scala 164:19]
  reg [15:0] V1_16; // @[SWChisel.scala 164:19]
  reg [15:0] V1_17; // @[SWChisel.scala 164:19]
  reg [15:0] V1_18; // @[SWChisel.scala 164:19]
  reg [15:0] V1_19; // @[SWChisel.scala 164:19]
  reg [15:0] V1_20; // @[SWChisel.scala 164:19]
  reg [15:0] V1_21; // @[SWChisel.scala 164:19]
  reg [15:0] V1_22; // @[SWChisel.scala 164:19]
  reg [15:0] V1_23; // @[SWChisel.scala 164:19]
  reg [15:0] V1_24; // @[SWChisel.scala 164:19]
  reg [15:0] V1_25; // @[SWChisel.scala 164:19]
  reg [15:0] V1_26; // @[SWChisel.scala 164:19]
  reg [15:0] V1_27; // @[SWChisel.scala 164:19]
  reg [15:0] V1_28; // @[SWChisel.scala 164:19]
  reg [15:0] V1_29; // @[SWChisel.scala 164:19]
  reg [15:0] V1_30; // @[SWChisel.scala 164:19]
  reg [15:0] V1_31; // @[SWChisel.scala 164:19]
  reg [15:0] V1_32; // @[SWChisel.scala 164:19]
  reg [15:0] V1_33; // @[SWChisel.scala 164:19]
  reg [15:0] V1_34; // @[SWChisel.scala 164:19]
  reg [15:0] V1_35; // @[SWChisel.scala 164:19]
  reg [15:0] V1_36; // @[SWChisel.scala 164:19]
  reg [15:0] V1_37; // @[SWChisel.scala 164:19]
  reg [15:0] V1_38; // @[SWChisel.scala 164:19]
  reg [15:0] V1_39; // @[SWChisel.scala 164:19]
  reg [15:0] V1_40; // @[SWChisel.scala 164:19]
  reg [15:0] V2_0; // @[SWChisel.scala 166:19]
  reg [15:0] V2_1; // @[SWChisel.scala 166:19]
  reg [15:0] V2_2; // @[SWChisel.scala 166:19]
  reg [15:0] V2_3; // @[SWChisel.scala 166:19]
  reg [15:0] V2_4; // @[SWChisel.scala 166:19]
  reg [15:0] V2_5; // @[SWChisel.scala 166:19]
  reg [15:0] V2_6; // @[SWChisel.scala 166:19]
  reg [15:0] V2_7; // @[SWChisel.scala 166:19]
  reg [15:0] V2_8; // @[SWChisel.scala 166:19]
  reg [15:0] V2_9; // @[SWChisel.scala 166:19]
  reg [15:0] V2_10; // @[SWChisel.scala 166:19]
  reg [15:0] V2_11; // @[SWChisel.scala 166:19]
  reg [15:0] V2_12; // @[SWChisel.scala 166:19]
  reg [15:0] V2_13; // @[SWChisel.scala 166:19]
  reg [15:0] V2_14; // @[SWChisel.scala 166:19]
  reg [15:0] V2_15; // @[SWChisel.scala 166:19]
  reg [15:0] V2_16; // @[SWChisel.scala 166:19]
  reg [15:0] V2_17; // @[SWChisel.scala 166:19]
  reg [15:0] V2_18; // @[SWChisel.scala 166:19]
  reg [15:0] V2_19; // @[SWChisel.scala 166:19]
  reg [15:0] V2_20; // @[SWChisel.scala 166:19]
  reg [15:0] V2_21; // @[SWChisel.scala 166:19]
  reg [15:0] V2_22; // @[SWChisel.scala 166:19]
  reg [15:0] V2_23; // @[SWChisel.scala 166:19]
  reg [15:0] V2_24; // @[SWChisel.scala 166:19]
  reg [15:0] V2_25; // @[SWChisel.scala 166:19]
  reg [15:0] V2_26; // @[SWChisel.scala 166:19]
  reg [15:0] V2_27; // @[SWChisel.scala 166:19]
  reg [15:0] V2_28; // @[SWChisel.scala 166:19]
  reg [15:0] V2_29; // @[SWChisel.scala 166:19]
  reg [15:0] V2_30; // @[SWChisel.scala 166:19]
  reg [15:0] V2_31; // @[SWChisel.scala 166:19]
  reg [15:0] V2_32; // @[SWChisel.scala 166:19]
  reg [15:0] V2_33; // @[SWChisel.scala 166:19]
  reg [15:0] V2_34; // @[SWChisel.scala 166:19]
  reg [15:0] V2_35; // @[SWChisel.scala 166:19]
  reg [15:0] V2_36; // @[SWChisel.scala 166:19]
  reg [15:0] V2_37; // @[SWChisel.scala 166:19]
  reg [15:0] V2_38; // @[SWChisel.scala 166:19]
  reg [15:0] V2_39; // @[SWChisel.scala 166:19]
  reg  start_reg_0; // @[SWChisel.scala 167:26]
  reg  start_reg_1; // @[SWChisel.scala 167:26]
  reg  start_reg_2; // @[SWChisel.scala 167:26]
  reg  start_reg_3; // @[SWChisel.scala 167:26]
  reg  start_reg_4; // @[SWChisel.scala 167:26]
  reg  start_reg_5; // @[SWChisel.scala 167:26]
  reg  start_reg_6; // @[SWChisel.scala 167:26]
  reg  start_reg_7; // @[SWChisel.scala 167:26]
  reg  start_reg_8; // @[SWChisel.scala 167:26]
  reg  start_reg_9; // @[SWChisel.scala 167:26]
  reg  start_reg_10; // @[SWChisel.scala 167:26]
  reg  start_reg_11; // @[SWChisel.scala 167:26]
  reg  start_reg_12; // @[SWChisel.scala 167:26]
  reg  start_reg_13; // @[SWChisel.scala 167:26]
  reg  start_reg_14; // @[SWChisel.scala 167:26]
  reg  start_reg_15; // @[SWChisel.scala 167:26]
  reg  start_reg_16; // @[SWChisel.scala 167:26]
  reg  start_reg_17; // @[SWChisel.scala 167:26]
  reg  start_reg_18; // @[SWChisel.scala 167:26]
  reg  start_reg_19; // @[SWChisel.scala 167:26]
  reg  start_reg_20; // @[SWChisel.scala 167:26]
  reg  start_reg_21; // @[SWChisel.scala 167:26]
  reg  start_reg_22; // @[SWChisel.scala 167:26]
  reg  start_reg_23; // @[SWChisel.scala 167:26]
  reg  start_reg_24; // @[SWChisel.scala 167:26]
  reg  start_reg_25; // @[SWChisel.scala 167:26]
  reg  start_reg_26; // @[SWChisel.scala 167:26]
  reg  start_reg_27; // @[SWChisel.scala 167:26]
  reg  start_reg_28; // @[SWChisel.scala 167:26]
  reg  start_reg_29; // @[SWChisel.scala 167:26]
  reg  start_reg_30; // @[SWChisel.scala 167:26]
  reg  start_reg_31; // @[SWChisel.scala 167:26]
  reg  start_reg_32; // @[SWChisel.scala 167:26]
  reg  start_reg_33; // @[SWChisel.scala 167:26]
  reg  start_reg_34; // @[SWChisel.scala 167:26]
  reg  start_reg_35; // @[SWChisel.scala 167:26]
  reg  start_reg_36; // @[SWChisel.scala 167:26]
  reg  start_reg_37; // @[SWChisel.scala 167:26]
  reg  start_reg_38; // @[SWChisel.scala 167:26]
  reg  start_reg_39; // @[SWChisel.scala 167:26]
  wire [1:0] _GEN_121 = 8'h1 == r_count_0_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_122 = 8'h2 == r_count_0_io_out ? io_r_2_b : _GEN_121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_123 = 8'h3 == r_count_0_io_out ? io_r_3_b : _GEN_122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_124 = 8'h4 == r_count_0_io_out ? io_r_4_b : _GEN_123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_125 = 8'h5 == r_count_0_io_out ? io_r_5_b : _GEN_124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_126 = 8'h6 == r_count_0_io_out ? io_r_6_b : _GEN_125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_127 = 8'h7 == r_count_0_io_out ? io_r_7_b : _GEN_126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_128 = 8'h8 == r_count_0_io_out ? io_r_8_b : _GEN_127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_129 = 8'h9 == r_count_0_io_out ? io_r_9_b : _GEN_128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_130 = 8'ha == r_count_0_io_out ? io_r_10_b : _GEN_129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_131 = 8'hb == r_count_0_io_out ? io_r_11_b : _GEN_130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_132 = 8'hc == r_count_0_io_out ? io_r_12_b : _GEN_131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_133 = 8'hd == r_count_0_io_out ? io_r_13_b : _GEN_132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_134 = 8'he == r_count_0_io_out ? io_r_14_b : _GEN_133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_135 = 8'hf == r_count_0_io_out ? io_r_15_b : _GEN_134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_136 = 8'h10 == r_count_0_io_out ? io_r_16_b : _GEN_135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_137 = 8'h11 == r_count_0_io_out ? io_r_17_b : _GEN_136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_138 = 8'h12 == r_count_0_io_out ? io_r_18_b : _GEN_137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_139 = 8'h13 == r_count_0_io_out ? io_r_19_b : _GEN_138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_140 = 8'h14 == r_count_0_io_out ? io_r_20_b : _GEN_139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_141 = 8'h15 == r_count_0_io_out ? io_r_21_b : _GEN_140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_142 = 8'h16 == r_count_0_io_out ? io_r_22_b : _GEN_141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_143 = 8'h17 == r_count_0_io_out ? io_r_23_b : _GEN_142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_144 = 8'h18 == r_count_0_io_out ? io_r_24_b : _GEN_143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_145 = 8'h19 == r_count_0_io_out ? io_r_25_b : _GEN_144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_146 = 8'h1a == r_count_0_io_out ? io_r_26_b : _GEN_145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_147 = 8'h1b == r_count_0_io_out ? io_r_27_b : _GEN_146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_148 = 8'h1c == r_count_0_io_out ? io_r_28_b : _GEN_147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_149 = 8'h1d == r_count_0_io_out ? io_r_29_b : _GEN_148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_150 = 8'h1e == r_count_0_io_out ? io_r_30_b : _GEN_149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_151 = 8'h1f == r_count_0_io_out ? io_r_31_b : _GEN_150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_152 = 8'h20 == r_count_0_io_out ? io_r_32_b : _GEN_151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_153 = 8'h21 == r_count_0_io_out ? io_r_33_b : _GEN_152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_154 = 8'h22 == r_count_0_io_out ? io_r_34_b : _GEN_153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_155 = 8'h23 == r_count_0_io_out ? io_r_35_b : _GEN_154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_156 = 8'h24 == r_count_0_io_out ? io_r_36_b : _GEN_155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_157 = 8'h25 == r_count_0_io_out ? io_r_37_b : _GEN_156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_158 = 8'h26 == r_count_0_io_out ? io_r_38_b : _GEN_157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_159 = 8'h27 == r_count_0_io_out ? io_r_39_b : _GEN_158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_160 = 8'h28 == r_count_0_io_out ? io_r_40_b : _GEN_159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_161 = 8'h29 == r_count_0_io_out ? io_r_41_b : _GEN_160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_162 = 8'h2a == r_count_0_io_out ? io_r_42_b : _GEN_161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_163 = 8'h2b == r_count_0_io_out ? io_r_43_b : _GEN_162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_164 = 8'h2c == r_count_0_io_out ? io_r_44_b : _GEN_163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_165 = 8'h2d == r_count_0_io_out ? io_r_45_b : _GEN_164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_166 = 8'h2e == r_count_0_io_out ? io_r_46_b : _GEN_165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_167 = 8'h2f == r_count_0_io_out ? io_r_47_b : _GEN_166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_168 = 8'h30 == r_count_0_io_out ? io_r_48_b : _GEN_167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_169 = 8'h31 == r_count_0_io_out ? io_r_49_b : _GEN_168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_170 = 8'h32 == r_count_0_io_out ? io_r_50_b : _GEN_169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_171 = 8'h33 == r_count_0_io_out ? io_r_51_b : _GEN_170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_172 = 8'h34 == r_count_0_io_out ? io_r_52_b : _GEN_171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_173 = 8'h35 == r_count_0_io_out ? io_r_53_b : _GEN_172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_174 = 8'h36 == r_count_0_io_out ? io_r_54_b : _GEN_173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_175 = 8'h37 == r_count_0_io_out ? io_r_55_b : _GEN_174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_176 = 8'h38 == r_count_0_io_out ? io_r_56_b : _GEN_175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_177 = 8'h39 == r_count_0_io_out ? io_r_57_b : _GEN_176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_178 = 8'h3a == r_count_0_io_out ? io_r_58_b : _GEN_177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_179 = 8'h3b == r_count_0_io_out ? io_r_59_b : _GEN_178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_180 = 8'h3c == r_count_0_io_out ? io_r_60_b : _GEN_179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_181 = 8'h3d == r_count_0_io_out ? io_r_61_b : _GEN_180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_182 = 8'h3e == r_count_0_io_out ? io_r_62_b : _GEN_181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_183 = 8'h3f == r_count_0_io_out ? io_r_63_b : _GEN_182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_184 = 8'h40 == r_count_0_io_out ? io_r_64_b : _GEN_183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_185 = 8'h41 == r_count_0_io_out ? io_r_65_b : _GEN_184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_186 = 8'h42 == r_count_0_io_out ? io_r_66_b : _GEN_185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_187 = 8'h43 == r_count_0_io_out ? io_r_67_b : _GEN_186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_188 = 8'h44 == r_count_0_io_out ? io_r_68_b : _GEN_187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_189 = 8'h45 == r_count_0_io_out ? io_r_69_b : _GEN_188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_190 = 8'h46 == r_count_0_io_out ? io_r_70_b : _GEN_189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_191 = 8'h47 == r_count_0_io_out ? io_r_71_b : _GEN_190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_192 = 8'h48 == r_count_0_io_out ? io_r_72_b : _GEN_191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_193 = 8'h49 == r_count_0_io_out ? io_r_73_b : _GEN_192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_194 = 8'h4a == r_count_0_io_out ? io_r_74_b : _GEN_193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_195 = 8'h4b == r_count_0_io_out ? io_r_75_b : _GEN_194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_196 = 8'h4c == r_count_0_io_out ? io_r_76_b : _GEN_195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_197 = 8'h4d == r_count_0_io_out ? io_r_77_b : _GEN_196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_198 = 8'h4e == r_count_0_io_out ? io_r_78_b : _GEN_197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_199 = 8'h4f == r_count_0_io_out ? io_r_79_b : _GEN_198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_200 = 8'h50 == r_count_0_io_out ? io_r_80_b : _GEN_199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_201 = 8'h51 == r_count_0_io_out ? io_r_81_b : _GEN_200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_202 = 8'h52 == r_count_0_io_out ? io_r_82_b : _GEN_201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_203 = 8'h53 == r_count_0_io_out ? io_r_83_b : _GEN_202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_204 = 8'h54 == r_count_0_io_out ? io_r_84_b : _GEN_203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_205 = 8'h55 == r_count_0_io_out ? io_r_85_b : _GEN_204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_206 = 8'h56 == r_count_0_io_out ? io_r_86_b : _GEN_205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_207 = 8'h57 == r_count_0_io_out ? io_r_87_b : _GEN_206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_208 = 8'h58 == r_count_0_io_out ? io_r_88_b : _GEN_207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_209 = 8'h59 == r_count_0_io_out ? io_r_89_b : _GEN_208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_210 = 8'h5a == r_count_0_io_out ? io_r_90_b : _GEN_209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_211 = 8'h5b == r_count_0_io_out ? io_r_91_b : _GEN_210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_212 = 8'h5c == r_count_0_io_out ? io_r_92_b : _GEN_211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_213 = 8'h5d == r_count_0_io_out ? io_r_93_b : _GEN_212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_214 = 8'h5e == r_count_0_io_out ? io_r_94_b : _GEN_213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_215 = 8'h5f == r_count_0_io_out ? io_r_95_b : _GEN_214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_216 = 8'h60 == r_count_0_io_out ? io_r_96_b : _GEN_215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_217 = 8'h61 == r_count_0_io_out ? io_r_97_b : _GEN_216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_218 = 8'h62 == r_count_0_io_out ? io_r_98_b : _GEN_217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_219 = 8'h63 == r_count_0_io_out ? io_r_99_b : _GEN_218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_220 = 8'h64 == r_count_0_io_out ? io_r_100_b : _GEN_219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_221 = 8'h65 == r_count_0_io_out ? io_r_101_b : _GEN_220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_222 = 8'h66 == r_count_0_io_out ? io_r_102_b : _GEN_221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_223 = 8'h67 == r_count_0_io_out ? io_r_103_b : _GEN_222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_224 = 8'h68 == r_count_0_io_out ? io_r_104_b : _GEN_223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_225 = 8'h69 == r_count_0_io_out ? io_r_105_b : _GEN_224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_226 = 8'h6a == r_count_0_io_out ? io_r_106_b : _GEN_225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_227 = 8'h6b == r_count_0_io_out ? io_r_107_b : _GEN_226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_228 = 8'h6c == r_count_0_io_out ? io_r_108_b : _GEN_227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_229 = 8'h6d == r_count_0_io_out ? io_r_109_b : _GEN_228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_230 = 8'h6e == r_count_0_io_out ? io_r_110_b : _GEN_229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_231 = 8'h6f == r_count_0_io_out ? io_r_111_b : _GEN_230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_232 = 8'h70 == r_count_0_io_out ? io_r_112_b : _GEN_231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_233 = 8'h71 == r_count_0_io_out ? io_r_113_b : _GEN_232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_234 = 8'h72 == r_count_0_io_out ? io_r_114_b : _GEN_233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_235 = 8'h73 == r_count_0_io_out ? io_r_115_b : _GEN_234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_236 = 8'h74 == r_count_0_io_out ? io_r_116_b : _GEN_235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_237 = 8'h75 == r_count_0_io_out ? io_r_117_b : _GEN_236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_238 = 8'h76 == r_count_0_io_out ? io_r_118_b : _GEN_237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_239 = 8'h77 == r_count_0_io_out ? io_r_119_b : _GEN_238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_240 = 8'h78 == r_count_0_io_out ? io_r_120_b : _GEN_239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_241 = 8'h79 == r_count_0_io_out ? io_r_121_b : _GEN_240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_242 = 8'h7a == r_count_0_io_out ? io_r_122_b : _GEN_241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_243 = 8'h7b == r_count_0_io_out ? io_r_123_b : _GEN_242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_244 = 8'h7c == r_count_0_io_out ? io_r_124_b : _GEN_243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_245 = 8'h7d == r_count_0_io_out ? io_r_125_b : _GEN_244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_246 = 8'h7e == r_count_0_io_out ? io_r_126_b : _GEN_245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_247 = 8'h7f == r_count_0_io_out ? io_r_127_b : _GEN_246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_248 = 8'h80 == r_count_0_io_out ? io_r_128_b : _GEN_247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_249 = 8'h81 == r_count_0_io_out ? io_r_129_b : _GEN_248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_250 = 8'h82 == r_count_0_io_out ? io_r_130_b : _GEN_249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_251 = 8'h83 == r_count_0_io_out ? io_r_131_b : _GEN_250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_252 = 8'h84 == r_count_0_io_out ? io_r_132_b : _GEN_251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_253 = 8'h85 == r_count_0_io_out ? io_r_133_b : _GEN_252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_254 = 8'h86 == r_count_0_io_out ? io_r_134_b : _GEN_253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_255 = 8'h87 == r_count_0_io_out ? io_r_135_b : _GEN_254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_256 = 8'h88 == r_count_0_io_out ? io_r_136_b : _GEN_255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_257 = 8'h89 == r_count_0_io_out ? io_r_137_b : _GEN_256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_258 = 8'h8a == r_count_0_io_out ? io_r_138_b : _GEN_257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_259 = 8'h8b == r_count_0_io_out ? io_r_139_b : _GEN_258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_260 = 8'h8c == r_count_0_io_out ? io_r_140_b : _GEN_259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_261 = 8'h8d == r_count_0_io_out ? io_r_141_b : _GEN_260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_262 = 8'h8e == r_count_0_io_out ? io_r_142_b : _GEN_261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_263 = 8'h8f == r_count_0_io_out ? io_r_143_b : _GEN_262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_264 = 8'h90 == r_count_0_io_out ? io_r_144_b : _GEN_263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_265 = 8'h91 == r_count_0_io_out ? io_r_145_b : _GEN_264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_266 = 8'h92 == r_count_0_io_out ? io_r_146_b : _GEN_265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_267 = 8'h93 == r_count_0_io_out ? io_r_147_b : _GEN_266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_268 = 8'h94 == r_count_0_io_out ? io_r_148_b : _GEN_267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_269 = 8'h95 == r_count_0_io_out ? io_r_149_b : _GEN_268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_270 = 8'h96 == r_count_0_io_out ? io_r_150_b : _GEN_269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_271 = 8'h97 == r_count_0_io_out ? io_r_151_b : _GEN_270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_272 = 8'h98 == r_count_0_io_out ? io_r_152_b : _GEN_271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_273 = 8'h99 == r_count_0_io_out ? io_r_153_b : _GEN_272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_274 = 8'h9a == r_count_0_io_out ? io_r_154_b : _GEN_273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_275 = 8'h9b == r_count_0_io_out ? io_r_155_b : _GEN_274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_276 = 8'h9c == r_count_0_io_out ? io_r_156_b : _GEN_275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_277 = 8'h9d == r_count_0_io_out ? io_r_157_b : _GEN_276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_278 = 8'h9e == r_count_0_io_out ? io_r_158_b : _GEN_277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_279 = 8'h9f == r_count_0_io_out ? io_r_159_b : _GEN_278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_280 = 8'ha0 == r_count_0_io_out ? io_r_160_b : _GEN_279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_281 = 8'ha1 == r_count_0_io_out ? io_r_161_b : _GEN_280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_282 = 8'ha2 == r_count_0_io_out ? io_r_162_b : _GEN_281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_283 = 8'ha3 == r_count_0_io_out ? io_r_163_b : _GEN_282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_284 = 8'ha4 == r_count_0_io_out ? io_r_164_b : _GEN_283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_285 = 8'ha5 == r_count_0_io_out ? io_r_165_b : _GEN_284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_286 = 8'ha6 == r_count_0_io_out ? io_r_166_b : _GEN_285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_287 = 8'ha7 == r_count_0_io_out ? io_r_167_b : _GEN_286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_288 = 8'ha8 == r_count_0_io_out ? io_r_168_b : _GEN_287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_289 = 8'ha9 == r_count_0_io_out ? io_r_169_b : _GEN_288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_290 = 8'haa == r_count_0_io_out ? io_r_170_b : _GEN_289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_291 = 8'hab == r_count_0_io_out ? io_r_171_b : _GEN_290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_292 = 8'hac == r_count_0_io_out ? io_r_172_b : _GEN_291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_293 = 8'had == r_count_0_io_out ? io_r_173_b : _GEN_292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_294 = 8'hae == r_count_0_io_out ? io_r_174_b : _GEN_293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_295 = 8'haf == r_count_0_io_out ? io_r_175_b : _GEN_294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_296 = 8'hb0 == r_count_0_io_out ? io_r_176_b : _GEN_295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_297 = 8'hb1 == r_count_0_io_out ? io_r_177_b : _GEN_296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_298 = 8'hb2 == r_count_0_io_out ? io_r_178_b : _GEN_297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_299 = 8'hb3 == r_count_0_io_out ? io_r_179_b : _GEN_298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_300 = 8'hb4 == r_count_0_io_out ? io_r_180_b : _GEN_299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_301 = 8'hb5 == r_count_0_io_out ? io_r_181_b : _GEN_300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_302 = 8'hb6 == r_count_0_io_out ? io_r_182_b : _GEN_301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_303 = 8'hb7 == r_count_0_io_out ? io_r_183_b : _GEN_302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_304 = 8'hb8 == r_count_0_io_out ? io_r_184_b : _GEN_303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_305 = 8'hb9 == r_count_0_io_out ? io_r_185_b : _GEN_304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_306 = 8'hba == r_count_0_io_out ? io_r_186_b : _GEN_305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_307 = 8'hbb == r_count_0_io_out ? io_r_187_b : _GEN_306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_308 = 8'hbc == r_count_0_io_out ? io_r_188_b : _GEN_307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_309 = 8'hbd == r_count_0_io_out ? io_r_189_b : _GEN_308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_310 = 8'hbe == r_count_0_io_out ? io_r_190_b : _GEN_309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_311 = 8'hbf == r_count_0_io_out ? io_r_191_b : _GEN_310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_312 = 8'hc0 == r_count_0_io_out ? io_r_192_b : _GEN_311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_313 = 8'hc1 == r_count_0_io_out ? io_r_193_b : _GEN_312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_314 = 8'hc2 == r_count_0_io_out ? io_r_194_b : _GEN_313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_315 = 8'hc3 == r_count_0_io_out ? io_r_195_b : _GEN_314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_316 = 8'hc4 == r_count_0_io_out ? io_r_196_b : _GEN_315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_317 = 8'hc5 == r_count_0_io_out ? io_r_197_b : _GEN_316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_318 = 8'hc6 == r_count_0_io_out ? io_r_198_b : _GEN_317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_321 = 8'h1 == r_count_1_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_322 = 8'h2 == r_count_1_io_out ? io_r_2_b : _GEN_321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_323 = 8'h3 == r_count_1_io_out ? io_r_3_b : _GEN_322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_324 = 8'h4 == r_count_1_io_out ? io_r_4_b : _GEN_323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_325 = 8'h5 == r_count_1_io_out ? io_r_5_b : _GEN_324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_326 = 8'h6 == r_count_1_io_out ? io_r_6_b : _GEN_325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_327 = 8'h7 == r_count_1_io_out ? io_r_7_b : _GEN_326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_328 = 8'h8 == r_count_1_io_out ? io_r_8_b : _GEN_327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_329 = 8'h9 == r_count_1_io_out ? io_r_9_b : _GEN_328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_330 = 8'ha == r_count_1_io_out ? io_r_10_b : _GEN_329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_331 = 8'hb == r_count_1_io_out ? io_r_11_b : _GEN_330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_332 = 8'hc == r_count_1_io_out ? io_r_12_b : _GEN_331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_333 = 8'hd == r_count_1_io_out ? io_r_13_b : _GEN_332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_334 = 8'he == r_count_1_io_out ? io_r_14_b : _GEN_333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_335 = 8'hf == r_count_1_io_out ? io_r_15_b : _GEN_334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_336 = 8'h10 == r_count_1_io_out ? io_r_16_b : _GEN_335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_337 = 8'h11 == r_count_1_io_out ? io_r_17_b : _GEN_336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_338 = 8'h12 == r_count_1_io_out ? io_r_18_b : _GEN_337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_339 = 8'h13 == r_count_1_io_out ? io_r_19_b : _GEN_338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_340 = 8'h14 == r_count_1_io_out ? io_r_20_b : _GEN_339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_341 = 8'h15 == r_count_1_io_out ? io_r_21_b : _GEN_340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_342 = 8'h16 == r_count_1_io_out ? io_r_22_b : _GEN_341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_343 = 8'h17 == r_count_1_io_out ? io_r_23_b : _GEN_342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_344 = 8'h18 == r_count_1_io_out ? io_r_24_b : _GEN_343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_345 = 8'h19 == r_count_1_io_out ? io_r_25_b : _GEN_344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_346 = 8'h1a == r_count_1_io_out ? io_r_26_b : _GEN_345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_347 = 8'h1b == r_count_1_io_out ? io_r_27_b : _GEN_346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_348 = 8'h1c == r_count_1_io_out ? io_r_28_b : _GEN_347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_349 = 8'h1d == r_count_1_io_out ? io_r_29_b : _GEN_348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_350 = 8'h1e == r_count_1_io_out ? io_r_30_b : _GEN_349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_351 = 8'h1f == r_count_1_io_out ? io_r_31_b : _GEN_350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_352 = 8'h20 == r_count_1_io_out ? io_r_32_b : _GEN_351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_353 = 8'h21 == r_count_1_io_out ? io_r_33_b : _GEN_352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_354 = 8'h22 == r_count_1_io_out ? io_r_34_b : _GEN_353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_355 = 8'h23 == r_count_1_io_out ? io_r_35_b : _GEN_354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_356 = 8'h24 == r_count_1_io_out ? io_r_36_b : _GEN_355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_357 = 8'h25 == r_count_1_io_out ? io_r_37_b : _GEN_356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_358 = 8'h26 == r_count_1_io_out ? io_r_38_b : _GEN_357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_359 = 8'h27 == r_count_1_io_out ? io_r_39_b : _GEN_358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_360 = 8'h28 == r_count_1_io_out ? io_r_40_b : _GEN_359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_361 = 8'h29 == r_count_1_io_out ? io_r_41_b : _GEN_360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_362 = 8'h2a == r_count_1_io_out ? io_r_42_b : _GEN_361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_363 = 8'h2b == r_count_1_io_out ? io_r_43_b : _GEN_362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_364 = 8'h2c == r_count_1_io_out ? io_r_44_b : _GEN_363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_365 = 8'h2d == r_count_1_io_out ? io_r_45_b : _GEN_364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_366 = 8'h2e == r_count_1_io_out ? io_r_46_b : _GEN_365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_367 = 8'h2f == r_count_1_io_out ? io_r_47_b : _GEN_366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_368 = 8'h30 == r_count_1_io_out ? io_r_48_b : _GEN_367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_369 = 8'h31 == r_count_1_io_out ? io_r_49_b : _GEN_368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_370 = 8'h32 == r_count_1_io_out ? io_r_50_b : _GEN_369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_371 = 8'h33 == r_count_1_io_out ? io_r_51_b : _GEN_370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_372 = 8'h34 == r_count_1_io_out ? io_r_52_b : _GEN_371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_373 = 8'h35 == r_count_1_io_out ? io_r_53_b : _GEN_372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_374 = 8'h36 == r_count_1_io_out ? io_r_54_b : _GEN_373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_375 = 8'h37 == r_count_1_io_out ? io_r_55_b : _GEN_374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_376 = 8'h38 == r_count_1_io_out ? io_r_56_b : _GEN_375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_377 = 8'h39 == r_count_1_io_out ? io_r_57_b : _GEN_376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_378 = 8'h3a == r_count_1_io_out ? io_r_58_b : _GEN_377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_379 = 8'h3b == r_count_1_io_out ? io_r_59_b : _GEN_378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_380 = 8'h3c == r_count_1_io_out ? io_r_60_b : _GEN_379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_381 = 8'h3d == r_count_1_io_out ? io_r_61_b : _GEN_380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_382 = 8'h3e == r_count_1_io_out ? io_r_62_b : _GEN_381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_383 = 8'h3f == r_count_1_io_out ? io_r_63_b : _GEN_382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_384 = 8'h40 == r_count_1_io_out ? io_r_64_b : _GEN_383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_385 = 8'h41 == r_count_1_io_out ? io_r_65_b : _GEN_384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_386 = 8'h42 == r_count_1_io_out ? io_r_66_b : _GEN_385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_387 = 8'h43 == r_count_1_io_out ? io_r_67_b : _GEN_386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_388 = 8'h44 == r_count_1_io_out ? io_r_68_b : _GEN_387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_389 = 8'h45 == r_count_1_io_out ? io_r_69_b : _GEN_388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_390 = 8'h46 == r_count_1_io_out ? io_r_70_b : _GEN_389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_391 = 8'h47 == r_count_1_io_out ? io_r_71_b : _GEN_390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_392 = 8'h48 == r_count_1_io_out ? io_r_72_b : _GEN_391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_393 = 8'h49 == r_count_1_io_out ? io_r_73_b : _GEN_392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_394 = 8'h4a == r_count_1_io_out ? io_r_74_b : _GEN_393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_395 = 8'h4b == r_count_1_io_out ? io_r_75_b : _GEN_394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_396 = 8'h4c == r_count_1_io_out ? io_r_76_b : _GEN_395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_397 = 8'h4d == r_count_1_io_out ? io_r_77_b : _GEN_396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_398 = 8'h4e == r_count_1_io_out ? io_r_78_b : _GEN_397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_399 = 8'h4f == r_count_1_io_out ? io_r_79_b : _GEN_398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_400 = 8'h50 == r_count_1_io_out ? io_r_80_b : _GEN_399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_401 = 8'h51 == r_count_1_io_out ? io_r_81_b : _GEN_400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_402 = 8'h52 == r_count_1_io_out ? io_r_82_b : _GEN_401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_403 = 8'h53 == r_count_1_io_out ? io_r_83_b : _GEN_402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_404 = 8'h54 == r_count_1_io_out ? io_r_84_b : _GEN_403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_405 = 8'h55 == r_count_1_io_out ? io_r_85_b : _GEN_404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_406 = 8'h56 == r_count_1_io_out ? io_r_86_b : _GEN_405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_407 = 8'h57 == r_count_1_io_out ? io_r_87_b : _GEN_406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_408 = 8'h58 == r_count_1_io_out ? io_r_88_b : _GEN_407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_409 = 8'h59 == r_count_1_io_out ? io_r_89_b : _GEN_408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_410 = 8'h5a == r_count_1_io_out ? io_r_90_b : _GEN_409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_411 = 8'h5b == r_count_1_io_out ? io_r_91_b : _GEN_410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_412 = 8'h5c == r_count_1_io_out ? io_r_92_b : _GEN_411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_413 = 8'h5d == r_count_1_io_out ? io_r_93_b : _GEN_412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_414 = 8'h5e == r_count_1_io_out ? io_r_94_b : _GEN_413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_415 = 8'h5f == r_count_1_io_out ? io_r_95_b : _GEN_414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_416 = 8'h60 == r_count_1_io_out ? io_r_96_b : _GEN_415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_417 = 8'h61 == r_count_1_io_out ? io_r_97_b : _GEN_416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_418 = 8'h62 == r_count_1_io_out ? io_r_98_b : _GEN_417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_419 = 8'h63 == r_count_1_io_out ? io_r_99_b : _GEN_418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_420 = 8'h64 == r_count_1_io_out ? io_r_100_b : _GEN_419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_421 = 8'h65 == r_count_1_io_out ? io_r_101_b : _GEN_420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_422 = 8'h66 == r_count_1_io_out ? io_r_102_b : _GEN_421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_423 = 8'h67 == r_count_1_io_out ? io_r_103_b : _GEN_422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_424 = 8'h68 == r_count_1_io_out ? io_r_104_b : _GEN_423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_425 = 8'h69 == r_count_1_io_out ? io_r_105_b : _GEN_424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_426 = 8'h6a == r_count_1_io_out ? io_r_106_b : _GEN_425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_427 = 8'h6b == r_count_1_io_out ? io_r_107_b : _GEN_426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_428 = 8'h6c == r_count_1_io_out ? io_r_108_b : _GEN_427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_429 = 8'h6d == r_count_1_io_out ? io_r_109_b : _GEN_428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_430 = 8'h6e == r_count_1_io_out ? io_r_110_b : _GEN_429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_431 = 8'h6f == r_count_1_io_out ? io_r_111_b : _GEN_430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_432 = 8'h70 == r_count_1_io_out ? io_r_112_b : _GEN_431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_433 = 8'h71 == r_count_1_io_out ? io_r_113_b : _GEN_432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_434 = 8'h72 == r_count_1_io_out ? io_r_114_b : _GEN_433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_435 = 8'h73 == r_count_1_io_out ? io_r_115_b : _GEN_434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_436 = 8'h74 == r_count_1_io_out ? io_r_116_b : _GEN_435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_437 = 8'h75 == r_count_1_io_out ? io_r_117_b : _GEN_436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_438 = 8'h76 == r_count_1_io_out ? io_r_118_b : _GEN_437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_439 = 8'h77 == r_count_1_io_out ? io_r_119_b : _GEN_438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_440 = 8'h78 == r_count_1_io_out ? io_r_120_b : _GEN_439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_441 = 8'h79 == r_count_1_io_out ? io_r_121_b : _GEN_440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_442 = 8'h7a == r_count_1_io_out ? io_r_122_b : _GEN_441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_443 = 8'h7b == r_count_1_io_out ? io_r_123_b : _GEN_442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_444 = 8'h7c == r_count_1_io_out ? io_r_124_b : _GEN_443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_445 = 8'h7d == r_count_1_io_out ? io_r_125_b : _GEN_444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_446 = 8'h7e == r_count_1_io_out ? io_r_126_b : _GEN_445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_447 = 8'h7f == r_count_1_io_out ? io_r_127_b : _GEN_446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_448 = 8'h80 == r_count_1_io_out ? io_r_128_b : _GEN_447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_449 = 8'h81 == r_count_1_io_out ? io_r_129_b : _GEN_448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_450 = 8'h82 == r_count_1_io_out ? io_r_130_b : _GEN_449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_451 = 8'h83 == r_count_1_io_out ? io_r_131_b : _GEN_450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_452 = 8'h84 == r_count_1_io_out ? io_r_132_b : _GEN_451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_453 = 8'h85 == r_count_1_io_out ? io_r_133_b : _GEN_452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_454 = 8'h86 == r_count_1_io_out ? io_r_134_b : _GEN_453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_455 = 8'h87 == r_count_1_io_out ? io_r_135_b : _GEN_454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_456 = 8'h88 == r_count_1_io_out ? io_r_136_b : _GEN_455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_457 = 8'h89 == r_count_1_io_out ? io_r_137_b : _GEN_456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_458 = 8'h8a == r_count_1_io_out ? io_r_138_b : _GEN_457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_459 = 8'h8b == r_count_1_io_out ? io_r_139_b : _GEN_458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_460 = 8'h8c == r_count_1_io_out ? io_r_140_b : _GEN_459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_461 = 8'h8d == r_count_1_io_out ? io_r_141_b : _GEN_460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_462 = 8'h8e == r_count_1_io_out ? io_r_142_b : _GEN_461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_463 = 8'h8f == r_count_1_io_out ? io_r_143_b : _GEN_462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_464 = 8'h90 == r_count_1_io_out ? io_r_144_b : _GEN_463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_465 = 8'h91 == r_count_1_io_out ? io_r_145_b : _GEN_464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_466 = 8'h92 == r_count_1_io_out ? io_r_146_b : _GEN_465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_467 = 8'h93 == r_count_1_io_out ? io_r_147_b : _GEN_466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_468 = 8'h94 == r_count_1_io_out ? io_r_148_b : _GEN_467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_469 = 8'h95 == r_count_1_io_out ? io_r_149_b : _GEN_468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_470 = 8'h96 == r_count_1_io_out ? io_r_150_b : _GEN_469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_471 = 8'h97 == r_count_1_io_out ? io_r_151_b : _GEN_470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_472 = 8'h98 == r_count_1_io_out ? io_r_152_b : _GEN_471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_473 = 8'h99 == r_count_1_io_out ? io_r_153_b : _GEN_472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_474 = 8'h9a == r_count_1_io_out ? io_r_154_b : _GEN_473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_475 = 8'h9b == r_count_1_io_out ? io_r_155_b : _GEN_474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_476 = 8'h9c == r_count_1_io_out ? io_r_156_b : _GEN_475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_477 = 8'h9d == r_count_1_io_out ? io_r_157_b : _GEN_476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_478 = 8'h9e == r_count_1_io_out ? io_r_158_b : _GEN_477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_479 = 8'h9f == r_count_1_io_out ? io_r_159_b : _GEN_478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_480 = 8'ha0 == r_count_1_io_out ? io_r_160_b : _GEN_479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_481 = 8'ha1 == r_count_1_io_out ? io_r_161_b : _GEN_480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_482 = 8'ha2 == r_count_1_io_out ? io_r_162_b : _GEN_481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_483 = 8'ha3 == r_count_1_io_out ? io_r_163_b : _GEN_482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_484 = 8'ha4 == r_count_1_io_out ? io_r_164_b : _GEN_483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_485 = 8'ha5 == r_count_1_io_out ? io_r_165_b : _GEN_484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_486 = 8'ha6 == r_count_1_io_out ? io_r_166_b : _GEN_485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_487 = 8'ha7 == r_count_1_io_out ? io_r_167_b : _GEN_486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_488 = 8'ha8 == r_count_1_io_out ? io_r_168_b : _GEN_487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_489 = 8'ha9 == r_count_1_io_out ? io_r_169_b : _GEN_488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_490 = 8'haa == r_count_1_io_out ? io_r_170_b : _GEN_489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_491 = 8'hab == r_count_1_io_out ? io_r_171_b : _GEN_490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_492 = 8'hac == r_count_1_io_out ? io_r_172_b : _GEN_491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_493 = 8'had == r_count_1_io_out ? io_r_173_b : _GEN_492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_494 = 8'hae == r_count_1_io_out ? io_r_174_b : _GEN_493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_495 = 8'haf == r_count_1_io_out ? io_r_175_b : _GEN_494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_496 = 8'hb0 == r_count_1_io_out ? io_r_176_b : _GEN_495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_497 = 8'hb1 == r_count_1_io_out ? io_r_177_b : _GEN_496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_498 = 8'hb2 == r_count_1_io_out ? io_r_178_b : _GEN_497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_499 = 8'hb3 == r_count_1_io_out ? io_r_179_b : _GEN_498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_500 = 8'hb4 == r_count_1_io_out ? io_r_180_b : _GEN_499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_501 = 8'hb5 == r_count_1_io_out ? io_r_181_b : _GEN_500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_502 = 8'hb6 == r_count_1_io_out ? io_r_182_b : _GEN_501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_503 = 8'hb7 == r_count_1_io_out ? io_r_183_b : _GEN_502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_504 = 8'hb8 == r_count_1_io_out ? io_r_184_b : _GEN_503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_505 = 8'hb9 == r_count_1_io_out ? io_r_185_b : _GEN_504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_506 = 8'hba == r_count_1_io_out ? io_r_186_b : _GEN_505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_507 = 8'hbb == r_count_1_io_out ? io_r_187_b : _GEN_506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_508 = 8'hbc == r_count_1_io_out ? io_r_188_b : _GEN_507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_509 = 8'hbd == r_count_1_io_out ? io_r_189_b : _GEN_508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_510 = 8'hbe == r_count_1_io_out ? io_r_190_b : _GEN_509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_511 = 8'hbf == r_count_1_io_out ? io_r_191_b : _GEN_510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_512 = 8'hc0 == r_count_1_io_out ? io_r_192_b : _GEN_511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_513 = 8'hc1 == r_count_1_io_out ? io_r_193_b : _GEN_512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_514 = 8'hc2 == r_count_1_io_out ? io_r_194_b : _GEN_513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_515 = 8'hc3 == r_count_1_io_out ? io_r_195_b : _GEN_514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_516 = 8'hc4 == r_count_1_io_out ? io_r_196_b : _GEN_515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_517 = 8'hc5 == r_count_1_io_out ? io_r_197_b : _GEN_516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_518 = 8'hc6 == r_count_1_io_out ? io_r_198_b : _GEN_517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_521 = 8'h1 == r_count_2_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_522 = 8'h2 == r_count_2_io_out ? io_r_2_b : _GEN_521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_523 = 8'h3 == r_count_2_io_out ? io_r_3_b : _GEN_522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_524 = 8'h4 == r_count_2_io_out ? io_r_4_b : _GEN_523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_525 = 8'h5 == r_count_2_io_out ? io_r_5_b : _GEN_524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_526 = 8'h6 == r_count_2_io_out ? io_r_6_b : _GEN_525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_527 = 8'h7 == r_count_2_io_out ? io_r_7_b : _GEN_526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_528 = 8'h8 == r_count_2_io_out ? io_r_8_b : _GEN_527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_529 = 8'h9 == r_count_2_io_out ? io_r_9_b : _GEN_528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_530 = 8'ha == r_count_2_io_out ? io_r_10_b : _GEN_529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_531 = 8'hb == r_count_2_io_out ? io_r_11_b : _GEN_530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_532 = 8'hc == r_count_2_io_out ? io_r_12_b : _GEN_531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_533 = 8'hd == r_count_2_io_out ? io_r_13_b : _GEN_532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_534 = 8'he == r_count_2_io_out ? io_r_14_b : _GEN_533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_535 = 8'hf == r_count_2_io_out ? io_r_15_b : _GEN_534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_536 = 8'h10 == r_count_2_io_out ? io_r_16_b : _GEN_535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_537 = 8'h11 == r_count_2_io_out ? io_r_17_b : _GEN_536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_538 = 8'h12 == r_count_2_io_out ? io_r_18_b : _GEN_537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_539 = 8'h13 == r_count_2_io_out ? io_r_19_b : _GEN_538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_540 = 8'h14 == r_count_2_io_out ? io_r_20_b : _GEN_539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_541 = 8'h15 == r_count_2_io_out ? io_r_21_b : _GEN_540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_542 = 8'h16 == r_count_2_io_out ? io_r_22_b : _GEN_541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_543 = 8'h17 == r_count_2_io_out ? io_r_23_b : _GEN_542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_544 = 8'h18 == r_count_2_io_out ? io_r_24_b : _GEN_543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_545 = 8'h19 == r_count_2_io_out ? io_r_25_b : _GEN_544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_546 = 8'h1a == r_count_2_io_out ? io_r_26_b : _GEN_545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_547 = 8'h1b == r_count_2_io_out ? io_r_27_b : _GEN_546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_548 = 8'h1c == r_count_2_io_out ? io_r_28_b : _GEN_547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_549 = 8'h1d == r_count_2_io_out ? io_r_29_b : _GEN_548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_550 = 8'h1e == r_count_2_io_out ? io_r_30_b : _GEN_549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_551 = 8'h1f == r_count_2_io_out ? io_r_31_b : _GEN_550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_552 = 8'h20 == r_count_2_io_out ? io_r_32_b : _GEN_551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_553 = 8'h21 == r_count_2_io_out ? io_r_33_b : _GEN_552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_554 = 8'h22 == r_count_2_io_out ? io_r_34_b : _GEN_553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_555 = 8'h23 == r_count_2_io_out ? io_r_35_b : _GEN_554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_556 = 8'h24 == r_count_2_io_out ? io_r_36_b : _GEN_555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_557 = 8'h25 == r_count_2_io_out ? io_r_37_b : _GEN_556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_558 = 8'h26 == r_count_2_io_out ? io_r_38_b : _GEN_557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_559 = 8'h27 == r_count_2_io_out ? io_r_39_b : _GEN_558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_560 = 8'h28 == r_count_2_io_out ? io_r_40_b : _GEN_559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_561 = 8'h29 == r_count_2_io_out ? io_r_41_b : _GEN_560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_562 = 8'h2a == r_count_2_io_out ? io_r_42_b : _GEN_561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_563 = 8'h2b == r_count_2_io_out ? io_r_43_b : _GEN_562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_564 = 8'h2c == r_count_2_io_out ? io_r_44_b : _GEN_563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_565 = 8'h2d == r_count_2_io_out ? io_r_45_b : _GEN_564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_566 = 8'h2e == r_count_2_io_out ? io_r_46_b : _GEN_565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_567 = 8'h2f == r_count_2_io_out ? io_r_47_b : _GEN_566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_568 = 8'h30 == r_count_2_io_out ? io_r_48_b : _GEN_567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_569 = 8'h31 == r_count_2_io_out ? io_r_49_b : _GEN_568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_570 = 8'h32 == r_count_2_io_out ? io_r_50_b : _GEN_569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_571 = 8'h33 == r_count_2_io_out ? io_r_51_b : _GEN_570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_572 = 8'h34 == r_count_2_io_out ? io_r_52_b : _GEN_571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_573 = 8'h35 == r_count_2_io_out ? io_r_53_b : _GEN_572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_574 = 8'h36 == r_count_2_io_out ? io_r_54_b : _GEN_573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_575 = 8'h37 == r_count_2_io_out ? io_r_55_b : _GEN_574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_576 = 8'h38 == r_count_2_io_out ? io_r_56_b : _GEN_575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_577 = 8'h39 == r_count_2_io_out ? io_r_57_b : _GEN_576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_578 = 8'h3a == r_count_2_io_out ? io_r_58_b : _GEN_577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_579 = 8'h3b == r_count_2_io_out ? io_r_59_b : _GEN_578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_580 = 8'h3c == r_count_2_io_out ? io_r_60_b : _GEN_579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_581 = 8'h3d == r_count_2_io_out ? io_r_61_b : _GEN_580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_582 = 8'h3e == r_count_2_io_out ? io_r_62_b : _GEN_581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_583 = 8'h3f == r_count_2_io_out ? io_r_63_b : _GEN_582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_584 = 8'h40 == r_count_2_io_out ? io_r_64_b : _GEN_583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_585 = 8'h41 == r_count_2_io_out ? io_r_65_b : _GEN_584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_586 = 8'h42 == r_count_2_io_out ? io_r_66_b : _GEN_585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_587 = 8'h43 == r_count_2_io_out ? io_r_67_b : _GEN_586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_588 = 8'h44 == r_count_2_io_out ? io_r_68_b : _GEN_587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_589 = 8'h45 == r_count_2_io_out ? io_r_69_b : _GEN_588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_590 = 8'h46 == r_count_2_io_out ? io_r_70_b : _GEN_589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_591 = 8'h47 == r_count_2_io_out ? io_r_71_b : _GEN_590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_592 = 8'h48 == r_count_2_io_out ? io_r_72_b : _GEN_591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_593 = 8'h49 == r_count_2_io_out ? io_r_73_b : _GEN_592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_594 = 8'h4a == r_count_2_io_out ? io_r_74_b : _GEN_593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_595 = 8'h4b == r_count_2_io_out ? io_r_75_b : _GEN_594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_596 = 8'h4c == r_count_2_io_out ? io_r_76_b : _GEN_595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_597 = 8'h4d == r_count_2_io_out ? io_r_77_b : _GEN_596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_598 = 8'h4e == r_count_2_io_out ? io_r_78_b : _GEN_597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_599 = 8'h4f == r_count_2_io_out ? io_r_79_b : _GEN_598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_600 = 8'h50 == r_count_2_io_out ? io_r_80_b : _GEN_599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_601 = 8'h51 == r_count_2_io_out ? io_r_81_b : _GEN_600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_602 = 8'h52 == r_count_2_io_out ? io_r_82_b : _GEN_601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_603 = 8'h53 == r_count_2_io_out ? io_r_83_b : _GEN_602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_604 = 8'h54 == r_count_2_io_out ? io_r_84_b : _GEN_603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_605 = 8'h55 == r_count_2_io_out ? io_r_85_b : _GEN_604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_606 = 8'h56 == r_count_2_io_out ? io_r_86_b : _GEN_605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_607 = 8'h57 == r_count_2_io_out ? io_r_87_b : _GEN_606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_608 = 8'h58 == r_count_2_io_out ? io_r_88_b : _GEN_607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_609 = 8'h59 == r_count_2_io_out ? io_r_89_b : _GEN_608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_610 = 8'h5a == r_count_2_io_out ? io_r_90_b : _GEN_609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_611 = 8'h5b == r_count_2_io_out ? io_r_91_b : _GEN_610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_612 = 8'h5c == r_count_2_io_out ? io_r_92_b : _GEN_611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_613 = 8'h5d == r_count_2_io_out ? io_r_93_b : _GEN_612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_614 = 8'h5e == r_count_2_io_out ? io_r_94_b : _GEN_613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_615 = 8'h5f == r_count_2_io_out ? io_r_95_b : _GEN_614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_616 = 8'h60 == r_count_2_io_out ? io_r_96_b : _GEN_615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_617 = 8'h61 == r_count_2_io_out ? io_r_97_b : _GEN_616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_618 = 8'h62 == r_count_2_io_out ? io_r_98_b : _GEN_617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_619 = 8'h63 == r_count_2_io_out ? io_r_99_b : _GEN_618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_620 = 8'h64 == r_count_2_io_out ? io_r_100_b : _GEN_619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_621 = 8'h65 == r_count_2_io_out ? io_r_101_b : _GEN_620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_622 = 8'h66 == r_count_2_io_out ? io_r_102_b : _GEN_621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_623 = 8'h67 == r_count_2_io_out ? io_r_103_b : _GEN_622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_624 = 8'h68 == r_count_2_io_out ? io_r_104_b : _GEN_623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_625 = 8'h69 == r_count_2_io_out ? io_r_105_b : _GEN_624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_626 = 8'h6a == r_count_2_io_out ? io_r_106_b : _GEN_625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_627 = 8'h6b == r_count_2_io_out ? io_r_107_b : _GEN_626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_628 = 8'h6c == r_count_2_io_out ? io_r_108_b : _GEN_627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_629 = 8'h6d == r_count_2_io_out ? io_r_109_b : _GEN_628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_630 = 8'h6e == r_count_2_io_out ? io_r_110_b : _GEN_629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_631 = 8'h6f == r_count_2_io_out ? io_r_111_b : _GEN_630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_632 = 8'h70 == r_count_2_io_out ? io_r_112_b : _GEN_631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_633 = 8'h71 == r_count_2_io_out ? io_r_113_b : _GEN_632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_634 = 8'h72 == r_count_2_io_out ? io_r_114_b : _GEN_633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_635 = 8'h73 == r_count_2_io_out ? io_r_115_b : _GEN_634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_636 = 8'h74 == r_count_2_io_out ? io_r_116_b : _GEN_635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_637 = 8'h75 == r_count_2_io_out ? io_r_117_b : _GEN_636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_638 = 8'h76 == r_count_2_io_out ? io_r_118_b : _GEN_637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_639 = 8'h77 == r_count_2_io_out ? io_r_119_b : _GEN_638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_640 = 8'h78 == r_count_2_io_out ? io_r_120_b : _GEN_639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_641 = 8'h79 == r_count_2_io_out ? io_r_121_b : _GEN_640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_642 = 8'h7a == r_count_2_io_out ? io_r_122_b : _GEN_641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_643 = 8'h7b == r_count_2_io_out ? io_r_123_b : _GEN_642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_644 = 8'h7c == r_count_2_io_out ? io_r_124_b : _GEN_643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_645 = 8'h7d == r_count_2_io_out ? io_r_125_b : _GEN_644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_646 = 8'h7e == r_count_2_io_out ? io_r_126_b : _GEN_645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_647 = 8'h7f == r_count_2_io_out ? io_r_127_b : _GEN_646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_648 = 8'h80 == r_count_2_io_out ? io_r_128_b : _GEN_647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_649 = 8'h81 == r_count_2_io_out ? io_r_129_b : _GEN_648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_650 = 8'h82 == r_count_2_io_out ? io_r_130_b : _GEN_649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_651 = 8'h83 == r_count_2_io_out ? io_r_131_b : _GEN_650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_652 = 8'h84 == r_count_2_io_out ? io_r_132_b : _GEN_651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_653 = 8'h85 == r_count_2_io_out ? io_r_133_b : _GEN_652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_654 = 8'h86 == r_count_2_io_out ? io_r_134_b : _GEN_653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_655 = 8'h87 == r_count_2_io_out ? io_r_135_b : _GEN_654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_656 = 8'h88 == r_count_2_io_out ? io_r_136_b : _GEN_655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_657 = 8'h89 == r_count_2_io_out ? io_r_137_b : _GEN_656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_658 = 8'h8a == r_count_2_io_out ? io_r_138_b : _GEN_657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_659 = 8'h8b == r_count_2_io_out ? io_r_139_b : _GEN_658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_660 = 8'h8c == r_count_2_io_out ? io_r_140_b : _GEN_659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_661 = 8'h8d == r_count_2_io_out ? io_r_141_b : _GEN_660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_662 = 8'h8e == r_count_2_io_out ? io_r_142_b : _GEN_661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_663 = 8'h8f == r_count_2_io_out ? io_r_143_b : _GEN_662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_664 = 8'h90 == r_count_2_io_out ? io_r_144_b : _GEN_663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_665 = 8'h91 == r_count_2_io_out ? io_r_145_b : _GEN_664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_666 = 8'h92 == r_count_2_io_out ? io_r_146_b : _GEN_665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_667 = 8'h93 == r_count_2_io_out ? io_r_147_b : _GEN_666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_668 = 8'h94 == r_count_2_io_out ? io_r_148_b : _GEN_667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_669 = 8'h95 == r_count_2_io_out ? io_r_149_b : _GEN_668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_670 = 8'h96 == r_count_2_io_out ? io_r_150_b : _GEN_669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_671 = 8'h97 == r_count_2_io_out ? io_r_151_b : _GEN_670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_672 = 8'h98 == r_count_2_io_out ? io_r_152_b : _GEN_671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_673 = 8'h99 == r_count_2_io_out ? io_r_153_b : _GEN_672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_674 = 8'h9a == r_count_2_io_out ? io_r_154_b : _GEN_673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_675 = 8'h9b == r_count_2_io_out ? io_r_155_b : _GEN_674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_676 = 8'h9c == r_count_2_io_out ? io_r_156_b : _GEN_675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_677 = 8'h9d == r_count_2_io_out ? io_r_157_b : _GEN_676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_678 = 8'h9e == r_count_2_io_out ? io_r_158_b : _GEN_677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_679 = 8'h9f == r_count_2_io_out ? io_r_159_b : _GEN_678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_680 = 8'ha0 == r_count_2_io_out ? io_r_160_b : _GEN_679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_681 = 8'ha1 == r_count_2_io_out ? io_r_161_b : _GEN_680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_682 = 8'ha2 == r_count_2_io_out ? io_r_162_b : _GEN_681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_683 = 8'ha3 == r_count_2_io_out ? io_r_163_b : _GEN_682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_684 = 8'ha4 == r_count_2_io_out ? io_r_164_b : _GEN_683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_685 = 8'ha5 == r_count_2_io_out ? io_r_165_b : _GEN_684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_686 = 8'ha6 == r_count_2_io_out ? io_r_166_b : _GEN_685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_687 = 8'ha7 == r_count_2_io_out ? io_r_167_b : _GEN_686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_688 = 8'ha8 == r_count_2_io_out ? io_r_168_b : _GEN_687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_689 = 8'ha9 == r_count_2_io_out ? io_r_169_b : _GEN_688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_690 = 8'haa == r_count_2_io_out ? io_r_170_b : _GEN_689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_691 = 8'hab == r_count_2_io_out ? io_r_171_b : _GEN_690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_692 = 8'hac == r_count_2_io_out ? io_r_172_b : _GEN_691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_693 = 8'had == r_count_2_io_out ? io_r_173_b : _GEN_692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_694 = 8'hae == r_count_2_io_out ? io_r_174_b : _GEN_693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_695 = 8'haf == r_count_2_io_out ? io_r_175_b : _GEN_694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_696 = 8'hb0 == r_count_2_io_out ? io_r_176_b : _GEN_695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_697 = 8'hb1 == r_count_2_io_out ? io_r_177_b : _GEN_696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_698 = 8'hb2 == r_count_2_io_out ? io_r_178_b : _GEN_697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_699 = 8'hb3 == r_count_2_io_out ? io_r_179_b : _GEN_698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_700 = 8'hb4 == r_count_2_io_out ? io_r_180_b : _GEN_699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_701 = 8'hb5 == r_count_2_io_out ? io_r_181_b : _GEN_700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_702 = 8'hb6 == r_count_2_io_out ? io_r_182_b : _GEN_701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_703 = 8'hb7 == r_count_2_io_out ? io_r_183_b : _GEN_702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_704 = 8'hb8 == r_count_2_io_out ? io_r_184_b : _GEN_703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_705 = 8'hb9 == r_count_2_io_out ? io_r_185_b : _GEN_704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_706 = 8'hba == r_count_2_io_out ? io_r_186_b : _GEN_705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_707 = 8'hbb == r_count_2_io_out ? io_r_187_b : _GEN_706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_708 = 8'hbc == r_count_2_io_out ? io_r_188_b : _GEN_707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_709 = 8'hbd == r_count_2_io_out ? io_r_189_b : _GEN_708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_710 = 8'hbe == r_count_2_io_out ? io_r_190_b : _GEN_709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_711 = 8'hbf == r_count_2_io_out ? io_r_191_b : _GEN_710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_712 = 8'hc0 == r_count_2_io_out ? io_r_192_b : _GEN_711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_713 = 8'hc1 == r_count_2_io_out ? io_r_193_b : _GEN_712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_714 = 8'hc2 == r_count_2_io_out ? io_r_194_b : _GEN_713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_715 = 8'hc3 == r_count_2_io_out ? io_r_195_b : _GEN_714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_716 = 8'hc4 == r_count_2_io_out ? io_r_196_b : _GEN_715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_717 = 8'hc5 == r_count_2_io_out ? io_r_197_b : _GEN_716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_718 = 8'hc6 == r_count_2_io_out ? io_r_198_b : _GEN_717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_721 = 8'h1 == r_count_3_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_722 = 8'h2 == r_count_3_io_out ? io_r_2_b : _GEN_721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_723 = 8'h3 == r_count_3_io_out ? io_r_3_b : _GEN_722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_724 = 8'h4 == r_count_3_io_out ? io_r_4_b : _GEN_723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_725 = 8'h5 == r_count_3_io_out ? io_r_5_b : _GEN_724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_726 = 8'h6 == r_count_3_io_out ? io_r_6_b : _GEN_725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_727 = 8'h7 == r_count_3_io_out ? io_r_7_b : _GEN_726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_728 = 8'h8 == r_count_3_io_out ? io_r_8_b : _GEN_727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_729 = 8'h9 == r_count_3_io_out ? io_r_9_b : _GEN_728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_730 = 8'ha == r_count_3_io_out ? io_r_10_b : _GEN_729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_731 = 8'hb == r_count_3_io_out ? io_r_11_b : _GEN_730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_732 = 8'hc == r_count_3_io_out ? io_r_12_b : _GEN_731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_733 = 8'hd == r_count_3_io_out ? io_r_13_b : _GEN_732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_734 = 8'he == r_count_3_io_out ? io_r_14_b : _GEN_733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_735 = 8'hf == r_count_3_io_out ? io_r_15_b : _GEN_734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_736 = 8'h10 == r_count_3_io_out ? io_r_16_b : _GEN_735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_737 = 8'h11 == r_count_3_io_out ? io_r_17_b : _GEN_736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_738 = 8'h12 == r_count_3_io_out ? io_r_18_b : _GEN_737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_739 = 8'h13 == r_count_3_io_out ? io_r_19_b : _GEN_738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_740 = 8'h14 == r_count_3_io_out ? io_r_20_b : _GEN_739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_741 = 8'h15 == r_count_3_io_out ? io_r_21_b : _GEN_740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_742 = 8'h16 == r_count_3_io_out ? io_r_22_b : _GEN_741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_743 = 8'h17 == r_count_3_io_out ? io_r_23_b : _GEN_742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_744 = 8'h18 == r_count_3_io_out ? io_r_24_b : _GEN_743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_745 = 8'h19 == r_count_3_io_out ? io_r_25_b : _GEN_744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_746 = 8'h1a == r_count_3_io_out ? io_r_26_b : _GEN_745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_747 = 8'h1b == r_count_3_io_out ? io_r_27_b : _GEN_746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_748 = 8'h1c == r_count_3_io_out ? io_r_28_b : _GEN_747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_749 = 8'h1d == r_count_3_io_out ? io_r_29_b : _GEN_748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_750 = 8'h1e == r_count_3_io_out ? io_r_30_b : _GEN_749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_751 = 8'h1f == r_count_3_io_out ? io_r_31_b : _GEN_750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_752 = 8'h20 == r_count_3_io_out ? io_r_32_b : _GEN_751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_753 = 8'h21 == r_count_3_io_out ? io_r_33_b : _GEN_752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_754 = 8'h22 == r_count_3_io_out ? io_r_34_b : _GEN_753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_755 = 8'h23 == r_count_3_io_out ? io_r_35_b : _GEN_754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_756 = 8'h24 == r_count_3_io_out ? io_r_36_b : _GEN_755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_757 = 8'h25 == r_count_3_io_out ? io_r_37_b : _GEN_756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_758 = 8'h26 == r_count_3_io_out ? io_r_38_b : _GEN_757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_759 = 8'h27 == r_count_3_io_out ? io_r_39_b : _GEN_758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_760 = 8'h28 == r_count_3_io_out ? io_r_40_b : _GEN_759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_761 = 8'h29 == r_count_3_io_out ? io_r_41_b : _GEN_760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_762 = 8'h2a == r_count_3_io_out ? io_r_42_b : _GEN_761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_763 = 8'h2b == r_count_3_io_out ? io_r_43_b : _GEN_762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_764 = 8'h2c == r_count_3_io_out ? io_r_44_b : _GEN_763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_765 = 8'h2d == r_count_3_io_out ? io_r_45_b : _GEN_764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_766 = 8'h2e == r_count_3_io_out ? io_r_46_b : _GEN_765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_767 = 8'h2f == r_count_3_io_out ? io_r_47_b : _GEN_766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_768 = 8'h30 == r_count_3_io_out ? io_r_48_b : _GEN_767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_769 = 8'h31 == r_count_3_io_out ? io_r_49_b : _GEN_768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_770 = 8'h32 == r_count_3_io_out ? io_r_50_b : _GEN_769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_771 = 8'h33 == r_count_3_io_out ? io_r_51_b : _GEN_770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_772 = 8'h34 == r_count_3_io_out ? io_r_52_b : _GEN_771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_773 = 8'h35 == r_count_3_io_out ? io_r_53_b : _GEN_772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_774 = 8'h36 == r_count_3_io_out ? io_r_54_b : _GEN_773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_775 = 8'h37 == r_count_3_io_out ? io_r_55_b : _GEN_774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_776 = 8'h38 == r_count_3_io_out ? io_r_56_b : _GEN_775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_777 = 8'h39 == r_count_3_io_out ? io_r_57_b : _GEN_776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_778 = 8'h3a == r_count_3_io_out ? io_r_58_b : _GEN_777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_779 = 8'h3b == r_count_3_io_out ? io_r_59_b : _GEN_778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_780 = 8'h3c == r_count_3_io_out ? io_r_60_b : _GEN_779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_781 = 8'h3d == r_count_3_io_out ? io_r_61_b : _GEN_780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_782 = 8'h3e == r_count_3_io_out ? io_r_62_b : _GEN_781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_783 = 8'h3f == r_count_3_io_out ? io_r_63_b : _GEN_782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_784 = 8'h40 == r_count_3_io_out ? io_r_64_b : _GEN_783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_785 = 8'h41 == r_count_3_io_out ? io_r_65_b : _GEN_784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_786 = 8'h42 == r_count_3_io_out ? io_r_66_b : _GEN_785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_787 = 8'h43 == r_count_3_io_out ? io_r_67_b : _GEN_786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_788 = 8'h44 == r_count_3_io_out ? io_r_68_b : _GEN_787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_789 = 8'h45 == r_count_3_io_out ? io_r_69_b : _GEN_788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_790 = 8'h46 == r_count_3_io_out ? io_r_70_b : _GEN_789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_791 = 8'h47 == r_count_3_io_out ? io_r_71_b : _GEN_790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_792 = 8'h48 == r_count_3_io_out ? io_r_72_b : _GEN_791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_793 = 8'h49 == r_count_3_io_out ? io_r_73_b : _GEN_792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_794 = 8'h4a == r_count_3_io_out ? io_r_74_b : _GEN_793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_795 = 8'h4b == r_count_3_io_out ? io_r_75_b : _GEN_794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_796 = 8'h4c == r_count_3_io_out ? io_r_76_b : _GEN_795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_797 = 8'h4d == r_count_3_io_out ? io_r_77_b : _GEN_796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_798 = 8'h4e == r_count_3_io_out ? io_r_78_b : _GEN_797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_799 = 8'h4f == r_count_3_io_out ? io_r_79_b : _GEN_798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_800 = 8'h50 == r_count_3_io_out ? io_r_80_b : _GEN_799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_801 = 8'h51 == r_count_3_io_out ? io_r_81_b : _GEN_800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_802 = 8'h52 == r_count_3_io_out ? io_r_82_b : _GEN_801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_803 = 8'h53 == r_count_3_io_out ? io_r_83_b : _GEN_802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_804 = 8'h54 == r_count_3_io_out ? io_r_84_b : _GEN_803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_805 = 8'h55 == r_count_3_io_out ? io_r_85_b : _GEN_804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_806 = 8'h56 == r_count_3_io_out ? io_r_86_b : _GEN_805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_807 = 8'h57 == r_count_3_io_out ? io_r_87_b : _GEN_806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_808 = 8'h58 == r_count_3_io_out ? io_r_88_b : _GEN_807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_809 = 8'h59 == r_count_3_io_out ? io_r_89_b : _GEN_808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_810 = 8'h5a == r_count_3_io_out ? io_r_90_b : _GEN_809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_811 = 8'h5b == r_count_3_io_out ? io_r_91_b : _GEN_810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_812 = 8'h5c == r_count_3_io_out ? io_r_92_b : _GEN_811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_813 = 8'h5d == r_count_3_io_out ? io_r_93_b : _GEN_812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_814 = 8'h5e == r_count_3_io_out ? io_r_94_b : _GEN_813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_815 = 8'h5f == r_count_3_io_out ? io_r_95_b : _GEN_814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_816 = 8'h60 == r_count_3_io_out ? io_r_96_b : _GEN_815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_817 = 8'h61 == r_count_3_io_out ? io_r_97_b : _GEN_816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_818 = 8'h62 == r_count_3_io_out ? io_r_98_b : _GEN_817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_819 = 8'h63 == r_count_3_io_out ? io_r_99_b : _GEN_818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_820 = 8'h64 == r_count_3_io_out ? io_r_100_b : _GEN_819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_821 = 8'h65 == r_count_3_io_out ? io_r_101_b : _GEN_820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_822 = 8'h66 == r_count_3_io_out ? io_r_102_b : _GEN_821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_823 = 8'h67 == r_count_3_io_out ? io_r_103_b : _GEN_822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_824 = 8'h68 == r_count_3_io_out ? io_r_104_b : _GEN_823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_825 = 8'h69 == r_count_3_io_out ? io_r_105_b : _GEN_824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_826 = 8'h6a == r_count_3_io_out ? io_r_106_b : _GEN_825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_827 = 8'h6b == r_count_3_io_out ? io_r_107_b : _GEN_826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_828 = 8'h6c == r_count_3_io_out ? io_r_108_b : _GEN_827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_829 = 8'h6d == r_count_3_io_out ? io_r_109_b : _GEN_828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_830 = 8'h6e == r_count_3_io_out ? io_r_110_b : _GEN_829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_831 = 8'h6f == r_count_3_io_out ? io_r_111_b : _GEN_830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_832 = 8'h70 == r_count_3_io_out ? io_r_112_b : _GEN_831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_833 = 8'h71 == r_count_3_io_out ? io_r_113_b : _GEN_832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_834 = 8'h72 == r_count_3_io_out ? io_r_114_b : _GEN_833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_835 = 8'h73 == r_count_3_io_out ? io_r_115_b : _GEN_834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_836 = 8'h74 == r_count_3_io_out ? io_r_116_b : _GEN_835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_837 = 8'h75 == r_count_3_io_out ? io_r_117_b : _GEN_836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_838 = 8'h76 == r_count_3_io_out ? io_r_118_b : _GEN_837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_839 = 8'h77 == r_count_3_io_out ? io_r_119_b : _GEN_838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_840 = 8'h78 == r_count_3_io_out ? io_r_120_b : _GEN_839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_841 = 8'h79 == r_count_3_io_out ? io_r_121_b : _GEN_840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_842 = 8'h7a == r_count_3_io_out ? io_r_122_b : _GEN_841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_843 = 8'h7b == r_count_3_io_out ? io_r_123_b : _GEN_842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_844 = 8'h7c == r_count_3_io_out ? io_r_124_b : _GEN_843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_845 = 8'h7d == r_count_3_io_out ? io_r_125_b : _GEN_844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_846 = 8'h7e == r_count_3_io_out ? io_r_126_b : _GEN_845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_847 = 8'h7f == r_count_3_io_out ? io_r_127_b : _GEN_846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_848 = 8'h80 == r_count_3_io_out ? io_r_128_b : _GEN_847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_849 = 8'h81 == r_count_3_io_out ? io_r_129_b : _GEN_848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_850 = 8'h82 == r_count_3_io_out ? io_r_130_b : _GEN_849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_851 = 8'h83 == r_count_3_io_out ? io_r_131_b : _GEN_850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_852 = 8'h84 == r_count_3_io_out ? io_r_132_b : _GEN_851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_853 = 8'h85 == r_count_3_io_out ? io_r_133_b : _GEN_852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_854 = 8'h86 == r_count_3_io_out ? io_r_134_b : _GEN_853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_855 = 8'h87 == r_count_3_io_out ? io_r_135_b : _GEN_854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_856 = 8'h88 == r_count_3_io_out ? io_r_136_b : _GEN_855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_857 = 8'h89 == r_count_3_io_out ? io_r_137_b : _GEN_856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_858 = 8'h8a == r_count_3_io_out ? io_r_138_b : _GEN_857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_859 = 8'h8b == r_count_3_io_out ? io_r_139_b : _GEN_858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_860 = 8'h8c == r_count_3_io_out ? io_r_140_b : _GEN_859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_861 = 8'h8d == r_count_3_io_out ? io_r_141_b : _GEN_860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_862 = 8'h8e == r_count_3_io_out ? io_r_142_b : _GEN_861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_863 = 8'h8f == r_count_3_io_out ? io_r_143_b : _GEN_862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_864 = 8'h90 == r_count_3_io_out ? io_r_144_b : _GEN_863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_865 = 8'h91 == r_count_3_io_out ? io_r_145_b : _GEN_864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_866 = 8'h92 == r_count_3_io_out ? io_r_146_b : _GEN_865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_867 = 8'h93 == r_count_3_io_out ? io_r_147_b : _GEN_866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_868 = 8'h94 == r_count_3_io_out ? io_r_148_b : _GEN_867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_869 = 8'h95 == r_count_3_io_out ? io_r_149_b : _GEN_868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_870 = 8'h96 == r_count_3_io_out ? io_r_150_b : _GEN_869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_871 = 8'h97 == r_count_3_io_out ? io_r_151_b : _GEN_870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_872 = 8'h98 == r_count_3_io_out ? io_r_152_b : _GEN_871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_873 = 8'h99 == r_count_3_io_out ? io_r_153_b : _GEN_872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_874 = 8'h9a == r_count_3_io_out ? io_r_154_b : _GEN_873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_875 = 8'h9b == r_count_3_io_out ? io_r_155_b : _GEN_874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_876 = 8'h9c == r_count_3_io_out ? io_r_156_b : _GEN_875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_877 = 8'h9d == r_count_3_io_out ? io_r_157_b : _GEN_876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_878 = 8'h9e == r_count_3_io_out ? io_r_158_b : _GEN_877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_879 = 8'h9f == r_count_3_io_out ? io_r_159_b : _GEN_878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_880 = 8'ha0 == r_count_3_io_out ? io_r_160_b : _GEN_879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_881 = 8'ha1 == r_count_3_io_out ? io_r_161_b : _GEN_880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_882 = 8'ha2 == r_count_3_io_out ? io_r_162_b : _GEN_881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_883 = 8'ha3 == r_count_3_io_out ? io_r_163_b : _GEN_882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_884 = 8'ha4 == r_count_3_io_out ? io_r_164_b : _GEN_883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_885 = 8'ha5 == r_count_3_io_out ? io_r_165_b : _GEN_884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_886 = 8'ha6 == r_count_3_io_out ? io_r_166_b : _GEN_885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_887 = 8'ha7 == r_count_3_io_out ? io_r_167_b : _GEN_886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_888 = 8'ha8 == r_count_3_io_out ? io_r_168_b : _GEN_887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_889 = 8'ha9 == r_count_3_io_out ? io_r_169_b : _GEN_888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_890 = 8'haa == r_count_3_io_out ? io_r_170_b : _GEN_889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_891 = 8'hab == r_count_3_io_out ? io_r_171_b : _GEN_890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_892 = 8'hac == r_count_3_io_out ? io_r_172_b : _GEN_891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_893 = 8'had == r_count_3_io_out ? io_r_173_b : _GEN_892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_894 = 8'hae == r_count_3_io_out ? io_r_174_b : _GEN_893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_895 = 8'haf == r_count_3_io_out ? io_r_175_b : _GEN_894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_896 = 8'hb0 == r_count_3_io_out ? io_r_176_b : _GEN_895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_897 = 8'hb1 == r_count_3_io_out ? io_r_177_b : _GEN_896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_898 = 8'hb2 == r_count_3_io_out ? io_r_178_b : _GEN_897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_899 = 8'hb3 == r_count_3_io_out ? io_r_179_b : _GEN_898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_900 = 8'hb4 == r_count_3_io_out ? io_r_180_b : _GEN_899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_901 = 8'hb5 == r_count_3_io_out ? io_r_181_b : _GEN_900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_902 = 8'hb6 == r_count_3_io_out ? io_r_182_b : _GEN_901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_903 = 8'hb7 == r_count_3_io_out ? io_r_183_b : _GEN_902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_904 = 8'hb8 == r_count_3_io_out ? io_r_184_b : _GEN_903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_905 = 8'hb9 == r_count_3_io_out ? io_r_185_b : _GEN_904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_906 = 8'hba == r_count_3_io_out ? io_r_186_b : _GEN_905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_907 = 8'hbb == r_count_3_io_out ? io_r_187_b : _GEN_906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_908 = 8'hbc == r_count_3_io_out ? io_r_188_b : _GEN_907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_909 = 8'hbd == r_count_3_io_out ? io_r_189_b : _GEN_908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_910 = 8'hbe == r_count_3_io_out ? io_r_190_b : _GEN_909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_911 = 8'hbf == r_count_3_io_out ? io_r_191_b : _GEN_910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_912 = 8'hc0 == r_count_3_io_out ? io_r_192_b : _GEN_911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_913 = 8'hc1 == r_count_3_io_out ? io_r_193_b : _GEN_912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_914 = 8'hc2 == r_count_3_io_out ? io_r_194_b : _GEN_913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_915 = 8'hc3 == r_count_3_io_out ? io_r_195_b : _GEN_914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_916 = 8'hc4 == r_count_3_io_out ? io_r_196_b : _GEN_915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_917 = 8'hc5 == r_count_3_io_out ? io_r_197_b : _GEN_916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_918 = 8'hc6 == r_count_3_io_out ? io_r_198_b : _GEN_917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_921 = 8'h1 == r_count_4_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_922 = 8'h2 == r_count_4_io_out ? io_r_2_b : _GEN_921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_923 = 8'h3 == r_count_4_io_out ? io_r_3_b : _GEN_922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_924 = 8'h4 == r_count_4_io_out ? io_r_4_b : _GEN_923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_925 = 8'h5 == r_count_4_io_out ? io_r_5_b : _GEN_924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_926 = 8'h6 == r_count_4_io_out ? io_r_6_b : _GEN_925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_927 = 8'h7 == r_count_4_io_out ? io_r_7_b : _GEN_926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_928 = 8'h8 == r_count_4_io_out ? io_r_8_b : _GEN_927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_929 = 8'h9 == r_count_4_io_out ? io_r_9_b : _GEN_928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_930 = 8'ha == r_count_4_io_out ? io_r_10_b : _GEN_929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_931 = 8'hb == r_count_4_io_out ? io_r_11_b : _GEN_930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_932 = 8'hc == r_count_4_io_out ? io_r_12_b : _GEN_931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_933 = 8'hd == r_count_4_io_out ? io_r_13_b : _GEN_932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_934 = 8'he == r_count_4_io_out ? io_r_14_b : _GEN_933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_935 = 8'hf == r_count_4_io_out ? io_r_15_b : _GEN_934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_936 = 8'h10 == r_count_4_io_out ? io_r_16_b : _GEN_935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_937 = 8'h11 == r_count_4_io_out ? io_r_17_b : _GEN_936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_938 = 8'h12 == r_count_4_io_out ? io_r_18_b : _GEN_937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_939 = 8'h13 == r_count_4_io_out ? io_r_19_b : _GEN_938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_940 = 8'h14 == r_count_4_io_out ? io_r_20_b : _GEN_939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_941 = 8'h15 == r_count_4_io_out ? io_r_21_b : _GEN_940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_942 = 8'h16 == r_count_4_io_out ? io_r_22_b : _GEN_941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_943 = 8'h17 == r_count_4_io_out ? io_r_23_b : _GEN_942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_944 = 8'h18 == r_count_4_io_out ? io_r_24_b : _GEN_943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_945 = 8'h19 == r_count_4_io_out ? io_r_25_b : _GEN_944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_946 = 8'h1a == r_count_4_io_out ? io_r_26_b : _GEN_945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_947 = 8'h1b == r_count_4_io_out ? io_r_27_b : _GEN_946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_948 = 8'h1c == r_count_4_io_out ? io_r_28_b : _GEN_947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_949 = 8'h1d == r_count_4_io_out ? io_r_29_b : _GEN_948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_950 = 8'h1e == r_count_4_io_out ? io_r_30_b : _GEN_949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_951 = 8'h1f == r_count_4_io_out ? io_r_31_b : _GEN_950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_952 = 8'h20 == r_count_4_io_out ? io_r_32_b : _GEN_951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_953 = 8'h21 == r_count_4_io_out ? io_r_33_b : _GEN_952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_954 = 8'h22 == r_count_4_io_out ? io_r_34_b : _GEN_953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_955 = 8'h23 == r_count_4_io_out ? io_r_35_b : _GEN_954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_956 = 8'h24 == r_count_4_io_out ? io_r_36_b : _GEN_955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_957 = 8'h25 == r_count_4_io_out ? io_r_37_b : _GEN_956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_958 = 8'h26 == r_count_4_io_out ? io_r_38_b : _GEN_957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_959 = 8'h27 == r_count_4_io_out ? io_r_39_b : _GEN_958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_960 = 8'h28 == r_count_4_io_out ? io_r_40_b : _GEN_959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_961 = 8'h29 == r_count_4_io_out ? io_r_41_b : _GEN_960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_962 = 8'h2a == r_count_4_io_out ? io_r_42_b : _GEN_961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_963 = 8'h2b == r_count_4_io_out ? io_r_43_b : _GEN_962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_964 = 8'h2c == r_count_4_io_out ? io_r_44_b : _GEN_963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_965 = 8'h2d == r_count_4_io_out ? io_r_45_b : _GEN_964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_966 = 8'h2e == r_count_4_io_out ? io_r_46_b : _GEN_965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_967 = 8'h2f == r_count_4_io_out ? io_r_47_b : _GEN_966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_968 = 8'h30 == r_count_4_io_out ? io_r_48_b : _GEN_967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_969 = 8'h31 == r_count_4_io_out ? io_r_49_b : _GEN_968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_970 = 8'h32 == r_count_4_io_out ? io_r_50_b : _GEN_969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_971 = 8'h33 == r_count_4_io_out ? io_r_51_b : _GEN_970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_972 = 8'h34 == r_count_4_io_out ? io_r_52_b : _GEN_971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_973 = 8'h35 == r_count_4_io_out ? io_r_53_b : _GEN_972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_974 = 8'h36 == r_count_4_io_out ? io_r_54_b : _GEN_973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_975 = 8'h37 == r_count_4_io_out ? io_r_55_b : _GEN_974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_976 = 8'h38 == r_count_4_io_out ? io_r_56_b : _GEN_975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_977 = 8'h39 == r_count_4_io_out ? io_r_57_b : _GEN_976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_978 = 8'h3a == r_count_4_io_out ? io_r_58_b : _GEN_977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_979 = 8'h3b == r_count_4_io_out ? io_r_59_b : _GEN_978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_980 = 8'h3c == r_count_4_io_out ? io_r_60_b : _GEN_979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_981 = 8'h3d == r_count_4_io_out ? io_r_61_b : _GEN_980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_982 = 8'h3e == r_count_4_io_out ? io_r_62_b : _GEN_981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_983 = 8'h3f == r_count_4_io_out ? io_r_63_b : _GEN_982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_984 = 8'h40 == r_count_4_io_out ? io_r_64_b : _GEN_983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_985 = 8'h41 == r_count_4_io_out ? io_r_65_b : _GEN_984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_986 = 8'h42 == r_count_4_io_out ? io_r_66_b : _GEN_985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_987 = 8'h43 == r_count_4_io_out ? io_r_67_b : _GEN_986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_988 = 8'h44 == r_count_4_io_out ? io_r_68_b : _GEN_987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_989 = 8'h45 == r_count_4_io_out ? io_r_69_b : _GEN_988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_990 = 8'h46 == r_count_4_io_out ? io_r_70_b : _GEN_989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_991 = 8'h47 == r_count_4_io_out ? io_r_71_b : _GEN_990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_992 = 8'h48 == r_count_4_io_out ? io_r_72_b : _GEN_991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_993 = 8'h49 == r_count_4_io_out ? io_r_73_b : _GEN_992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_994 = 8'h4a == r_count_4_io_out ? io_r_74_b : _GEN_993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_995 = 8'h4b == r_count_4_io_out ? io_r_75_b : _GEN_994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_996 = 8'h4c == r_count_4_io_out ? io_r_76_b : _GEN_995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_997 = 8'h4d == r_count_4_io_out ? io_r_77_b : _GEN_996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_998 = 8'h4e == r_count_4_io_out ? io_r_78_b : _GEN_997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_999 = 8'h4f == r_count_4_io_out ? io_r_79_b : _GEN_998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1000 = 8'h50 == r_count_4_io_out ? io_r_80_b : _GEN_999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1001 = 8'h51 == r_count_4_io_out ? io_r_81_b : _GEN_1000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1002 = 8'h52 == r_count_4_io_out ? io_r_82_b : _GEN_1001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1003 = 8'h53 == r_count_4_io_out ? io_r_83_b : _GEN_1002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1004 = 8'h54 == r_count_4_io_out ? io_r_84_b : _GEN_1003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1005 = 8'h55 == r_count_4_io_out ? io_r_85_b : _GEN_1004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1006 = 8'h56 == r_count_4_io_out ? io_r_86_b : _GEN_1005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1007 = 8'h57 == r_count_4_io_out ? io_r_87_b : _GEN_1006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1008 = 8'h58 == r_count_4_io_out ? io_r_88_b : _GEN_1007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1009 = 8'h59 == r_count_4_io_out ? io_r_89_b : _GEN_1008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1010 = 8'h5a == r_count_4_io_out ? io_r_90_b : _GEN_1009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1011 = 8'h5b == r_count_4_io_out ? io_r_91_b : _GEN_1010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1012 = 8'h5c == r_count_4_io_out ? io_r_92_b : _GEN_1011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1013 = 8'h5d == r_count_4_io_out ? io_r_93_b : _GEN_1012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1014 = 8'h5e == r_count_4_io_out ? io_r_94_b : _GEN_1013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1015 = 8'h5f == r_count_4_io_out ? io_r_95_b : _GEN_1014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1016 = 8'h60 == r_count_4_io_out ? io_r_96_b : _GEN_1015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1017 = 8'h61 == r_count_4_io_out ? io_r_97_b : _GEN_1016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1018 = 8'h62 == r_count_4_io_out ? io_r_98_b : _GEN_1017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1019 = 8'h63 == r_count_4_io_out ? io_r_99_b : _GEN_1018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1020 = 8'h64 == r_count_4_io_out ? io_r_100_b : _GEN_1019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1021 = 8'h65 == r_count_4_io_out ? io_r_101_b : _GEN_1020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1022 = 8'h66 == r_count_4_io_out ? io_r_102_b : _GEN_1021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1023 = 8'h67 == r_count_4_io_out ? io_r_103_b : _GEN_1022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1024 = 8'h68 == r_count_4_io_out ? io_r_104_b : _GEN_1023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1025 = 8'h69 == r_count_4_io_out ? io_r_105_b : _GEN_1024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1026 = 8'h6a == r_count_4_io_out ? io_r_106_b : _GEN_1025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1027 = 8'h6b == r_count_4_io_out ? io_r_107_b : _GEN_1026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1028 = 8'h6c == r_count_4_io_out ? io_r_108_b : _GEN_1027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1029 = 8'h6d == r_count_4_io_out ? io_r_109_b : _GEN_1028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1030 = 8'h6e == r_count_4_io_out ? io_r_110_b : _GEN_1029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1031 = 8'h6f == r_count_4_io_out ? io_r_111_b : _GEN_1030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1032 = 8'h70 == r_count_4_io_out ? io_r_112_b : _GEN_1031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1033 = 8'h71 == r_count_4_io_out ? io_r_113_b : _GEN_1032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1034 = 8'h72 == r_count_4_io_out ? io_r_114_b : _GEN_1033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1035 = 8'h73 == r_count_4_io_out ? io_r_115_b : _GEN_1034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1036 = 8'h74 == r_count_4_io_out ? io_r_116_b : _GEN_1035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1037 = 8'h75 == r_count_4_io_out ? io_r_117_b : _GEN_1036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1038 = 8'h76 == r_count_4_io_out ? io_r_118_b : _GEN_1037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1039 = 8'h77 == r_count_4_io_out ? io_r_119_b : _GEN_1038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1040 = 8'h78 == r_count_4_io_out ? io_r_120_b : _GEN_1039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1041 = 8'h79 == r_count_4_io_out ? io_r_121_b : _GEN_1040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1042 = 8'h7a == r_count_4_io_out ? io_r_122_b : _GEN_1041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1043 = 8'h7b == r_count_4_io_out ? io_r_123_b : _GEN_1042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1044 = 8'h7c == r_count_4_io_out ? io_r_124_b : _GEN_1043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1045 = 8'h7d == r_count_4_io_out ? io_r_125_b : _GEN_1044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1046 = 8'h7e == r_count_4_io_out ? io_r_126_b : _GEN_1045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1047 = 8'h7f == r_count_4_io_out ? io_r_127_b : _GEN_1046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1048 = 8'h80 == r_count_4_io_out ? io_r_128_b : _GEN_1047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1049 = 8'h81 == r_count_4_io_out ? io_r_129_b : _GEN_1048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1050 = 8'h82 == r_count_4_io_out ? io_r_130_b : _GEN_1049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1051 = 8'h83 == r_count_4_io_out ? io_r_131_b : _GEN_1050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1052 = 8'h84 == r_count_4_io_out ? io_r_132_b : _GEN_1051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1053 = 8'h85 == r_count_4_io_out ? io_r_133_b : _GEN_1052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1054 = 8'h86 == r_count_4_io_out ? io_r_134_b : _GEN_1053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1055 = 8'h87 == r_count_4_io_out ? io_r_135_b : _GEN_1054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1056 = 8'h88 == r_count_4_io_out ? io_r_136_b : _GEN_1055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1057 = 8'h89 == r_count_4_io_out ? io_r_137_b : _GEN_1056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1058 = 8'h8a == r_count_4_io_out ? io_r_138_b : _GEN_1057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1059 = 8'h8b == r_count_4_io_out ? io_r_139_b : _GEN_1058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1060 = 8'h8c == r_count_4_io_out ? io_r_140_b : _GEN_1059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1061 = 8'h8d == r_count_4_io_out ? io_r_141_b : _GEN_1060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1062 = 8'h8e == r_count_4_io_out ? io_r_142_b : _GEN_1061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1063 = 8'h8f == r_count_4_io_out ? io_r_143_b : _GEN_1062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1064 = 8'h90 == r_count_4_io_out ? io_r_144_b : _GEN_1063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1065 = 8'h91 == r_count_4_io_out ? io_r_145_b : _GEN_1064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1066 = 8'h92 == r_count_4_io_out ? io_r_146_b : _GEN_1065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1067 = 8'h93 == r_count_4_io_out ? io_r_147_b : _GEN_1066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1068 = 8'h94 == r_count_4_io_out ? io_r_148_b : _GEN_1067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1069 = 8'h95 == r_count_4_io_out ? io_r_149_b : _GEN_1068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1070 = 8'h96 == r_count_4_io_out ? io_r_150_b : _GEN_1069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1071 = 8'h97 == r_count_4_io_out ? io_r_151_b : _GEN_1070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1072 = 8'h98 == r_count_4_io_out ? io_r_152_b : _GEN_1071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1073 = 8'h99 == r_count_4_io_out ? io_r_153_b : _GEN_1072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1074 = 8'h9a == r_count_4_io_out ? io_r_154_b : _GEN_1073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1075 = 8'h9b == r_count_4_io_out ? io_r_155_b : _GEN_1074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1076 = 8'h9c == r_count_4_io_out ? io_r_156_b : _GEN_1075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1077 = 8'h9d == r_count_4_io_out ? io_r_157_b : _GEN_1076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1078 = 8'h9e == r_count_4_io_out ? io_r_158_b : _GEN_1077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1079 = 8'h9f == r_count_4_io_out ? io_r_159_b : _GEN_1078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1080 = 8'ha0 == r_count_4_io_out ? io_r_160_b : _GEN_1079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1081 = 8'ha1 == r_count_4_io_out ? io_r_161_b : _GEN_1080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1082 = 8'ha2 == r_count_4_io_out ? io_r_162_b : _GEN_1081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1083 = 8'ha3 == r_count_4_io_out ? io_r_163_b : _GEN_1082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1084 = 8'ha4 == r_count_4_io_out ? io_r_164_b : _GEN_1083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1085 = 8'ha5 == r_count_4_io_out ? io_r_165_b : _GEN_1084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1086 = 8'ha6 == r_count_4_io_out ? io_r_166_b : _GEN_1085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1087 = 8'ha7 == r_count_4_io_out ? io_r_167_b : _GEN_1086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1088 = 8'ha8 == r_count_4_io_out ? io_r_168_b : _GEN_1087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1089 = 8'ha9 == r_count_4_io_out ? io_r_169_b : _GEN_1088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1090 = 8'haa == r_count_4_io_out ? io_r_170_b : _GEN_1089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1091 = 8'hab == r_count_4_io_out ? io_r_171_b : _GEN_1090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1092 = 8'hac == r_count_4_io_out ? io_r_172_b : _GEN_1091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1093 = 8'had == r_count_4_io_out ? io_r_173_b : _GEN_1092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1094 = 8'hae == r_count_4_io_out ? io_r_174_b : _GEN_1093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1095 = 8'haf == r_count_4_io_out ? io_r_175_b : _GEN_1094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1096 = 8'hb0 == r_count_4_io_out ? io_r_176_b : _GEN_1095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1097 = 8'hb1 == r_count_4_io_out ? io_r_177_b : _GEN_1096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1098 = 8'hb2 == r_count_4_io_out ? io_r_178_b : _GEN_1097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1099 = 8'hb3 == r_count_4_io_out ? io_r_179_b : _GEN_1098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1100 = 8'hb4 == r_count_4_io_out ? io_r_180_b : _GEN_1099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1101 = 8'hb5 == r_count_4_io_out ? io_r_181_b : _GEN_1100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1102 = 8'hb6 == r_count_4_io_out ? io_r_182_b : _GEN_1101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1103 = 8'hb7 == r_count_4_io_out ? io_r_183_b : _GEN_1102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1104 = 8'hb8 == r_count_4_io_out ? io_r_184_b : _GEN_1103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1105 = 8'hb9 == r_count_4_io_out ? io_r_185_b : _GEN_1104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1106 = 8'hba == r_count_4_io_out ? io_r_186_b : _GEN_1105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1107 = 8'hbb == r_count_4_io_out ? io_r_187_b : _GEN_1106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1108 = 8'hbc == r_count_4_io_out ? io_r_188_b : _GEN_1107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1109 = 8'hbd == r_count_4_io_out ? io_r_189_b : _GEN_1108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1110 = 8'hbe == r_count_4_io_out ? io_r_190_b : _GEN_1109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1111 = 8'hbf == r_count_4_io_out ? io_r_191_b : _GEN_1110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1112 = 8'hc0 == r_count_4_io_out ? io_r_192_b : _GEN_1111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1113 = 8'hc1 == r_count_4_io_out ? io_r_193_b : _GEN_1112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1114 = 8'hc2 == r_count_4_io_out ? io_r_194_b : _GEN_1113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1115 = 8'hc3 == r_count_4_io_out ? io_r_195_b : _GEN_1114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1116 = 8'hc4 == r_count_4_io_out ? io_r_196_b : _GEN_1115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1117 = 8'hc5 == r_count_4_io_out ? io_r_197_b : _GEN_1116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1118 = 8'hc6 == r_count_4_io_out ? io_r_198_b : _GEN_1117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1121 = 8'h1 == r_count_5_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1122 = 8'h2 == r_count_5_io_out ? io_r_2_b : _GEN_1121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1123 = 8'h3 == r_count_5_io_out ? io_r_3_b : _GEN_1122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1124 = 8'h4 == r_count_5_io_out ? io_r_4_b : _GEN_1123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1125 = 8'h5 == r_count_5_io_out ? io_r_5_b : _GEN_1124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1126 = 8'h6 == r_count_5_io_out ? io_r_6_b : _GEN_1125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1127 = 8'h7 == r_count_5_io_out ? io_r_7_b : _GEN_1126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1128 = 8'h8 == r_count_5_io_out ? io_r_8_b : _GEN_1127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1129 = 8'h9 == r_count_5_io_out ? io_r_9_b : _GEN_1128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1130 = 8'ha == r_count_5_io_out ? io_r_10_b : _GEN_1129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1131 = 8'hb == r_count_5_io_out ? io_r_11_b : _GEN_1130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1132 = 8'hc == r_count_5_io_out ? io_r_12_b : _GEN_1131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1133 = 8'hd == r_count_5_io_out ? io_r_13_b : _GEN_1132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1134 = 8'he == r_count_5_io_out ? io_r_14_b : _GEN_1133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1135 = 8'hf == r_count_5_io_out ? io_r_15_b : _GEN_1134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1136 = 8'h10 == r_count_5_io_out ? io_r_16_b : _GEN_1135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1137 = 8'h11 == r_count_5_io_out ? io_r_17_b : _GEN_1136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1138 = 8'h12 == r_count_5_io_out ? io_r_18_b : _GEN_1137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1139 = 8'h13 == r_count_5_io_out ? io_r_19_b : _GEN_1138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1140 = 8'h14 == r_count_5_io_out ? io_r_20_b : _GEN_1139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1141 = 8'h15 == r_count_5_io_out ? io_r_21_b : _GEN_1140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1142 = 8'h16 == r_count_5_io_out ? io_r_22_b : _GEN_1141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1143 = 8'h17 == r_count_5_io_out ? io_r_23_b : _GEN_1142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1144 = 8'h18 == r_count_5_io_out ? io_r_24_b : _GEN_1143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1145 = 8'h19 == r_count_5_io_out ? io_r_25_b : _GEN_1144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1146 = 8'h1a == r_count_5_io_out ? io_r_26_b : _GEN_1145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1147 = 8'h1b == r_count_5_io_out ? io_r_27_b : _GEN_1146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1148 = 8'h1c == r_count_5_io_out ? io_r_28_b : _GEN_1147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1149 = 8'h1d == r_count_5_io_out ? io_r_29_b : _GEN_1148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1150 = 8'h1e == r_count_5_io_out ? io_r_30_b : _GEN_1149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1151 = 8'h1f == r_count_5_io_out ? io_r_31_b : _GEN_1150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1152 = 8'h20 == r_count_5_io_out ? io_r_32_b : _GEN_1151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1153 = 8'h21 == r_count_5_io_out ? io_r_33_b : _GEN_1152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1154 = 8'h22 == r_count_5_io_out ? io_r_34_b : _GEN_1153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1155 = 8'h23 == r_count_5_io_out ? io_r_35_b : _GEN_1154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1156 = 8'h24 == r_count_5_io_out ? io_r_36_b : _GEN_1155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1157 = 8'h25 == r_count_5_io_out ? io_r_37_b : _GEN_1156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1158 = 8'h26 == r_count_5_io_out ? io_r_38_b : _GEN_1157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1159 = 8'h27 == r_count_5_io_out ? io_r_39_b : _GEN_1158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1160 = 8'h28 == r_count_5_io_out ? io_r_40_b : _GEN_1159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1161 = 8'h29 == r_count_5_io_out ? io_r_41_b : _GEN_1160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1162 = 8'h2a == r_count_5_io_out ? io_r_42_b : _GEN_1161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1163 = 8'h2b == r_count_5_io_out ? io_r_43_b : _GEN_1162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1164 = 8'h2c == r_count_5_io_out ? io_r_44_b : _GEN_1163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1165 = 8'h2d == r_count_5_io_out ? io_r_45_b : _GEN_1164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1166 = 8'h2e == r_count_5_io_out ? io_r_46_b : _GEN_1165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1167 = 8'h2f == r_count_5_io_out ? io_r_47_b : _GEN_1166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1168 = 8'h30 == r_count_5_io_out ? io_r_48_b : _GEN_1167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1169 = 8'h31 == r_count_5_io_out ? io_r_49_b : _GEN_1168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1170 = 8'h32 == r_count_5_io_out ? io_r_50_b : _GEN_1169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1171 = 8'h33 == r_count_5_io_out ? io_r_51_b : _GEN_1170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1172 = 8'h34 == r_count_5_io_out ? io_r_52_b : _GEN_1171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1173 = 8'h35 == r_count_5_io_out ? io_r_53_b : _GEN_1172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1174 = 8'h36 == r_count_5_io_out ? io_r_54_b : _GEN_1173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1175 = 8'h37 == r_count_5_io_out ? io_r_55_b : _GEN_1174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1176 = 8'h38 == r_count_5_io_out ? io_r_56_b : _GEN_1175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1177 = 8'h39 == r_count_5_io_out ? io_r_57_b : _GEN_1176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1178 = 8'h3a == r_count_5_io_out ? io_r_58_b : _GEN_1177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1179 = 8'h3b == r_count_5_io_out ? io_r_59_b : _GEN_1178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1180 = 8'h3c == r_count_5_io_out ? io_r_60_b : _GEN_1179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1181 = 8'h3d == r_count_5_io_out ? io_r_61_b : _GEN_1180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1182 = 8'h3e == r_count_5_io_out ? io_r_62_b : _GEN_1181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1183 = 8'h3f == r_count_5_io_out ? io_r_63_b : _GEN_1182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1184 = 8'h40 == r_count_5_io_out ? io_r_64_b : _GEN_1183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1185 = 8'h41 == r_count_5_io_out ? io_r_65_b : _GEN_1184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1186 = 8'h42 == r_count_5_io_out ? io_r_66_b : _GEN_1185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1187 = 8'h43 == r_count_5_io_out ? io_r_67_b : _GEN_1186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1188 = 8'h44 == r_count_5_io_out ? io_r_68_b : _GEN_1187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1189 = 8'h45 == r_count_5_io_out ? io_r_69_b : _GEN_1188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1190 = 8'h46 == r_count_5_io_out ? io_r_70_b : _GEN_1189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1191 = 8'h47 == r_count_5_io_out ? io_r_71_b : _GEN_1190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1192 = 8'h48 == r_count_5_io_out ? io_r_72_b : _GEN_1191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1193 = 8'h49 == r_count_5_io_out ? io_r_73_b : _GEN_1192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1194 = 8'h4a == r_count_5_io_out ? io_r_74_b : _GEN_1193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1195 = 8'h4b == r_count_5_io_out ? io_r_75_b : _GEN_1194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1196 = 8'h4c == r_count_5_io_out ? io_r_76_b : _GEN_1195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1197 = 8'h4d == r_count_5_io_out ? io_r_77_b : _GEN_1196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1198 = 8'h4e == r_count_5_io_out ? io_r_78_b : _GEN_1197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1199 = 8'h4f == r_count_5_io_out ? io_r_79_b : _GEN_1198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1200 = 8'h50 == r_count_5_io_out ? io_r_80_b : _GEN_1199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1201 = 8'h51 == r_count_5_io_out ? io_r_81_b : _GEN_1200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1202 = 8'h52 == r_count_5_io_out ? io_r_82_b : _GEN_1201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1203 = 8'h53 == r_count_5_io_out ? io_r_83_b : _GEN_1202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1204 = 8'h54 == r_count_5_io_out ? io_r_84_b : _GEN_1203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1205 = 8'h55 == r_count_5_io_out ? io_r_85_b : _GEN_1204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1206 = 8'h56 == r_count_5_io_out ? io_r_86_b : _GEN_1205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1207 = 8'h57 == r_count_5_io_out ? io_r_87_b : _GEN_1206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1208 = 8'h58 == r_count_5_io_out ? io_r_88_b : _GEN_1207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1209 = 8'h59 == r_count_5_io_out ? io_r_89_b : _GEN_1208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1210 = 8'h5a == r_count_5_io_out ? io_r_90_b : _GEN_1209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1211 = 8'h5b == r_count_5_io_out ? io_r_91_b : _GEN_1210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1212 = 8'h5c == r_count_5_io_out ? io_r_92_b : _GEN_1211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1213 = 8'h5d == r_count_5_io_out ? io_r_93_b : _GEN_1212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1214 = 8'h5e == r_count_5_io_out ? io_r_94_b : _GEN_1213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1215 = 8'h5f == r_count_5_io_out ? io_r_95_b : _GEN_1214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1216 = 8'h60 == r_count_5_io_out ? io_r_96_b : _GEN_1215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1217 = 8'h61 == r_count_5_io_out ? io_r_97_b : _GEN_1216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1218 = 8'h62 == r_count_5_io_out ? io_r_98_b : _GEN_1217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1219 = 8'h63 == r_count_5_io_out ? io_r_99_b : _GEN_1218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1220 = 8'h64 == r_count_5_io_out ? io_r_100_b : _GEN_1219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1221 = 8'h65 == r_count_5_io_out ? io_r_101_b : _GEN_1220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1222 = 8'h66 == r_count_5_io_out ? io_r_102_b : _GEN_1221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1223 = 8'h67 == r_count_5_io_out ? io_r_103_b : _GEN_1222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1224 = 8'h68 == r_count_5_io_out ? io_r_104_b : _GEN_1223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1225 = 8'h69 == r_count_5_io_out ? io_r_105_b : _GEN_1224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1226 = 8'h6a == r_count_5_io_out ? io_r_106_b : _GEN_1225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1227 = 8'h6b == r_count_5_io_out ? io_r_107_b : _GEN_1226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1228 = 8'h6c == r_count_5_io_out ? io_r_108_b : _GEN_1227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1229 = 8'h6d == r_count_5_io_out ? io_r_109_b : _GEN_1228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1230 = 8'h6e == r_count_5_io_out ? io_r_110_b : _GEN_1229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1231 = 8'h6f == r_count_5_io_out ? io_r_111_b : _GEN_1230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1232 = 8'h70 == r_count_5_io_out ? io_r_112_b : _GEN_1231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1233 = 8'h71 == r_count_5_io_out ? io_r_113_b : _GEN_1232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1234 = 8'h72 == r_count_5_io_out ? io_r_114_b : _GEN_1233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1235 = 8'h73 == r_count_5_io_out ? io_r_115_b : _GEN_1234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1236 = 8'h74 == r_count_5_io_out ? io_r_116_b : _GEN_1235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1237 = 8'h75 == r_count_5_io_out ? io_r_117_b : _GEN_1236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1238 = 8'h76 == r_count_5_io_out ? io_r_118_b : _GEN_1237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1239 = 8'h77 == r_count_5_io_out ? io_r_119_b : _GEN_1238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1240 = 8'h78 == r_count_5_io_out ? io_r_120_b : _GEN_1239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1241 = 8'h79 == r_count_5_io_out ? io_r_121_b : _GEN_1240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1242 = 8'h7a == r_count_5_io_out ? io_r_122_b : _GEN_1241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1243 = 8'h7b == r_count_5_io_out ? io_r_123_b : _GEN_1242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1244 = 8'h7c == r_count_5_io_out ? io_r_124_b : _GEN_1243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1245 = 8'h7d == r_count_5_io_out ? io_r_125_b : _GEN_1244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1246 = 8'h7e == r_count_5_io_out ? io_r_126_b : _GEN_1245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1247 = 8'h7f == r_count_5_io_out ? io_r_127_b : _GEN_1246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1248 = 8'h80 == r_count_5_io_out ? io_r_128_b : _GEN_1247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1249 = 8'h81 == r_count_5_io_out ? io_r_129_b : _GEN_1248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1250 = 8'h82 == r_count_5_io_out ? io_r_130_b : _GEN_1249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1251 = 8'h83 == r_count_5_io_out ? io_r_131_b : _GEN_1250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1252 = 8'h84 == r_count_5_io_out ? io_r_132_b : _GEN_1251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1253 = 8'h85 == r_count_5_io_out ? io_r_133_b : _GEN_1252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1254 = 8'h86 == r_count_5_io_out ? io_r_134_b : _GEN_1253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1255 = 8'h87 == r_count_5_io_out ? io_r_135_b : _GEN_1254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1256 = 8'h88 == r_count_5_io_out ? io_r_136_b : _GEN_1255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1257 = 8'h89 == r_count_5_io_out ? io_r_137_b : _GEN_1256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1258 = 8'h8a == r_count_5_io_out ? io_r_138_b : _GEN_1257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1259 = 8'h8b == r_count_5_io_out ? io_r_139_b : _GEN_1258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1260 = 8'h8c == r_count_5_io_out ? io_r_140_b : _GEN_1259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1261 = 8'h8d == r_count_5_io_out ? io_r_141_b : _GEN_1260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1262 = 8'h8e == r_count_5_io_out ? io_r_142_b : _GEN_1261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1263 = 8'h8f == r_count_5_io_out ? io_r_143_b : _GEN_1262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1264 = 8'h90 == r_count_5_io_out ? io_r_144_b : _GEN_1263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1265 = 8'h91 == r_count_5_io_out ? io_r_145_b : _GEN_1264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1266 = 8'h92 == r_count_5_io_out ? io_r_146_b : _GEN_1265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1267 = 8'h93 == r_count_5_io_out ? io_r_147_b : _GEN_1266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1268 = 8'h94 == r_count_5_io_out ? io_r_148_b : _GEN_1267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1269 = 8'h95 == r_count_5_io_out ? io_r_149_b : _GEN_1268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1270 = 8'h96 == r_count_5_io_out ? io_r_150_b : _GEN_1269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1271 = 8'h97 == r_count_5_io_out ? io_r_151_b : _GEN_1270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1272 = 8'h98 == r_count_5_io_out ? io_r_152_b : _GEN_1271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1273 = 8'h99 == r_count_5_io_out ? io_r_153_b : _GEN_1272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1274 = 8'h9a == r_count_5_io_out ? io_r_154_b : _GEN_1273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1275 = 8'h9b == r_count_5_io_out ? io_r_155_b : _GEN_1274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1276 = 8'h9c == r_count_5_io_out ? io_r_156_b : _GEN_1275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1277 = 8'h9d == r_count_5_io_out ? io_r_157_b : _GEN_1276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1278 = 8'h9e == r_count_5_io_out ? io_r_158_b : _GEN_1277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1279 = 8'h9f == r_count_5_io_out ? io_r_159_b : _GEN_1278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1280 = 8'ha0 == r_count_5_io_out ? io_r_160_b : _GEN_1279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1281 = 8'ha1 == r_count_5_io_out ? io_r_161_b : _GEN_1280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1282 = 8'ha2 == r_count_5_io_out ? io_r_162_b : _GEN_1281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1283 = 8'ha3 == r_count_5_io_out ? io_r_163_b : _GEN_1282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1284 = 8'ha4 == r_count_5_io_out ? io_r_164_b : _GEN_1283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1285 = 8'ha5 == r_count_5_io_out ? io_r_165_b : _GEN_1284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1286 = 8'ha6 == r_count_5_io_out ? io_r_166_b : _GEN_1285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1287 = 8'ha7 == r_count_5_io_out ? io_r_167_b : _GEN_1286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1288 = 8'ha8 == r_count_5_io_out ? io_r_168_b : _GEN_1287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1289 = 8'ha9 == r_count_5_io_out ? io_r_169_b : _GEN_1288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1290 = 8'haa == r_count_5_io_out ? io_r_170_b : _GEN_1289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1291 = 8'hab == r_count_5_io_out ? io_r_171_b : _GEN_1290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1292 = 8'hac == r_count_5_io_out ? io_r_172_b : _GEN_1291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1293 = 8'had == r_count_5_io_out ? io_r_173_b : _GEN_1292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1294 = 8'hae == r_count_5_io_out ? io_r_174_b : _GEN_1293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1295 = 8'haf == r_count_5_io_out ? io_r_175_b : _GEN_1294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1296 = 8'hb0 == r_count_5_io_out ? io_r_176_b : _GEN_1295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1297 = 8'hb1 == r_count_5_io_out ? io_r_177_b : _GEN_1296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1298 = 8'hb2 == r_count_5_io_out ? io_r_178_b : _GEN_1297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1299 = 8'hb3 == r_count_5_io_out ? io_r_179_b : _GEN_1298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1300 = 8'hb4 == r_count_5_io_out ? io_r_180_b : _GEN_1299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1301 = 8'hb5 == r_count_5_io_out ? io_r_181_b : _GEN_1300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1302 = 8'hb6 == r_count_5_io_out ? io_r_182_b : _GEN_1301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1303 = 8'hb7 == r_count_5_io_out ? io_r_183_b : _GEN_1302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1304 = 8'hb8 == r_count_5_io_out ? io_r_184_b : _GEN_1303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1305 = 8'hb9 == r_count_5_io_out ? io_r_185_b : _GEN_1304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1306 = 8'hba == r_count_5_io_out ? io_r_186_b : _GEN_1305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1307 = 8'hbb == r_count_5_io_out ? io_r_187_b : _GEN_1306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1308 = 8'hbc == r_count_5_io_out ? io_r_188_b : _GEN_1307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1309 = 8'hbd == r_count_5_io_out ? io_r_189_b : _GEN_1308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1310 = 8'hbe == r_count_5_io_out ? io_r_190_b : _GEN_1309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1311 = 8'hbf == r_count_5_io_out ? io_r_191_b : _GEN_1310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1312 = 8'hc0 == r_count_5_io_out ? io_r_192_b : _GEN_1311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1313 = 8'hc1 == r_count_5_io_out ? io_r_193_b : _GEN_1312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1314 = 8'hc2 == r_count_5_io_out ? io_r_194_b : _GEN_1313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1315 = 8'hc3 == r_count_5_io_out ? io_r_195_b : _GEN_1314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1316 = 8'hc4 == r_count_5_io_out ? io_r_196_b : _GEN_1315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1317 = 8'hc5 == r_count_5_io_out ? io_r_197_b : _GEN_1316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1318 = 8'hc6 == r_count_5_io_out ? io_r_198_b : _GEN_1317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1321 = 8'h1 == r_count_6_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1322 = 8'h2 == r_count_6_io_out ? io_r_2_b : _GEN_1321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1323 = 8'h3 == r_count_6_io_out ? io_r_3_b : _GEN_1322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1324 = 8'h4 == r_count_6_io_out ? io_r_4_b : _GEN_1323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1325 = 8'h5 == r_count_6_io_out ? io_r_5_b : _GEN_1324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1326 = 8'h6 == r_count_6_io_out ? io_r_6_b : _GEN_1325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1327 = 8'h7 == r_count_6_io_out ? io_r_7_b : _GEN_1326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1328 = 8'h8 == r_count_6_io_out ? io_r_8_b : _GEN_1327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1329 = 8'h9 == r_count_6_io_out ? io_r_9_b : _GEN_1328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1330 = 8'ha == r_count_6_io_out ? io_r_10_b : _GEN_1329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1331 = 8'hb == r_count_6_io_out ? io_r_11_b : _GEN_1330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1332 = 8'hc == r_count_6_io_out ? io_r_12_b : _GEN_1331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1333 = 8'hd == r_count_6_io_out ? io_r_13_b : _GEN_1332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1334 = 8'he == r_count_6_io_out ? io_r_14_b : _GEN_1333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1335 = 8'hf == r_count_6_io_out ? io_r_15_b : _GEN_1334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1336 = 8'h10 == r_count_6_io_out ? io_r_16_b : _GEN_1335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1337 = 8'h11 == r_count_6_io_out ? io_r_17_b : _GEN_1336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1338 = 8'h12 == r_count_6_io_out ? io_r_18_b : _GEN_1337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1339 = 8'h13 == r_count_6_io_out ? io_r_19_b : _GEN_1338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1340 = 8'h14 == r_count_6_io_out ? io_r_20_b : _GEN_1339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1341 = 8'h15 == r_count_6_io_out ? io_r_21_b : _GEN_1340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1342 = 8'h16 == r_count_6_io_out ? io_r_22_b : _GEN_1341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1343 = 8'h17 == r_count_6_io_out ? io_r_23_b : _GEN_1342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1344 = 8'h18 == r_count_6_io_out ? io_r_24_b : _GEN_1343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1345 = 8'h19 == r_count_6_io_out ? io_r_25_b : _GEN_1344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1346 = 8'h1a == r_count_6_io_out ? io_r_26_b : _GEN_1345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1347 = 8'h1b == r_count_6_io_out ? io_r_27_b : _GEN_1346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1348 = 8'h1c == r_count_6_io_out ? io_r_28_b : _GEN_1347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1349 = 8'h1d == r_count_6_io_out ? io_r_29_b : _GEN_1348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1350 = 8'h1e == r_count_6_io_out ? io_r_30_b : _GEN_1349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1351 = 8'h1f == r_count_6_io_out ? io_r_31_b : _GEN_1350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1352 = 8'h20 == r_count_6_io_out ? io_r_32_b : _GEN_1351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1353 = 8'h21 == r_count_6_io_out ? io_r_33_b : _GEN_1352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1354 = 8'h22 == r_count_6_io_out ? io_r_34_b : _GEN_1353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1355 = 8'h23 == r_count_6_io_out ? io_r_35_b : _GEN_1354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1356 = 8'h24 == r_count_6_io_out ? io_r_36_b : _GEN_1355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1357 = 8'h25 == r_count_6_io_out ? io_r_37_b : _GEN_1356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1358 = 8'h26 == r_count_6_io_out ? io_r_38_b : _GEN_1357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1359 = 8'h27 == r_count_6_io_out ? io_r_39_b : _GEN_1358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1360 = 8'h28 == r_count_6_io_out ? io_r_40_b : _GEN_1359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1361 = 8'h29 == r_count_6_io_out ? io_r_41_b : _GEN_1360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1362 = 8'h2a == r_count_6_io_out ? io_r_42_b : _GEN_1361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1363 = 8'h2b == r_count_6_io_out ? io_r_43_b : _GEN_1362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1364 = 8'h2c == r_count_6_io_out ? io_r_44_b : _GEN_1363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1365 = 8'h2d == r_count_6_io_out ? io_r_45_b : _GEN_1364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1366 = 8'h2e == r_count_6_io_out ? io_r_46_b : _GEN_1365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1367 = 8'h2f == r_count_6_io_out ? io_r_47_b : _GEN_1366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1368 = 8'h30 == r_count_6_io_out ? io_r_48_b : _GEN_1367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1369 = 8'h31 == r_count_6_io_out ? io_r_49_b : _GEN_1368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1370 = 8'h32 == r_count_6_io_out ? io_r_50_b : _GEN_1369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1371 = 8'h33 == r_count_6_io_out ? io_r_51_b : _GEN_1370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1372 = 8'h34 == r_count_6_io_out ? io_r_52_b : _GEN_1371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1373 = 8'h35 == r_count_6_io_out ? io_r_53_b : _GEN_1372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1374 = 8'h36 == r_count_6_io_out ? io_r_54_b : _GEN_1373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1375 = 8'h37 == r_count_6_io_out ? io_r_55_b : _GEN_1374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1376 = 8'h38 == r_count_6_io_out ? io_r_56_b : _GEN_1375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1377 = 8'h39 == r_count_6_io_out ? io_r_57_b : _GEN_1376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1378 = 8'h3a == r_count_6_io_out ? io_r_58_b : _GEN_1377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1379 = 8'h3b == r_count_6_io_out ? io_r_59_b : _GEN_1378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1380 = 8'h3c == r_count_6_io_out ? io_r_60_b : _GEN_1379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1381 = 8'h3d == r_count_6_io_out ? io_r_61_b : _GEN_1380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1382 = 8'h3e == r_count_6_io_out ? io_r_62_b : _GEN_1381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1383 = 8'h3f == r_count_6_io_out ? io_r_63_b : _GEN_1382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1384 = 8'h40 == r_count_6_io_out ? io_r_64_b : _GEN_1383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1385 = 8'h41 == r_count_6_io_out ? io_r_65_b : _GEN_1384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1386 = 8'h42 == r_count_6_io_out ? io_r_66_b : _GEN_1385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1387 = 8'h43 == r_count_6_io_out ? io_r_67_b : _GEN_1386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1388 = 8'h44 == r_count_6_io_out ? io_r_68_b : _GEN_1387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1389 = 8'h45 == r_count_6_io_out ? io_r_69_b : _GEN_1388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1390 = 8'h46 == r_count_6_io_out ? io_r_70_b : _GEN_1389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1391 = 8'h47 == r_count_6_io_out ? io_r_71_b : _GEN_1390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1392 = 8'h48 == r_count_6_io_out ? io_r_72_b : _GEN_1391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1393 = 8'h49 == r_count_6_io_out ? io_r_73_b : _GEN_1392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1394 = 8'h4a == r_count_6_io_out ? io_r_74_b : _GEN_1393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1395 = 8'h4b == r_count_6_io_out ? io_r_75_b : _GEN_1394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1396 = 8'h4c == r_count_6_io_out ? io_r_76_b : _GEN_1395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1397 = 8'h4d == r_count_6_io_out ? io_r_77_b : _GEN_1396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1398 = 8'h4e == r_count_6_io_out ? io_r_78_b : _GEN_1397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1399 = 8'h4f == r_count_6_io_out ? io_r_79_b : _GEN_1398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1400 = 8'h50 == r_count_6_io_out ? io_r_80_b : _GEN_1399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1401 = 8'h51 == r_count_6_io_out ? io_r_81_b : _GEN_1400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1402 = 8'h52 == r_count_6_io_out ? io_r_82_b : _GEN_1401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1403 = 8'h53 == r_count_6_io_out ? io_r_83_b : _GEN_1402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1404 = 8'h54 == r_count_6_io_out ? io_r_84_b : _GEN_1403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1405 = 8'h55 == r_count_6_io_out ? io_r_85_b : _GEN_1404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1406 = 8'h56 == r_count_6_io_out ? io_r_86_b : _GEN_1405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1407 = 8'h57 == r_count_6_io_out ? io_r_87_b : _GEN_1406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1408 = 8'h58 == r_count_6_io_out ? io_r_88_b : _GEN_1407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1409 = 8'h59 == r_count_6_io_out ? io_r_89_b : _GEN_1408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1410 = 8'h5a == r_count_6_io_out ? io_r_90_b : _GEN_1409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1411 = 8'h5b == r_count_6_io_out ? io_r_91_b : _GEN_1410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1412 = 8'h5c == r_count_6_io_out ? io_r_92_b : _GEN_1411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1413 = 8'h5d == r_count_6_io_out ? io_r_93_b : _GEN_1412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1414 = 8'h5e == r_count_6_io_out ? io_r_94_b : _GEN_1413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1415 = 8'h5f == r_count_6_io_out ? io_r_95_b : _GEN_1414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1416 = 8'h60 == r_count_6_io_out ? io_r_96_b : _GEN_1415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1417 = 8'h61 == r_count_6_io_out ? io_r_97_b : _GEN_1416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1418 = 8'h62 == r_count_6_io_out ? io_r_98_b : _GEN_1417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1419 = 8'h63 == r_count_6_io_out ? io_r_99_b : _GEN_1418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1420 = 8'h64 == r_count_6_io_out ? io_r_100_b : _GEN_1419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1421 = 8'h65 == r_count_6_io_out ? io_r_101_b : _GEN_1420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1422 = 8'h66 == r_count_6_io_out ? io_r_102_b : _GEN_1421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1423 = 8'h67 == r_count_6_io_out ? io_r_103_b : _GEN_1422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1424 = 8'h68 == r_count_6_io_out ? io_r_104_b : _GEN_1423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1425 = 8'h69 == r_count_6_io_out ? io_r_105_b : _GEN_1424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1426 = 8'h6a == r_count_6_io_out ? io_r_106_b : _GEN_1425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1427 = 8'h6b == r_count_6_io_out ? io_r_107_b : _GEN_1426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1428 = 8'h6c == r_count_6_io_out ? io_r_108_b : _GEN_1427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1429 = 8'h6d == r_count_6_io_out ? io_r_109_b : _GEN_1428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1430 = 8'h6e == r_count_6_io_out ? io_r_110_b : _GEN_1429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1431 = 8'h6f == r_count_6_io_out ? io_r_111_b : _GEN_1430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1432 = 8'h70 == r_count_6_io_out ? io_r_112_b : _GEN_1431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1433 = 8'h71 == r_count_6_io_out ? io_r_113_b : _GEN_1432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1434 = 8'h72 == r_count_6_io_out ? io_r_114_b : _GEN_1433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1435 = 8'h73 == r_count_6_io_out ? io_r_115_b : _GEN_1434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1436 = 8'h74 == r_count_6_io_out ? io_r_116_b : _GEN_1435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1437 = 8'h75 == r_count_6_io_out ? io_r_117_b : _GEN_1436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1438 = 8'h76 == r_count_6_io_out ? io_r_118_b : _GEN_1437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1439 = 8'h77 == r_count_6_io_out ? io_r_119_b : _GEN_1438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1440 = 8'h78 == r_count_6_io_out ? io_r_120_b : _GEN_1439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1441 = 8'h79 == r_count_6_io_out ? io_r_121_b : _GEN_1440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1442 = 8'h7a == r_count_6_io_out ? io_r_122_b : _GEN_1441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1443 = 8'h7b == r_count_6_io_out ? io_r_123_b : _GEN_1442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1444 = 8'h7c == r_count_6_io_out ? io_r_124_b : _GEN_1443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1445 = 8'h7d == r_count_6_io_out ? io_r_125_b : _GEN_1444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1446 = 8'h7e == r_count_6_io_out ? io_r_126_b : _GEN_1445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1447 = 8'h7f == r_count_6_io_out ? io_r_127_b : _GEN_1446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1448 = 8'h80 == r_count_6_io_out ? io_r_128_b : _GEN_1447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1449 = 8'h81 == r_count_6_io_out ? io_r_129_b : _GEN_1448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1450 = 8'h82 == r_count_6_io_out ? io_r_130_b : _GEN_1449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1451 = 8'h83 == r_count_6_io_out ? io_r_131_b : _GEN_1450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1452 = 8'h84 == r_count_6_io_out ? io_r_132_b : _GEN_1451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1453 = 8'h85 == r_count_6_io_out ? io_r_133_b : _GEN_1452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1454 = 8'h86 == r_count_6_io_out ? io_r_134_b : _GEN_1453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1455 = 8'h87 == r_count_6_io_out ? io_r_135_b : _GEN_1454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1456 = 8'h88 == r_count_6_io_out ? io_r_136_b : _GEN_1455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1457 = 8'h89 == r_count_6_io_out ? io_r_137_b : _GEN_1456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1458 = 8'h8a == r_count_6_io_out ? io_r_138_b : _GEN_1457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1459 = 8'h8b == r_count_6_io_out ? io_r_139_b : _GEN_1458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1460 = 8'h8c == r_count_6_io_out ? io_r_140_b : _GEN_1459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1461 = 8'h8d == r_count_6_io_out ? io_r_141_b : _GEN_1460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1462 = 8'h8e == r_count_6_io_out ? io_r_142_b : _GEN_1461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1463 = 8'h8f == r_count_6_io_out ? io_r_143_b : _GEN_1462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1464 = 8'h90 == r_count_6_io_out ? io_r_144_b : _GEN_1463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1465 = 8'h91 == r_count_6_io_out ? io_r_145_b : _GEN_1464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1466 = 8'h92 == r_count_6_io_out ? io_r_146_b : _GEN_1465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1467 = 8'h93 == r_count_6_io_out ? io_r_147_b : _GEN_1466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1468 = 8'h94 == r_count_6_io_out ? io_r_148_b : _GEN_1467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1469 = 8'h95 == r_count_6_io_out ? io_r_149_b : _GEN_1468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1470 = 8'h96 == r_count_6_io_out ? io_r_150_b : _GEN_1469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1471 = 8'h97 == r_count_6_io_out ? io_r_151_b : _GEN_1470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1472 = 8'h98 == r_count_6_io_out ? io_r_152_b : _GEN_1471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1473 = 8'h99 == r_count_6_io_out ? io_r_153_b : _GEN_1472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1474 = 8'h9a == r_count_6_io_out ? io_r_154_b : _GEN_1473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1475 = 8'h9b == r_count_6_io_out ? io_r_155_b : _GEN_1474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1476 = 8'h9c == r_count_6_io_out ? io_r_156_b : _GEN_1475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1477 = 8'h9d == r_count_6_io_out ? io_r_157_b : _GEN_1476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1478 = 8'h9e == r_count_6_io_out ? io_r_158_b : _GEN_1477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1479 = 8'h9f == r_count_6_io_out ? io_r_159_b : _GEN_1478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1480 = 8'ha0 == r_count_6_io_out ? io_r_160_b : _GEN_1479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1481 = 8'ha1 == r_count_6_io_out ? io_r_161_b : _GEN_1480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1482 = 8'ha2 == r_count_6_io_out ? io_r_162_b : _GEN_1481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1483 = 8'ha3 == r_count_6_io_out ? io_r_163_b : _GEN_1482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1484 = 8'ha4 == r_count_6_io_out ? io_r_164_b : _GEN_1483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1485 = 8'ha5 == r_count_6_io_out ? io_r_165_b : _GEN_1484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1486 = 8'ha6 == r_count_6_io_out ? io_r_166_b : _GEN_1485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1487 = 8'ha7 == r_count_6_io_out ? io_r_167_b : _GEN_1486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1488 = 8'ha8 == r_count_6_io_out ? io_r_168_b : _GEN_1487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1489 = 8'ha9 == r_count_6_io_out ? io_r_169_b : _GEN_1488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1490 = 8'haa == r_count_6_io_out ? io_r_170_b : _GEN_1489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1491 = 8'hab == r_count_6_io_out ? io_r_171_b : _GEN_1490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1492 = 8'hac == r_count_6_io_out ? io_r_172_b : _GEN_1491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1493 = 8'had == r_count_6_io_out ? io_r_173_b : _GEN_1492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1494 = 8'hae == r_count_6_io_out ? io_r_174_b : _GEN_1493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1495 = 8'haf == r_count_6_io_out ? io_r_175_b : _GEN_1494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1496 = 8'hb0 == r_count_6_io_out ? io_r_176_b : _GEN_1495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1497 = 8'hb1 == r_count_6_io_out ? io_r_177_b : _GEN_1496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1498 = 8'hb2 == r_count_6_io_out ? io_r_178_b : _GEN_1497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1499 = 8'hb3 == r_count_6_io_out ? io_r_179_b : _GEN_1498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1500 = 8'hb4 == r_count_6_io_out ? io_r_180_b : _GEN_1499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1501 = 8'hb5 == r_count_6_io_out ? io_r_181_b : _GEN_1500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1502 = 8'hb6 == r_count_6_io_out ? io_r_182_b : _GEN_1501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1503 = 8'hb7 == r_count_6_io_out ? io_r_183_b : _GEN_1502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1504 = 8'hb8 == r_count_6_io_out ? io_r_184_b : _GEN_1503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1505 = 8'hb9 == r_count_6_io_out ? io_r_185_b : _GEN_1504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1506 = 8'hba == r_count_6_io_out ? io_r_186_b : _GEN_1505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1507 = 8'hbb == r_count_6_io_out ? io_r_187_b : _GEN_1506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1508 = 8'hbc == r_count_6_io_out ? io_r_188_b : _GEN_1507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1509 = 8'hbd == r_count_6_io_out ? io_r_189_b : _GEN_1508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1510 = 8'hbe == r_count_6_io_out ? io_r_190_b : _GEN_1509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1511 = 8'hbf == r_count_6_io_out ? io_r_191_b : _GEN_1510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1512 = 8'hc0 == r_count_6_io_out ? io_r_192_b : _GEN_1511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1513 = 8'hc1 == r_count_6_io_out ? io_r_193_b : _GEN_1512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1514 = 8'hc2 == r_count_6_io_out ? io_r_194_b : _GEN_1513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1515 = 8'hc3 == r_count_6_io_out ? io_r_195_b : _GEN_1514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1516 = 8'hc4 == r_count_6_io_out ? io_r_196_b : _GEN_1515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1517 = 8'hc5 == r_count_6_io_out ? io_r_197_b : _GEN_1516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1518 = 8'hc6 == r_count_6_io_out ? io_r_198_b : _GEN_1517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1521 = 8'h1 == r_count_7_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1522 = 8'h2 == r_count_7_io_out ? io_r_2_b : _GEN_1521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1523 = 8'h3 == r_count_7_io_out ? io_r_3_b : _GEN_1522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1524 = 8'h4 == r_count_7_io_out ? io_r_4_b : _GEN_1523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1525 = 8'h5 == r_count_7_io_out ? io_r_5_b : _GEN_1524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1526 = 8'h6 == r_count_7_io_out ? io_r_6_b : _GEN_1525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1527 = 8'h7 == r_count_7_io_out ? io_r_7_b : _GEN_1526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1528 = 8'h8 == r_count_7_io_out ? io_r_8_b : _GEN_1527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1529 = 8'h9 == r_count_7_io_out ? io_r_9_b : _GEN_1528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1530 = 8'ha == r_count_7_io_out ? io_r_10_b : _GEN_1529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1531 = 8'hb == r_count_7_io_out ? io_r_11_b : _GEN_1530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1532 = 8'hc == r_count_7_io_out ? io_r_12_b : _GEN_1531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1533 = 8'hd == r_count_7_io_out ? io_r_13_b : _GEN_1532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1534 = 8'he == r_count_7_io_out ? io_r_14_b : _GEN_1533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1535 = 8'hf == r_count_7_io_out ? io_r_15_b : _GEN_1534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1536 = 8'h10 == r_count_7_io_out ? io_r_16_b : _GEN_1535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1537 = 8'h11 == r_count_7_io_out ? io_r_17_b : _GEN_1536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1538 = 8'h12 == r_count_7_io_out ? io_r_18_b : _GEN_1537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1539 = 8'h13 == r_count_7_io_out ? io_r_19_b : _GEN_1538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1540 = 8'h14 == r_count_7_io_out ? io_r_20_b : _GEN_1539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1541 = 8'h15 == r_count_7_io_out ? io_r_21_b : _GEN_1540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1542 = 8'h16 == r_count_7_io_out ? io_r_22_b : _GEN_1541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1543 = 8'h17 == r_count_7_io_out ? io_r_23_b : _GEN_1542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1544 = 8'h18 == r_count_7_io_out ? io_r_24_b : _GEN_1543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1545 = 8'h19 == r_count_7_io_out ? io_r_25_b : _GEN_1544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1546 = 8'h1a == r_count_7_io_out ? io_r_26_b : _GEN_1545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1547 = 8'h1b == r_count_7_io_out ? io_r_27_b : _GEN_1546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1548 = 8'h1c == r_count_7_io_out ? io_r_28_b : _GEN_1547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1549 = 8'h1d == r_count_7_io_out ? io_r_29_b : _GEN_1548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1550 = 8'h1e == r_count_7_io_out ? io_r_30_b : _GEN_1549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1551 = 8'h1f == r_count_7_io_out ? io_r_31_b : _GEN_1550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1552 = 8'h20 == r_count_7_io_out ? io_r_32_b : _GEN_1551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1553 = 8'h21 == r_count_7_io_out ? io_r_33_b : _GEN_1552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1554 = 8'h22 == r_count_7_io_out ? io_r_34_b : _GEN_1553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1555 = 8'h23 == r_count_7_io_out ? io_r_35_b : _GEN_1554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1556 = 8'h24 == r_count_7_io_out ? io_r_36_b : _GEN_1555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1557 = 8'h25 == r_count_7_io_out ? io_r_37_b : _GEN_1556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1558 = 8'h26 == r_count_7_io_out ? io_r_38_b : _GEN_1557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1559 = 8'h27 == r_count_7_io_out ? io_r_39_b : _GEN_1558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1560 = 8'h28 == r_count_7_io_out ? io_r_40_b : _GEN_1559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1561 = 8'h29 == r_count_7_io_out ? io_r_41_b : _GEN_1560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1562 = 8'h2a == r_count_7_io_out ? io_r_42_b : _GEN_1561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1563 = 8'h2b == r_count_7_io_out ? io_r_43_b : _GEN_1562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1564 = 8'h2c == r_count_7_io_out ? io_r_44_b : _GEN_1563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1565 = 8'h2d == r_count_7_io_out ? io_r_45_b : _GEN_1564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1566 = 8'h2e == r_count_7_io_out ? io_r_46_b : _GEN_1565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1567 = 8'h2f == r_count_7_io_out ? io_r_47_b : _GEN_1566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1568 = 8'h30 == r_count_7_io_out ? io_r_48_b : _GEN_1567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1569 = 8'h31 == r_count_7_io_out ? io_r_49_b : _GEN_1568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1570 = 8'h32 == r_count_7_io_out ? io_r_50_b : _GEN_1569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1571 = 8'h33 == r_count_7_io_out ? io_r_51_b : _GEN_1570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1572 = 8'h34 == r_count_7_io_out ? io_r_52_b : _GEN_1571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1573 = 8'h35 == r_count_7_io_out ? io_r_53_b : _GEN_1572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1574 = 8'h36 == r_count_7_io_out ? io_r_54_b : _GEN_1573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1575 = 8'h37 == r_count_7_io_out ? io_r_55_b : _GEN_1574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1576 = 8'h38 == r_count_7_io_out ? io_r_56_b : _GEN_1575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1577 = 8'h39 == r_count_7_io_out ? io_r_57_b : _GEN_1576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1578 = 8'h3a == r_count_7_io_out ? io_r_58_b : _GEN_1577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1579 = 8'h3b == r_count_7_io_out ? io_r_59_b : _GEN_1578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1580 = 8'h3c == r_count_7_io_out ? io_r_60_b : _GEN_1579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1581 = 8'h3d == r_count_7_io_out ? io_r_61_b : _GEN_1580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1582 = 8'h3e == r_count_7_io_out ? io_r_62_b : _GEN_1581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1583 = 8'h3f == r_count_7_io_out ? io_r_63_b : _GEN_1582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1584 = 8'h40 == r_count_7_io_out ? io_r_64_b : _GEN_1583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1585 = 8'h41 == r_count_7_io_out ? io_r_65_b : _GEN_1584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1586 = 8'h42 == r_count_7_io_out ? io_r_66_b : _GEN_1585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1587 = 8'h43 == r_count_7_io_out ? io_r_67_b : _GEN_1586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1588 = 8'h44 == r_count_7_io_out ? io_r_68_b : _GEN_1587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1589 = 8'h45 == r_count_7_io_out ? io_r_69_b : _GEN_1588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1590 = 8'h46 == r_count_7_io_out ? io_r_70_b : _GEN_1589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1591 = 8'h47 == r_count_7_io_out ? io_r_71_b : _GEN_1590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1592 = 8'h48 == r_count_7_io_out ? io_r_72_b : _GEN_1591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1593 = 8'h49 == r_count_7_io_out ? io_r_73_b : _GEN_1592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1594 = 8'h4a == r_count_7_io_out ? io_r_74_b : _GEN_1593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1595 = 8'h4b == r_count_7_io_out ? io_r_75_b : _GEN_1594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1596 = 8'h4c == r_count_7_io_out ? io_r_76_b : _GEN_1595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1597 = 8'h4d == r_count_7_io_out ? io_r_77_b : _GEN_1596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1598 = 8'h4e == r_count_7_io_out ? io_r_78_b : _GEN_1597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1599 = 8'h4f == r_count_7_io_out ? io_r_79_b : _GEN_1598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1600 = 8'h50 == r_count_7_io_out ? io_r_80_b : _GEN_1599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1601 = 8'h51 == r_count_7_io_out ? io_r_81_b : _GEN_1600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1602 = 8'h52 == r_count_7_io_out ? io_r_82_b : _GEN_1601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1603 = 8'h53 == r_count_7_io_out ? io_r_83_b : _GEN_1602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1604 = 8'h54 == r_count_7_io_out ? io_r_84_b : _GEN_1603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1605 = 8'h55 == r_count_7_io_out ? io_r_85_b : _GEN_1604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1606 = 8'h56 == r_count_7_io_out ? io_r_86_b : _GEN_1605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1607 = 8'h57 == r_count_7_io_out ? io_r_87_b : _GEN_1606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1608 = 8'h58 == r_count_7_io_out ? io_r_88_b : _GEN_1607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1609 = 8'h59 == r_count_7_io_out ? io_r_89_b : _GEN_1608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1610 = 8'h5a == r_count_7_io_out ? io_r_90_b : _GEN_1609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1611 = 8'h5b == r_count_7_io_out ? io_r_91_b : _GEN_1610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1612 = 8'h5c == r_count_7_io_out ? io_r_92_b : _GEN_1611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1613 = 8'h5d == r_count_7_io_out ? io_r_93_b : _GEN_1612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1614 = 8'h5e == r_count_7_io_out ? io_r_94_b : _GEN_1613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1615 = 8'h5f == r_count_7_io_out ? io_r_95_b : _GEN_1614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1616 = 8'h60 == r_count_7_io_out ? io_r_96_b : _GEN_1615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1617 = 8'h61 == r_count_7_io_out ? io_r_97_b : _GEN_1616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1618 = 8'h62 == r_count_7_io_out ? io_r_98_b : _GEN_1617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1619 = 8'h63 == r_count_7_io_out ? io_r_99_b : _GEN_1618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1620 = 8'h64 == r_count_7_io_out ? io_r_100_b : _GEN_1619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1621 = 8'h65 == r_count_7_io_out ? io_r_101_b : _GEN_1620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1622 = 8'h66 == r_count_7_io_out ? io_r_102_b : _GEN_1621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1623 = 8'h67 == r_count_7_io_out ? io_r_103_b : _GEN_1622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1624 = 8'h68 == r_count_7_io_out ? io_r_104_b : _GEN_1623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1625 = 8'h69 == r_count_7_io_out ? io_r_105_b : _GEN_1624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1626 = 8'h6a == r_count_7_io_out ? io_r_106_b : _GEN_1625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1627 = 8'h6b == r_count_7_io_out ? io_r_107_b : _GEN_1626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1628 = 8'h6c == r_count_7_io_out ? io_r_108_b : _GEN_1627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1629 = 8'h6d == r_count_7_io_out ? io_r_109_b : _GEN_1628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1630 = 8'h6e == r_count_7_io_out ? io_r_110_b : _GEN_1629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1631 = 8'h6f == r_count_7_io_out ? io_r_111_b : _GEN_1630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1632 = 8'h70 == r_count_7_io_out ? io_r_112_b : _GEN_1631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1633 = 8'h71 == r_count_7_io_out ? io_r_113_b : _GEN_1632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1634 = 8'h72 == r_count_7_io_out ? io_r_114_b : _GEN_1633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1635 = 8'h73 == r_count_7_io_out ? io_r_115_b : _GEN_1634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1636 = 8'h74 == r_count_7_io_out ? io_r_116_b : _GEN_1635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1637 = 8'h75 == r_count_7_io_out ? io_r_117_b : _GEN_1636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1638 = 8'h76 == r_count_7_io_out ? io_r_118_b : _GEN_1637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1639 = 8'h77 == r_count_7_io_out ? io_r_119_b : _GEN_1638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1640 = 8'h78 == r_count_7_io_out ? io_r_120_b : _GEN_1639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1641 = 8'h79 == r_count_7_io_out ? io_r_121_b : _GEN_1640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1642 = 8'h7a == r_count_7_io_out ? io_r_122_b : _GEN_1641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1643 = 8'h7b == r_count_7_io_out ? io_r_123_b : _GEN_1642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1644 = 8'h7c == r_count_7_io_out ? io_r_124_b : _GEN_1643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1645 = 8'h7d == r_count_7_io_out ? io_r_125_b : _GEN_1644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1646 = 8'h7e == r_count_7_io_out ? io_r_126_b : _GEN_1645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1647 = 8'h7f == r_count_7_io_out ? io_r_127_b : _GEN_1646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1648 = 8'h80 == r_count_7_io_out ? io_r_128_b : _GEN_1647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1649 = 8'h81 == r_count_7_io_out ? io_r_129_b : _GEN_1648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1650 = 8'h82 == r_count_7_io_out ? io_r_130_b : _GEN_1649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1651 = 8'h83 == r_count_7_io_out ? io_r_131_b : _GEN_1650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1652 = 8'h84 == r_count_7_io_out ? io_r_132_b : _GEN_1651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1653 = 8'h85 == r_count_7_io_out ? io_r_133_b : _GEN_1652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1654 = 8'h86 == r_count_7_io_out ? io_r_134_b : _GEN_1653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1655 = 8'h87 == r_count_7_io_out ? io_r_135_b : _GEN_1654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1656 = 8'h88 == r_count_7_io_out ? io_r_136_b : _GEN_1655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1657 = 8'h89 == r_count_7_io_out ? io_r_137_b : _GEN_1656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1658 = 8'h8a == r_count_7_io_out ? io_r_138_b : _GEN_1657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1659 = 8'h8b == r_count_7_io_out ? io_r_139_b : _GEN_1658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1660 = 8'h8c == r_count_7_io_out ? io_r_140_b : _GEN_1659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1661 = 8'h8d == r_count_7_io_out ? io_r_141_b : _GEN_1660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1662 = 8'h8e == r_count_7_io_out ? io_r_142_b : _GEN_1661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1663 = 8'h8f == r_count_7_io_out ? io_r_143_b : _GEN_1662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1664 = 8'h90 == r_count_7_io_out ? io_r_144_b : _GEN_1663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1665 = 8'h91 == r_count_7_io_out ? io_r_145_b : _GEN_1664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1666 = 8'h92 == r_count_7_io_out ? io_r_146_b : _GEN_1665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1667 = 8'h93 == r_count_7_io_out ? io_r_147_b : _GEN_1666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1668 = 8'h94 == r_count_7_io_out ? io_r_148_b : _GEN_1667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1669 = 8'h95 == r_count_7_io_out ? io_r_149_b : _GEN_1668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1670 = 8'h96 == r_count_7_io_out ? io_r_150_b : _GEN_1669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1671 = 8'h97 == r_count_7_io_out ? io_r_151_b : _GEN_1670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1672 = 8'h98 == r_count_7_io_out ? io_r_152_b : _GEN_1671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1673 = 8'h99 == r_count_7_io_out ? io_r_153_b : _GEN_1672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1674 = 8'h9a == r_count_7_io_out ? io_r_154_b : _GEN_1673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1675 = 8'h9b == r_count_7_io_out ? io_r_155_b : _GEN_1674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1676 = 8'h9c == r_count_7_io_out ? io_r_156_b : _GEN_1675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1677 = 8'h9d == r_count_7_io_out ? io_r_157_b : _GEN_1676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1678 = 8'h9e == r_count_7_io_out ? io_r_158_b : _GEN_1677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1679 = 8'h9f == r_count_7_io_out ? io_r_159_b : _GEN_1678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1680 = 8'ha0 == r_count_7_io_out ? io_r_160_b : _GEN_1679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1681 = 8'ha1 == r_count_7_io_out ? io_r_161_b : _GEN_1680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1682 = 8'ha2 == r_count_7_io_out ? io_r_162_b : _GEN_1681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1683 = 8'ha3 == r_count_7_io_out ? io_r_163_b : _GEN_1682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1684 = 8'ha4 == r_count_7_io_out ? io_r_164_b : _GEN_1683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1685 = 8'ha5 == r_count_7_io_out ? io_r_165_b : _GEN_1684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1686 = 8'ha6 == r_count_7_io_out ? io_r_166_b : _GEN_1685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1687 = 8'ha7 == r_count_7_io_out ? io_r_167_b : _GEN_1686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1688 = 8'ha8 == r_count_7_io_out ? io_r_168_b : _GEN_1687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1689 = 8'ha9 == r_count_7_io_out ? io_r_169_b : _GEN_1688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1690 = 8'haa == r_count_7_io_out ? io_r_170_b : _GEN_1689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1691 = 8'hab == r_count_7_io_out ? io_r_171_b : _GEN_1690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1692 = 8'hac == r_count_7_io_out ? io_r_172_b : _GEN_1691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1693 = 8'had == r_count_7_io_out ? io_r_173_b : _GEN_1692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1694 = 8'hae == r_count_7_io_out ? io_r_174_b : _GEN_1693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1695 = 8'haf == r_count_7_io_out ? io_r_175_b : _GEN_1694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1696 = 8'hb0 == r_count_7_io_out ? io_r_176_b : _GEN_1695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1697 = 8'hb1 == r_count_7_io_out ? io_r_177_b : _GEN_1696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1698 = 8'hb2 == r_count_7_io_out ? io_r_178_b : _GEN_1697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1699 = 8'hb3 == r_count_7_io_out ? io_r_179_b : _GEN_1698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1700 = 8'hb4 == r_count_7_io_out ? io_r_180_b : _GEN_1699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1701 = 8'hb5 == r_count_7_io_out ? io_r_181_b : _GEN_1700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1702 = 8'hb6 == r_count_7_io_out ? io_r_182_b : _GEN_1701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1703 = 8'hb7 == r_count_7_io_out ? io_r_183_b : _GEN_1702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1704 = 8'hb8 == r_count_7_io_out ? io_r_184_b : _GEN_1703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1705 = 8'hb9 == r_count_7_io_out ? io_r_185_b : _GEN_1704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1706 = 8'hba == r_count_7_io_out ? io_r_186_b : _GEN_1705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1707 = 8'hbb == r_count_7_io_out ? io_r_187_b : _GEN_1706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1708 = 8'hbc == r_count_7_io_out ? io_r_188_b : _GEN_1707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1709 = 8'hbd == r_count_7_io_out ? io_r_189_b : _GEN_1708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1710 = 8'hbe == r_count_7_io_out ? io_r_190_b : _GEN_1709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1711 = 8'hbf == r_count_7_io_out ? io_r_191_b : _GEN_1710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1712 = 8'hc0 == r_count_7_io_out ? io_r_192_b : _GEN_1711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1713 = 8'hc1 == r_count_7_io_out ? io_r_193_b : _GEN_1712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1714 = 8'hc2 == r_count_7_io_out ? io_r_194_b : _GEN_1713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1715 = 8'hc3 == r_count_7_io_out ? io_r_195_b : _GEN_1714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1716 = 8'hc4 == r_count_7_io_out ? io_r_196_b : _GEN_1715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1717 = 8'hc5 == r_count_7_io_out ? io_r_197_b : _GEN_1716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1718 = 8'hc6 == r_count_7_io_out ? io_r_198_b : _GEN_1717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1721 = 8'h1 == r_count_8_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1722 = 8'h2 == r_count_8_io_out ? io_r_2_b : _GEN_1721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1723 = 8'h3 == r_count_8_io_out ? io_r_3_b : _GEN_1722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1724 = 8'h4 == r_count_8_io_out ? io_r_4_b : _GEN_1723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1725 = 8'h5 == r_count_8_io_out ? io_r_5_b : _GEN_1724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1726 = 8'h6 == r_count_8_io_out ? io_r_6_b : _GEN_1725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1727 = 8'h7 == r_count_8_io_out ? io_r_7_b : _GEN_1726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1728 = 8'h8 == r_count_8_io_out ? io_r_8_b : _GEN_1727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1729 = 8'h9 == r_count_8_io_out ? io_r_9_b : _GEN_1728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1730 = 8'ha == r_count_8_io_out ? io_r_10_b : _GEN_1729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1731 = 8'hb == r_count_8_io_out ? io_r_11_b : _GEN_1730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1732 = 8'hc == r_count_8_io_out ? io_r_12_b : _GEN_1731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1733 = 8'hd == r_count_8_io_out ? io_r_13_b : _GEN_1732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1734 = 8'he == r_count_8_io_out ? io_r_14_b : _GEN_1733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1735 = 8'hf == r_count_8_io_out ? io_r_15_b : _GEN_1734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1736 = 8'h10 == r_count_8_io_out ? io_r_16_b : _GEN_1735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1737 = 8'h11 == r_count_8_io_out ? io_r_17_b : _GEN_1736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1738 = 8'h12 == r_count_8_io_out ? io_r_18_b : _GEN_1737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1739 = 8'h13 == r_count_8_io_out ? io_r_19_b : _GEN_1738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1740 = 8'h14 == r_count_8_io_out ? io_r_20_b : _GEN_1739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1741 = 8'h15 == r_count_8_io_out ? io_r_21_b : _GEN_1740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1742 = 8'h16 == r_count_8_io_out ? io_r_22_b : _GEN_1741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1743 = 8'h17 == r_count_8_io_out ? io_r_23_b : _GEN_1742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1744 = 8'h18 == r_count_8_io_out ? io_r_24_b : _GEN_1743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1745 = 8'h19 == r_count_8_io_out ? io_r_25_b : _GEN_1744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1746 = 8'h1a == r_count_8_io_out ? io_r_26_b : _GEN_1745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1747 = 8'h1b == r_count_8_io_out ? io_r_27_b : _GEN_1746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1748 = 8'h1c == r_count_8_io_out ? io_r_28_b : _GEN_1747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1749 = 8'h1d == r_count_8_io_out ? io_r_29_b : _GEN_1748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1750 = 8'h1e == r_count_8_io_out ? io_r_30_b : _GEN_1749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1751 = 8'h1f == r_count_8_io_out ? io_r_31_b : _GEN_1750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1752 = 8'h20 == r_count_8_io_out ? io_r_32_b : _GEN_1751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1753 = 8'h21 == r_count_8_io_out ? io_r_33_b : _GEN_1752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1754 = 8'h22 == r_count_8_io_out ? io_r_34_b : _GEN_1753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1755 = 8'h23 == r_count_8_io_out ? io_r_35_b : _GEN_1754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1756 = 8'h24 == r_count_8_io_out ? io_r_36_b : _GEN_1755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1757 = 8'h25 == r_count_8_io_out ? io_r_37_b : _GEN_1756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1758 = 8'h26 == r_count_8_io_out ? io_r_38_b : _GEN_1757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1759 = 8'h27 == r_count_8_io_out ? io_r_39_b : _GEN_1758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1760 = 8'h28 == r_count_8_io_out ? io_r_40_b : _GEN_1759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1761 = 8'h29 == r_count_8_io_out ? io_r_41_b : _GEN_1760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1762 = 8'h2a == r_count_8_io_out ? io_r_42_b : _GEN_1761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1763 = 8'h2b == r_count_8_io_out ? io_r_43_b : _GEN_1762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1764 = 8'h2c == r_count_8_io_out ? io_r_44_b : _GEN_1763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1765 = 8'h2d == r_count_8_io_out ? io_r_45_b : _GEN_1764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1766 = 8'h2e == r_count_8_io_out ? io_r_46_b : _GEN_1765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1767 = 8'h2f == r_count_8_io_out ? io_r_47_b : _GEN_1766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1768 = 8'h30 == r_count_8_io_out ? io_r_48_b : _GEN_1767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1769 = 8'h31 == r_count_8_io_out ? io_r_49_b : _GEN_1768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1770 = 8'h32 == r_count_8_io_out ? io_r_50_b : _GEN_1769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1771 = 8'h33 == r_count_8_io_out ? io_r_51_b : _GEN_1770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1772 = 8'h34 == r_count_8_io_out ? io_r_52_b : _GEN_1771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1773 = 8'h35 == r_count_8_io_out ? io_r_53_b : _GEN_1772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1774 = 8'h36 == r_count_8_io_out ? io_r_54_b : _GEN_1773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1775 = 8'h37 == r_count_8_io_out ? io_r_55_b : _GEN_1774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1776 = 8'h38 == r_count_8_io_out ? io_r_56_b : _GEN_1775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1777 = 8'h39 == r_count_8_io_out ? io_r_57_b : _GEN_1776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1778 = 8'h3a == r_count_8_io_out ? io_r_58_b : _GEN_1777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1779 = 8'h3b == r_count_8_io_out ? io_r_59_b : _GEN_1778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1780 = 8'h3c == r_count_8_io_out ? io_r_60_b : _GEN_1779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1781 = 8'h3d == r_count_8_io_out ? io_r_61_b : _GEN_1780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1782 = 8'h3e == r_count_8_io_out ? io_r_62_b : _GEN_1781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1783 = 8'h3f == r_count_8_io_out ? io_r_63_b : _GEN_1782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1784 = 8'h40 == r_count_8_io_out ? io_r_64_b : _GEN_1783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1785 = 8'h41 == r_count_8_io_out ? io_r_65_b : _GEN_1784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1786 = 8'h42 == r_count_8_io_out ? io_r_66_b : _GEN_1785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1787 = 8'h43 == r_count_8_io_out ? io_r_67_b : _GEN_1786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1788 = 8'h44 == r_count_8_io_out ? io_r_68_b : _GEN_1787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1789 = 8'h45 == r_count_8_io_out ? io_r_69_b : _GEN_1788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1790 = 8'h46 == r_count_8_io_out ? io_r_70_b : _GEN_1789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1791 = 8'h47 == r_count_8_io_out ? io_r_71_b : _GEN_1790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1792 = 8'h48 == r_count_8_io_out ? io_r_72_b : _GEN_1791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1793 = 8'h49 == r_count_8_io_out ? io_r_73_b : _GEN_1792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1794 = 8'h4a == r_count_8_io_out ? io_r_74_b : _GEN_1793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1795 = 8'h4b == r_count_8_io_out ? io_r_75_b : _GEN_1794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1796 = 8'h4c == r_count_8_io_out ? io_r_76_b : _GEN_1795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1797 = 8'h4d == r_count_8_io_out ? io_r_77_b : _GEN_1796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1798 = 8'h4e == r_count_8_io_out ? io_r_78_b : _GEN_1797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1799 = 8'h4f == r_count_8_io_out ? io_r_79_b : _GEN_1798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1800 = 8'h50 == r_count_8_io_out ? io_r_80_b : _GEN_1799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1801 = 8'h51 == r_count_8_io_out ? io_r_81_b : _GEN_1800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1802 = 8'h52 == r_count_8_io_out ? io_r_82_b : _GEN_1801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1803 = 8'h53 == r_count_8_io_out ? io_r_83_b : _GEN_1802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1804 = 8'h54 == r_count_8_io_out ? io_r_84_b : _GEN_1803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1805 = 8'h55 == r_count_8_io_out ? io_r_85_b : _GEN_1804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1806 = 8'h56 == r_count_8_io_out ? io_r_86_b : _GEN_1805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1807 = 8'h57 == r_count_8_io_out ? io_r_87_b : _GEN_1806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1808 = 8'h58 == r_count_8_io_out ? io_r_88_b : _GEN_1807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1809 = 8'h59 == r_count_8_io_out ? io_r_89_b : _GEN_1808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1810 = 8'h5a == r_count_8_io_out ? io_r_90_b : _GEN_1809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1811 = 8'h5b == r_count_8_io_out ? io_r_91_b : _GEN_1810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1812 = 8'h5c == r_count_8_io_out ? io_r_92_b : _GEN_1811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1813 = 8'h5d == r_count_8_io_out ? io_r_93_b : _GEN_1812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1814 = 8'h5e == r_count_8_io_out ? io_r_94_b : _GEN_1813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1815 = 8'h5f == r_count_8_io_out ? io_r_95_b : _GEN_1814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1816 = 8'h60 == r_count_8_io_out ? io_r_96_b : _GEN_1815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1817 = 8'h61 == r_count_8_io_out ? io_r_97_b : _GEN_1816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1818 = 8'h62 == r_count_8_io_out ? io_r_98_b : _GEN_1817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1819 = 8'h63 == r_count_8_io_out ? io_r_99_b : _GEN_1818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1820 = 8'h64 == r_count_8_io_out ? io_r_100_b : _GEN_1819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1821 = 8'h65 == r_count_8_io_out ? io_r_101_b : _GEN_1820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1822 = 8'h66 == r_count_8_io_out ? io_r_102_b : _GEN_1821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1823 = 8'h67 == r_count_8_io_out ? io_r_103_b : _GEN_1822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1824 = 8'h68 == r_count_8_io_out ? io_r_104_b : _GEN_1823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1825 = 8'h69 == r_count_8_io_out ? io_r_105_b : _GEN_1824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1826 = 8'h6a == r_count_8_io_out ? io_r_106_b : _GEN_1825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1827 = 8'h6b == r_count_8_io_out ? io_r_107_b : _GEN_1826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1828 = 8'h6c == r_count_8_io_out ? io_r_108_b : _GEN_1827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1829 = 8'h6d == r_count_8_io_out ? io_r_109_b : _GEN_1828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1830 = 8'h6e == r_count_8_io_out ? io_r_110_b : _GEN_1829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1831 = 8'h6f == r_count_8_io_out ? io_r_111_b : _GEN_1830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1832 = 8'h70 == r_count_8_io_out ? io_r_112_b : _GEN_1831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1833 = 8'h71 == r_count_8_io_out ? io_r_113_b : _GEN_1832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1834 = 8'h72 == r_count_8_io_out ? io_r_114_b : _GEN_1833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1835 = 8'h73 == r_count_8_io_out ? io_r_115_b : _GEN_1834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1836 = 8'h74 == r_count_8_io_out ? io_r_116_b : _GEN_1835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1837 = 8'h75 == r_count_8_io_out ? io_r_117_b : _GEN_1836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1838 = 8'h76 == r_count_8_io_out ? io_r_118_b : _GEN_1837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1839 = 8'h77 == r_count_8_io_out ? io_r_119_b : _GEN_1838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1840 = 8'h78 == r_count_8_io_out ? io_r_120_b : _GEN_1839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1841 = 8'h79 == r_count_8_io_out ? io_r_121_b : _GEN_1840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1842 = 8'h7a == r_count_8_io_out ? io_r_122_b : _GEN_1841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1843 = 8'h7b == r_count_8_io_out ? io_r_123_b : _GEN_1842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1844 = 8'h7c == r_count_8_io_out ? io_r_124_b : _GEN_1843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1845 = 8'h7d == r_count_8_io_out ? io_r_125_b : _GEN_1844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1846 = 8'h7e == r_count_8_io_out ? io_r_126_b : _GEN_1845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1847 = 8'h7f == r_count_8_io_out ? io_r_127_b : _GEN_1846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1848 = 8'h80 == r_count_8_io_out ? io_r_128_b : _GEN_1847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1849 = 8'h81 == r_count_8_io_out ? io_r_129_b : _GEN_1848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1850 = 8'h82 == r_count_8_io_out ? io_r_130_b : _GEN_1849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1851 = 8'h83 == r_count_8_io_out ? io_r_131_b : _GEN_1850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1852 = 8'h84 == r_count_8_io_out ? io_r_132_b : _GEN_1851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1853 = 8'h85 == r_count_8_io_out ? io_r_133_b : _GEN_1852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1854 = 8'h86 == r_count_8_io_out ? io_r_134_b : _GEN_1853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1855 = 8'h87 == r_count_8_io_out ? io_r_135_b : _GEN_1854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1856 = 8'h88 == r_count_8_io_out ? io_r_136_b : _GEN_1855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1857 = 8'h89 == r_count_8_io_out ? io_r_137_b : _GEN_1856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1858 = 8'h8a == r_count_8_io_out ? io_r_138_b : _GEN_1857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1859 = 8'h8b == r_count_8_io_out ? io_r_139_b : _GEN_1858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1860 = 8'h8c == r_count_8_io_out ? io_r_140_b : _GEN_1859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1861 = 8'h8d == r_count_8_io_out ? io_r_141_b : _GEN_1860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1862 = 8'h8e == r_count_8_io_out ? io_r_142_b : _GEN_1861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1863 = 8'h8f == r_count_8_io_out ? io_r_143_b : _GEN_1862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1864 = 8'h90 == r_count_8_io_out ? io_r_144_b : _GEN_1863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1865 = 8'h91 == r_count_8_io_out ? io_r_145_b : _GEN_1864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1866 = 8'h92 == r_count_8_io_out ? io_r_146_b : _GEN_1865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1867 = 8'h93 == r_count_8_io_out ? io_r_147_b : _GEN_1866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1868 = 8'h94 == r_count_8_io_out ? io_r_148_b : _GEN_1867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1869 = 8'h95 == r_count_8_io_out ? io_r_149_b : _GEN_1868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1870 = 8'h96 == r_count_8_io_out ? io_r_150_b : _GEN_1869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1871 = 8'h97 == r_count_8_io_out ? io_r_151_b : _GEN_1870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1872 = 8'h98 == r_count_8_io_out ? io_r_152_b : _GEN_1871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1873 = 8'h99 == r_count_8_io_out ? io_r_153_b : _GEN_1872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1874 = 8'h9a == r_count_8_io_out ? io_r_154_b : _GEN_1873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1875 = 8'h9b == r_count_8_io_out ? io_r_155_b : _GEN_1874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1876 = 8'h9c == r_count_8_io_out ? io_r_156_b : _GEN_1875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1877 = 8'h9d == r_count_8_io_out ? io_r_157_b : _GEN_1876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1878 = 8'h9e == r_count_8_io_out ? io_r_158_b : _GEN_1877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1879 = 8'h9f == r_count_8_io_out ? io_r_159_b : _GEN_1878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1880 = 8'ha0 == r_count_8_io_out ? io_r_160_b : _GEN_1879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1881 = 8'ha1 == r_count_8_io_out ? io_r_161_b : _GEN_1880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1882 = 8'ha2 == r_count_8_io_out ? io_r_162_b : _GEN_1881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1883 = 8'ha3 == r_count_8_io_out ? io_r_163_b : _GEN_1882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1884 = 8'ha4 == r_count_8_io_out ? io_r_164_b : _GEN_1883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1885 = 8'ha5 == r_count_8_io_out ? io_r_165_b : _GEN_1884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1886 = 8'ha6 == r_count_8_io_out ? io_r_166_b : _GEN_1885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1887 = 8'ha7 == r_count_8_io_out ? io_r_167_b : _GEN_1886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1888 = 8'ha8 == r_count_8_io_out ? io_r_168_b : _GEN_1887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1889 = 8'ha9 == r_count_8_io_out ? io_r_169_b : _GEN_1888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1890 = 8'haa == r_count_8_io_out ? io_r_170_b : _GEN_1889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1891 = 8'hab == r_count_8_io_out ? io_r_171_b : _GEN_1890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1892 = 8'hac == r_count_8_io_out ? io_r_172_b : _GEN_1891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1893 = 8'had == r_count_8_io_out ? io_r_173_b : _GEN_1892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1894 = 8'hae == r_count_8_io_out ? io_r_174_b : _GEN_1893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1895 = 8'haf == r_count_8_io_out ? io_r_175_b : _GEN_1894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1896 = 8'hb0 == r_count_8_io_out ? io_r_176_b : _GEN_1895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1897 = 8'hb1 == r_count_8_io_out ? io_r_177_b : _GEN_1896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1898 = 8'hb2 == r_count_8_io_out ? io_r_178_b : _GEN_1897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1899 = 8'hb3 == r_count_8_io_out ? io_r_179_b : _GEN_1898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1900 = 8'hb4 == r_count_8_io_out ? io_r_180_b : _GEN_1899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1901 = 8'hb5 == r_count_8_io_out ? io_r_181_b : _GEN_1900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1902 = 8'hb6 == r_count_8_io_out ? io_r_182_b : _GEN_1901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1903 = 8'hb7 == r_count_8_io_out ? io_r_183_b : _GEN_1902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1904 = 8'hb8 == r_count_8_io_out ? io_r_184_b : _GEN_1903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1905 = 8'hb9 == r_count_8_io_out ? io_r_185_b : _GEN_1904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1906 = 8'hba == r_count_8_io_out ? io_r_186_b : _GEN_1905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1907 = 8'hbb == r_count_8_io_out ? io_r_187_b : _GEN_1906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1908 = 8'hbc == r_count_8_io_out ? io_r_188_b : _GEN_1907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1909 = 8'hbd == r_count_8_io_out ? io_r_189_b : _GEN_1908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1910 = 8'hbe == r_count_8_io_out ? io_r_190_b : _GEN_1909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1911 = 8'hbf == r_count_8_io_out ? io_r_191_b : _GEN_1910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1912 = 8'hc0 == r_count_8_io_out ? io_r_192_b : _GEN_1911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1913 = 8'hc1 == r_count_8_io_out ? io_r_193_b : _GEN_1912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1914 = 8'hc2 == r_count_8_io_out ? io_r_194_b : _GEN_1913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1915 = 8'hc3 == r_count_8_io_out ? io_r_195_b : _GEN_1914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1916 = 8'hc4 == r_count_8_io_out ? io_r_196_b : _GEN_1915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1917 = 8'hc5 == r_count_8_io_out ? io_r_197_b : _GEN_1916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1918 = 8'hc6 == r_count_8_io_out ? io_r_198_b : _GEN_1917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1921 = 8'h1 == r_count_9_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1922 = 8'h2 == r_count_9_io_out ? io_r_2_b : _GEN_1921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1923 = 8'h3 == r_count_9_io_out ? io_r_3_b : _GEN_1922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1924 = 8'h4 == r_count_9_io_out ? io_r_4_b : _GEN_1923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1925 = 8'h5 == r_count_9_io_out ? io_r_5_b : _GEN_1924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1926 = 8'h6 == r_count_9_io_out ? io_r_6_b : _GEN_1925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1927 = 8'h7 == r_count_9_io_out ? io_r_7_b : _GEN_1926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1928 = 8'h8 == r_count_9_io_out ? io_r_8_b : _GEN_1927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1929 = 8'h9 == r_count_9_io_out ? io_r_9_b : _GEN_1928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1930 = 8'ha == r_count_9_io_out ? io_r_10_b : _GEN_1929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1931 = 8'hb == r_count_9_io_out ? io_r_11_b : _GEN_1930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1932 = 8'hc == r_count_9_io_out ? io_r_12_b : _GEN_1931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1933 = 8'hd == r_count_9_io_out ? io_r_13_b : _GEN_1932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1934 = 8'he == r_count_9_io_out ? io_r_14_b : _GEN_1933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1935 = 8'hf == r_count_9_io_out ? io_r_15_b : _GEN_1934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1936 = 8'h10 == r_count_9_io_out ? io_r_16_b : _GEN_1935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1937 = 8'h11 == r_count_9_io_out ? io_r_17_b : _GEN_1936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1938 = 8'h12 == r_count_9_io_out ? io_r_18_b : _GEN_1937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1939 = 8'h13 == r_count_9_io_out ? io_r_19_b : _GEN_1938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1940 = 8'h14 == r_count_9_io_out ? io_r_20_b : _GEN_1939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1941 = 8'h15 == r_count_9_io_out ? io_r_21_b : _GEN_1940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1942 = 8'h16 == r_count_9_io_out ? io_r_22_b : _GEN_1941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1943 = 8'h17 == r_count_9_io_out ? io_r_23_b : _GEN_1942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1944 = 8'h18 == r_count_9_io_out ? io_r_24_b : _GEN_1943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1945 = 8'h19 == r_count_9_io_out ? io_r_25_b : _GEN_1944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1946 = 8'h1a == r_count_9_io_out ? io_r_26_b : _GEN_1945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1947 = 8'h1b == r_count_9_io_out ? io_r_27_b : _GEN_1946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1948 = 8'h1c == r_count_9_io_out ? io_r_28_b : _GEN_1947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1949 = 8'h1d == r_count_9_io_out ? io_r_29_b : _GEN_1948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1950 = 8'h1e == r_count_9_io_out ? io_r_30_b : _GEN_1949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1951 = 8'h1f == r_count_9_io_out ? io_r_31_b : _GEN_1950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1952 = 8'h20 == r_count_9_io_out ? io_r_32_b : _GEN_1951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1953 = 8'h21 == r_count_9_io_out ? io_r_33_b : _GEN_1952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1954 = 8'h22 == r_count_9_io_out ? io_r_34_b : _GEN_1953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1955 = 8'h23 == r_count_9_io_out ? io_r_35_b : _GEN_1954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1956 = 8'h24 == r_count_9_io_out ? io_r_36_b : _GEN_1955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1957 = 8'h25 == r_count_9_io_out ? io_r_37_b : _GEN_1956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1958 = 8'h26 == r_count_9_io_out ? io_r_38_b : _GEN_1957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1959 = 8'h27 == r_count_9_io_out ? io_r_39_b : _GEN_1958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1960 = 8'h28 == r_count_9_io_out ? io_r_40_b : _GEN_1959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1961 = 8'h29 == r_count_9_io_out ? io_r_41_b : _GEN_1960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1962 = 8'h2a == r_count_9_io_out ? io_r_42_b : _GEN_1961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1963 = 8'h2b == r_count_9_io_out ? io_r_43_b : _GEN_1962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1964 = 8'h2c == r_count_9_io_out ? io_r_44_b : _GEN_1963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1965 = 8'h2d == r_count_9_io_out ? io_r_45_b : _GEN_1964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1966 = 8'h2e == r_count_9_io_out ? io_r_46_b : _GEN_1965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1967 = 8'h2f == r_count_9_io_out ? io_r_47_b : _GEN_1966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1968 = 8'h30 == r_count_9_io_out ? io_r_48_b : _GEN_1967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1969 = 8'h31 == r_count_9_io_out ? io_r_49_b : _GEN_1968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1970 = 8'h32 == r_count_9_io_out ? io_r_50_b : _GEN_1969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1971 = 8'h33 == r_count_9_io_out ? io_r_51_b : _GEN_1970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1972 = 8'h34 == r_count_9_io_out ? io_r_52_b : _GEN_1971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1973 = 8'h35 == r_count_9_io_out ? io_r_53_b : _GEN_1972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1974 = 8'h36 == r_count_9_io_out ? io_r_54_b : _GEN_1973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1975 = 8'h37 == r_count_9_io_out ? io_r_55_b : _GEN_1974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1976 = 8'h38 == r_count_9_io_out ? io_r_56_b : _GEN_1975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1977 = 8'h39 == r_count_9_io_out ? io_r_57_b : _GEN_1976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1978 = 8'h3a == r_count_9_io_out ? io_r_58_b : _GEN_1977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1979 = 8'h3b == r_count_9_io_out ? io_r_59_b : _GEN_1978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1980 = 8'h3c == r_count_9_io_out ? io_r_60_b : _GEN_1979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1981 = 8'h3d == r_count_9_io_out ? io_r_61_b : _GEN_1980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1982 = 8'h3e == r_count_9_io_out ? io_r_62_b : _GEN_1981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1983 = 8'h3f == r_count_9_io_out ? io_r_63_b : _GEN_1982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1984 = 8'h40 == r_count_9_io_out ? io_r_64_b : _GEN_1983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1985 = 8'h41 == r_count_9_io_out ? io_r_65_b : _GEN_1984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1986 = 8'h42 == r_count_9_io_out ? io_r_66_b : _GEN_1985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1987 = 8'h43 == r_count_9_io_out ? io_r_67_b : _GEN_1986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1988 = 8'h44 == r_count_9_io_out ? io_r_68_b : _GEN_1987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1989 = 8'h45 == r_count_9_io_out ? io_r_69_b : _GEN_1988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1990 = 8'h46 == r_count_9_io_out ? io_r_70_b : _GEN_1989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1991 = 8'h47 == r_count_9_io_out ? io_r_71_b : _GEN_1990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1992 = 8'h48 == r_count_9_io_out ? io_r_72_b : _GEN_1991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1993 = 8'h49 == r_count_9_io_out ? io_r_73_b : _GEN_1992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1994 = 8'h4a == r_count_9_io_out ? io_r_74_b : _GEN_1993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1995 = 8'h4b == r_count_9_io_out ? io_r_75_b : _GEN_1994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1996 = 8'h4c == r_count_9_io_out ? io_r_76_b : _GEN_1995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1997 = 8'h4d == r_count_9_io_out ? io_r_77_b : _GEN_1996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1998 = 8'h4e == r_count_9_io_out ? io_r_78_b : _GEN_1997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1999 = 8'h4f == r_count_9_io_out ? io_r_79_b : _GEN_1998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2000 = 8'h50 == r_count_9_io_out ? io_r_80_b : _GEN_1999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2001 = 8'h51 == r_count_9_io_out ? io_r_81_b : _GEN_2000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2002 = 8'h52 == r_count_9_io_out ? io_r_82_b : _GEN_2001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2003 = 8'h53 == r_count_9_io_out ? io_r_83_b : _GEN_2002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2004 = 8'h54 == r_count_9_io_out ? io_r_84_b : _GEN_2003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2005 = 8'h55 == r_count_9_io_out ? io_r_85_b : _GEN_2004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2006 = 8'h56 == r_count_9_io_out ? io_r_86_b : _GEN_2005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2007 = 8'h57 == r_count_9_io_out ? io_r_87_b : _GEN_2006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2008 = 8'h58 == r_count_9_io_out ? io_r_88_b : _GEN_2007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2009 = 8'h59 == r_count_9_io_out ? io_r_89_b : _GEN_2008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2010 = 8'h5a == r_count_9_io_out ? io_r_90_b : _GEN_2009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2011 = 8'h5b == r_count_9_io_out ? io_r_91_b : _GEN_2010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2012 = 8'h5c == r_count_9_io_out ? io_r_92_b : _GEN_2011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2013 = 8'h5d == r_count_9_io_out ? io_r_93_b : _GEN_2012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2014 = 8'h5e == r_count_9_io_out ? io_r_94_b : _GEN_2013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2015 = 8'h5f == r_count_9_io_out ? io_r_95_b : _GEN_2014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2016 = 8'h60 == r_count_9_io_out ? io_r_96_b : _GEN_2015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2017 = 8'h61 == r_count_9_io_out ? io_r_97_b : _GEN_2016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2018 = 8'h62 == r_count_9_io_out ? io_r_98_b : _GEN_2017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2019 = 8'h63 == r_count_9_io_out ? io_r_99_b : _GEN_2018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2020 = 8'h64 == r_count_9_io_out ? io_r_100_b : _GEN_2019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2021 = 8'h65 == r_count_9_io_out ? io_r_101_b : _GEN_2020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2022 = 8'h66 == r_count_9_io_out ? io_r_102_b : _GEN_2021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2023 = 8'h67 == r_count_9_io_out ? io_r_103_b : _GEN_2022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2024 = 8'h68 == r_count_9_io_out ? io_r_104_b : _GEN_2023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2025 = 8'h69 == r_count_9_io_out ? io_r_105_b : _GEN_2024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2026 = 8'h6a == r_count_9_io_out ? io_r_106_b : _GEN_2025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2027 = 8'h6b == r_count_9_io_out ? io_r_107_b : _GEN_2026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2028 = 8'h6c == r_count_9_io_out ? io_r_108_b : _GEN_2027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2029 = 8'h6d == r_count_9_io_out ? io_r_109_b : _GEN_2028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2030 = 8'h6e == r_count_9_io_out ? io_r_110_b : _GEN_2029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2031 = 8'h6f == r_count_9_io_out ? io_r_111_b : _GEN_2030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2032 = 8'h70 == r_count_9_io_out ? io_r_112_b : _GEN_2031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2033 = 8'h71 == r_count_9_io_out ? io_r_113_b : _GEN_2032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2034 = 8'h72 == r_count_9_io_out ? io_r_114_b : _GEN_2033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2035 = 8'h73 == r_count_9_io_out ? io_r_115_b : _GEN_2034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2036 = 8'h74 == r_count_9_io_out ? io_r_116_b : _GEN_2035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2037 = 8'h75 == r_count_9_io_out ? io_r_117_b : _GEN_2036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2038 = 8'h76 == r_count_9_io_out ? io_r_118_b : _GEN_2037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2039 = 8'h77 == r_count_9_io_out ? io_r_119_b : _GEN_2038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2040 = 8'h78 == r_count_9_io_out ? io_r_120_b : _GEN_2039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2041 = 8'h79 == r_count_9_io_out ? io_r_121_b : _GEN_2040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2042 = 8'h7a == r_count_9_io_out ? io_r_122_b : _GEN_2041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2043 = 8'h7b == r_count_9_io_out ? io_r_123_b : _GEN_2042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2044 = 8'h7c == r_count_9_io_out ? io_r_124_b : _GEN_2043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2045 = 8'h7d == r_count_9_io_out ? io_r_125_b : _GEN_2044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2046 = 8'h7e == r_count_9_io_out ? io_r_126_b : _GEN_2045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2047 = 8'h7f == r_count_9_io_out ? io_r_127_b : _GEN_2046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2048 = 8'h80 == r_count_9_io_out ? io_r_128_b : _GEN_2047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2049 = 8'h81 == r_count_9_io_out ? io_r_129_b : _GEN_2048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2050 = 8'h82 == r_count_9_io_out ? io_r_130_b : _GEN_2049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2051 = 8'h83 == r_count_9_io_out ? io_r_131_b : _GEN_2050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2052 = 8'h84 == r_count_9_io_out ? io_r_132_b : _GEN_2051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2053 = 8'h85 == r_count_9_io_out ? io_r_133_b : _GEN_2052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2054 = 8'h86 == r_count_9_io_out ? io_r_134_b : _GEN_2053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2055 = 8'h87 == r_count_9_io_out ? io_r_135_b : _GEN_2054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2056 = 8'h88 == r_count_9_io_out ? io_r_136_b : _GEN_2055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2057 = 8'h89 == r_count_9_io_out ? io_r_137_b : _GEN_2056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2058 = 8'h8a == r_count_9_io_out ? io_r_138_b : _GEN_2057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2059 = 8'h8b == r_count_9_io_out ? io_r_139_b : _GEN_2058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2060 = 8'h8c == r_count_9_io_out ? io_r_140_b : _GEN_2059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2061 = 8'h8d == r_count_9_io_out ? io_r_141_b : _GEN_2060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2062 = 8'h8e == r_count_9_io_out ? io_r_142_b : _GEN_2061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2063 = 8'h8f == r_count_9_io_out ? io_r_143_b : _GEN_2062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2064 = 8'h90 == r_count_9_io_out ? io_r_144_b : _GEN_2063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2065 = 8'h91 == r_count_9_io_out ? io_r_145_b : _GEN_2064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2066 = 8'h92 == r_count_9_io_out ? io_r_146_b : _GEN_2065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2067 = 8'h93 == r_count_9_io_out ? io_r_147_b : _GEN_2066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2068 = 8'h94 == r_count_9_io_out ? io_r_148_b : _GEN_2067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2069 = 8'h95 == r_count_9_io_out ? io_r_149_b : _GEN_2068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2070 = 8'h96 == r_count_9_io_out ? io_r_150_b : _GEN_2069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2071 = 8'h97 == r_count_9_io_out ? io_r_151_b : _GEN_2070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2072 = 8'h98 == r_count_9_io_out ? io_r_152_b : _GEN_2071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2073 = 8'h99 == r_count_9_io_out ? io_r_153_b : _GEN_2072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2074 = 8'h9a == r_count_9_io_out ? io_r_154_b : _GEN_2073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2075 = 8'h9b == r_count_9_io_out ? io_r_155_b : _GEN_2074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2076 = 8'h9c == r_count_9_io_out ? io_r_156_b : _GEN_2075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2077 = 8'h9d == r_count_9_io_out ? io_r_157_b : _GEN_2076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2078 = 8'h9e == r_count_9_io_out ? io_r_158_b : _GEN_2077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2079 = 8'h9f == r_count_9_io_out ? io_r_159_b : _GEN_2078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2080 = 8'ha0 == r_count_9_io_out ? io_r_160_b : _GEN_2079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2081 = 8'ha1 == r_count_9_io_out ? io_r_161_b : _GEN_2080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2082 = 8'ha2 == r_count_9_io_out ? io_r_162_b : _GEN_2081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2083 = 8'ha3 == r_count_9_io_out ? io_r_163_b : _GEN_2082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2084 = 8'ha4 == r_count_9_io_out ? io_r_164_b : _GEN_2083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2085 = 8'ha5 == r_count_9_io_out ? io_r_165_b : _GEN_2084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2086 = 8'ha6 == r_count_9_io_out ? io_r_166_b : _GEN_2085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2087 = 8'ha7 == r_count_9_io_out ? io_r_167_b : _GEN_2086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2088 = 8'ha8 == r_count_9_io_out ? io_r_168_b : _GEN_2087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2089 = 8'ha9 == r_count_9_io_out ? io_r_169_b : _GEN_2088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2090 = 8'haa == r_count_9_io_out ? io_r_170_b : _GEN_2089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2091 = 8'hab == r_count_9_io_out ? io_r_171_b : _GEN_2090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2092 = 8'hac == r_count_9_io_out ? io_r_172_b : _GEN_2091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2093 = 8'had == r_count_9_io_out ? io_r_173_b : _GEN_2092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2094 = 8'hae == r_count_9_io_out ? io_r_174_b : _GEN_2093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2095 = 8'haf == r_count_9_io_out ? io_r_175_b : _GEN_2094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2096 = 8'hb0 == r_count_9_io_out ? io_r_176_b : _GEN_2095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2097 = 8'hb1 == r_count_9_io_out ? io_r_177_b : _GEN_2096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2098 = 8'hb2 == r_count_9_io_out ? io_r_178_b : _GEN_2097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2099 = 8'hb3 == r_count_9_io_out ? io_r_179_b : _GEN_2098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2100 = 8'hb4 == r_count_9_io_out ? io_r_180_b : _GEN_2099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2101 = 8'hb5 == r_count_9_io_out ? io_r_181_b : _GEN_2100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2102 = 8'hb6 == r_count_9_io_out ? io_r_182_b : _GEN_2101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2103 = 8'hb7 == r_count_9_io_out ? io_r_183_b : _GEN_2102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2104 = 8'hb8 == r_count_9_io_out ? io_r_184_b : _GEN_2103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2105 = 8'hb9 == r_count_9_io_out ? io_r_185_b : _GEN_2104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2106 = 8'hba == r_count_9_io_out ? io_r_186_b : _GEN_2105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2107 = 8'hbb == r_count_9_io_out ? io_r_187_b : _GEN_2106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2108 = 8'hbc == r_count_9_io_out ? io_r_188_b : _GEN_2107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2109 = 8'hbd == r_count_9_io_out ? io_r_189_b : _GEN_2108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2110 = 8'hbe == r_count_9_io_out ? io_r_190_b : _GEN_2109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2111 = 8'hbf == r_count_9_io_out ? io_r_191_b : _GEN_2110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2112 = 8'hc0 == r_count_9_io_out ? io_r_192_b : _GEN_2111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2113 = 8'hc1 == r_count_9_io_out ? io_r_193_b : _GEN_2112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2114 = 8'hc2 == r_count_9_io_out ? io_r_194_b : _GEN_2113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2115 = 8'hc3 == r_count_9_io_out ? io_r_195_b : _GEN_2114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2116 = 8'hc4 == r_count_9_io_out ? io_r_196_b : _GEN_2115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2117 = 8'hc5 == r_count_9_io_out ? io_r_197_b : _GEN_2116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2118 = 8'hc6 == r_count_9_io_out ? io_r_198_b : _GEN_2117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2121 = 8'h1 == r_count_10_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2122 = 8'h2 == r_count_10_io_out ? io_r_2_b : _GEN_2121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2123 = 8'h3 == r_count_10_io_out ? io_r_3_b : _GEN_2122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2124 = 8'h4 == r_count_10_io_out ? io_r_4_b : _GEN_2123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2125 = 8'h5 == r_count_10_io_out ? io_r_5_b : _GEN_2124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2126 = 8'h6 == r_count_10_io_out ? io_r_6_b : _GEN_2125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2127 = 8'h7 == r_count_10_io_out ? io_r_7_b : _GEN_2126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2128 = 8'h8 == r_count_10_io_out ? io_r_8_b : _GEN_2127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2129 = 8'h9 == r_count_10_io_out ? io_r_9_b : _GEN_2128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2130 = 8'ha == r_count_10_io_out ? io_r_10_b : _GEN_2129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2131 = 8'hb == r_count_10_io_out ? io_r_11_b : _GEN_2130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2132 = 8'hc == r_count_10_io_out ? io_r_12_b : _GEN_2131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2133 = 8'hd == r_count_10_io_out ? io_r_13_b : _GEN_2132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2134 = 8'he == r_count_10_io_out ? io_r_14_b : _GEN_2133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2135 = 8'hf == r_count_10_io_out ? io_r_15_b : _GEN_2134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2136 = 8'h10 == r_count_10_io_out ? io_r_16_b : _GEN_2135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2137 = 8'h11 == r_count_10_io_out ? io_r_17_b : _GEN_2136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2138 = 8'h12 == r_count_10_io_out ? io_r_18_b : _GEN_2137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2139 = 8'h13 == r_count_10_io_out ? io_r_19_b : _GEN_2138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2140 = 8'h14 == r_count_10_io_out ? io_r_20_b : _GEN_2139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2141 = 8'h15 == r_count_10_io_out ? io_r_21_b : _GEN_2140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2142 = 8'h16 == r_count_10_io_out ? io_r_22_b : _GEN_2141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2143 = 8'h17 == r_count_10_io_out ? io_r_23_b : _GEN_2142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2144 = 8'h18 == r_count_10_io_out ? io_r_24_b : _GEN_2143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2145 = 8'h19 == r_count_10_io_out ? io_r_25_b : _GEN_2144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2146 = 8'h1a == r_count_10_io_out ? io_r_26_b : _GEN_2145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2147 = 8'h1b == r_count_10_io_out ? io_r_27_b : _GEN_2146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2148 = 8'h1c == r_count_10_io_out ? io_r_28_b : _GEN_2147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2149 = 8'h1d == r_count_10_io_out ? io_r_29_b : _GEN_2148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2150 = 8'h1e == r_count_10_io_out ? io_r_30_b : _GEN_2149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2151 = 8'h1f == r_count_10_io_out ? io_r_31_b : _GEN_2150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2152 = 8'h20 == r_count_10_io_out ? io_r_32_b : _GEN_2151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2153 = 8'h21 == r_count_10_io_out ? io_r_33_b : _GEN_2152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2154 = 8'h22 == r_count_10_io_out ? io_r_34_b : _GEN_2153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2155 = 8'h23 == r_count_10_io_out ? io_r_35_b : _GEN_2154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2156 = 8'h24 == r_count_10_io_out ? io_r_36_b : _GEN_2155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2157 = 8'h25 == r_count_10_io_out ? io_r_37_b : _GEN_2156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2158 = 8'h26 == r_count_10_io_out ? io_r_38_b : _GEN_2157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2159 = 8'h27 == r_count_10_io_out ? io_r_39_b : _GEN_2158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2160 = 8'h28 == r_count_10_io_out ? io_r_40_b : _GEN_2159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2161 = 8'h29 == r_count_10_io_out ? io_r_41_b : _GEN_2160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2162 = 8'h2a == r_count_10_io_out ? io_r_42_b : _GEN_2161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2163 = 8'h2b == r_count_10_io_out ? io_r_43_b : _GEN_2162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2164 = 8'h2c == r_count_10_io_out ? io_r_44_b : _GEN_2163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2165 = 8'h2d == r_count_10_io_out ? io_r_45_b : _GEN_2164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2166 = 8'h2e == r_count_10_io_out ? io_r_46_b : _GEN_2165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2167 = 8'h2f == r_count_10_io_out ? io_r_47_b : _GEN_2166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2168 = 8'h30 == r_count_10_io_out ? io_r_48_b : _GEN_2167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2169 = 8'h31 == r_count_10_io_out ? io_r_49_b : _GEN_2168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2170 = 8'h32 == r_count_10_io_out ? io_r_50_b : _GEN_2169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2171 = 8'h33 == r_count_10_io_out ? io_r_51_b : _GEN_2170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2172 = 8'h34 == r_count_10_io_out ? io_r_52_b : _GEN_2171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2173 = 8'h35 == r_count_10_io_out ? io_r_53_b : _GEN_2172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2174 = 8'h36 == r_count_10_io_out ? io_r_54_b : _GEN_2173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2175 = 8'h37 == r_count_10_io_out ? io_r_55_b : _GEN_2174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2176 = 8'h38 == r_count_10_io_out ? io_r_56_b : _GEN_2175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2177 = 8'h39 == r_count_10_io_out ? io_r_57_b : _GEN_2176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2178 = 8'h3a == r_count_10_io_out ? io_r_58_b : _GEN_2177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2179 = 8'h3b == r_count_10_io_out ? io_r_59_b : _GEN_2178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2180 = 8'h3c == r_count_10_io_out ? io_r_60_b : _GEN_2179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2181 = 8'h3d == r_count_10_io_out ? io_r_61_b : _GEN_2180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2182 = 8'h3e == r_count_10_io_out ? io_r_62_b : _GEN_2181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2183 = 8'h3f == r_count_10_io_out ? io_r_63_b : _GEN_2182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2184 = 8'h40 == r_count_10_io_out ? io_r_64_b : _GEN_2183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2185 = 8'h41 == r_count_10_io_out ? io_r_65_b : _GEN_2184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2186 = 8'h42 == r_count_10_io_out ? io_r_66_b : _GEN_2185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2187 = 8'h43 == r_count_10_io_out ? io_r_67_b : _GEN_2186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2188 = 8'h44 == r_count_10_io_out ? io_r_68_b : _GEN_2187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2189 = 8'h45 == r_count_10_io_out ? io_r_69_b : _GEN_2188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2190 = 8'h46 == r_count_10_io_out ? io_r_70_b : _GEN_2189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2191 = 8'h47 == r_count_10_io_out ? io_r_71_b : _GEN_2190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2192 = 8'h48 == r_count_10_io_out ? io_r_72_b : _GEN_2191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2193 = 8'h49 == r_count_10_io_out ? io_r_73_b : _GEN_2192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2194 = 8'h4a == r_count_10_io_out ? io_r_74_b : _GEN_2193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2195 = 8'h4b == r_count_10_io_out ? io_r_75_b : _GEN_2194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2196 = 8'h4c == r_count_10_io_out ? io_r_76_b : _GEN_2195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2197 = 8'h4d == r_count_10_io_out ? io_r_77_b : _GEN_2196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2198 = 8'h4e == r_count_10_io_out ? io_r_78_b : _GEN_2197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2199 = 8'h4f == r_count_10_io_out ? io_r_79_b : _GEN_2198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2200 = 8'h50 == r_count_10_io_out ? io_r_80_b : _GEN_2199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2201 = 8'h51 == r_count_10_io_out ? io_r_81_b : _GEN_2200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2202 = 8'h52 == r_count_10_io_out ? io_r_82_b : _GEN_2201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2203 = 8'h53 == r_count_10_io_out ? io_r_83_b : _GEN_2202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2204 = 8'h54 == r_count_10_io_out ? io_r_84_b : _GEN_2203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2205 = 8'h55 == r_count_10_io_out ? io_r_85_b : _GEN_2204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2206 = 8'h56 == r_count_10_io_out ? io_r_86_b : _GEN_2205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2207 = 8'h57 == r_count_10_io_out ? io_r_87_b : _GEN_2206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2208 = 8'h58 == r_count_10_io_out ? io_r_88_b : _GEN_2207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2209 = 8'h59 == r_count_10_io_out ? io_r_89_b : _GEN_2208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2210 = 8'h5a == r_count_10_io_out ? io_r_90_b : _GEN_2209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2211 = 8'h5b == r_count_10_io_out ? io_r_91_b : _GEN_2210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2212 = 8'h5c == r_count_10_io_out ? io_r_92_b : _GEN_2211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2213 = 8'h5d == r_count_10_io_out ? io_r_93_b : _GEN_2212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2214 = 8'h5e == r_count_10_io_out ? io_r_94_b : _GEN_2213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2215 = 8'h5f == r_count_10_io_out ? io_r_95_b : _GEN_2214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2216 = 8'h60 == r_count_10_io_out ? io_r_96_b : _GEN_2215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2217 = 8'h61 == r_count_10_io_out ? io_r_97_b : _GEN_2216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2218 = 8'h62 == r_count_10_io_out ? io_r_98_b : _GEN_2217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2219 = 8'h63 == r_count_10_io_out ? io_r_99_b : _GEN_2218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2220 = 8'h64 == r_count_10_io_out ? io_r_100_b : _GEN_2219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2221 = 8'h65 == r_count_10_io_out ? io_r_101_b : _GEN_2220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2222 = 8'h66 == r_count_10_io_out ? io_r_102_b : _GEN_2221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2223 = 8'h67 == r_count_10_io_out ? io_r_103_b : _GEN_2222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2224 = 8'h68 == r_count_10_io_out ? io_r_104_b : _GEN_2223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2225 = 8'h69 == r_count_10_io_out ? io_r_105_b : _GEN_2224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2226 = 8'h6a == r_count_10_io_out ? io_r_106_b : _GEN_2225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2227 = 8'h6b == r_count_10_io_out ? io_r_107_b : _GEN_2226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2228 = 8'h6c == r_count_10_io_out ? io_r_108_b : _GEN_2227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2229 = 8'h6d == r_count_10_io_out ? io_r_109_b : _GEN_2228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2230 = 8'h6e == r_count_10_io_out ? io_r_110_b : _GEN_2229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2231 = 8'h6f == r_count_10_io_out ? io_r_111_b : _GEN_2230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2232 = 8'h70 == r_count_10_io_out ? io_r_112_b : _GEN_2231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2233 = 8'h71 == r_count_10_io_out ? io_r_113_b : _GEN_2232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2234 = 8'h72 == r_count_10_io_out ? io_r_114_b : _GEN_2233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2235 = 8'h73 == r_count_10_io_out ? io_r_115_b : _GEN_2234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2236 = 8'h74 == r_count_10_io_out ? io_r_116_b : _GEN_2235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2237 = 8'h75 == r_count_10_io_out ? io_r_117_b : _GEN_2236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2238 = 8'h76 == r_count_10_io_out ? io_r_118_b : _GEN_2237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2239 = 8'h77 == r_count_10_io_out ? io_r_119_b : _GEN_2238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2240 = 8'h78 == r_count_10_io_out ? io_r_120_b : _GEN_2239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2241 = 8'h79 == r_count_10_io_out ? io_r_121_b : _GEN_2240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2242 = 8'h7a == r_count_10_io_out ? io_r_122_b : _GEN_2241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2243 = 8'h7b == r_count_10_io_out ? io_r_123_b : _GEN_2242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2244 = 8'h7c == r_count_10_io_out ? io_r_124_b : _GEN_2243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2245 = 8'h7d == r_count_10_io_out ? io_r_125_b : _GEN_2244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2246 = 8'h7e == r_count_10_io_out ? io_r_126_b : _GEN_2245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2247 = 8'h7f == r_count_10_io_out ? io_r_127_b : _GEN_2246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2248 = 8'h80 == r_count_10_io_out ? io_r_128_b : _GEN_2247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2249 = 8'h81 == r_count_10_io_out ? io_r_129_b : _GEN_2248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2250 = 8'h82 == r_count_10_io_out ? io_r_130_b : _GEN_2249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2251 = 8'h83 == r_count_10_io_out ? io_r_131_b : _GEN_2250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2252 = 8'h84 == r_count_10_io_out ? io_r_132_b : _GEN_2251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2253 = 8'h85 == r_count_10_io_out ? io_r_133_b : _GEN_2252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2254 = 8'h86 == r_count_10_io_out ? io_r_134_b : _GEN_2253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2255 = 8'h87 == r_count_10_io_out ? io_r_135_b : _GEN_2254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2256 = 8'h88 == r_count_10_io_out ? io_r_136_b : _GEN_2255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2257 = 8'h89 == r_count_10_io_out ? io_r_137_b : _GEN_2256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2258 = 8'h8a == r_count_10_io_out ? io_r_138_b : _GEN_2257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2259 = 8'h8b == r_count_10_io_out ? io_r_139_b : _GEN_2258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2260 = 8'h8c == r_count_10_io_out ? io_r_140_b : _GEN_2259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2261 = 8'h8d == r_count_10_io_out ? io_r_141_b : _GEN_2260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2262 = 8'h8e == r_count_10_io_out ? io_r_142_b : _GEN_2261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2263 = 8'h8f == r_count_10_io_out ? io_r_143_b : _GEN_2262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2264 = 8'h90 == r_count_10_io_out ? io_r_144_b : _GEN_2263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2265 = 8'h91 == r_count_10_io_out ? io_r_145_b : _GEN_2264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2266 = 8'h92 == r_count_10_io_out ? io_r_146_b : _GEN_2265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2267 = 8'h93 == r_count_10_io_out ? io_r_147_b : _GEN_2266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2268 = 8'h94 == r_count_10_io_out ? io_r_148_b : _GEN_2267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2269 = 8'h95 == r_count_10_io_out ? io_r_149_b : _GEN_2268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2270 = 8'h96 == r_count_10_io_out ? io_r_150_b : _GEN_2269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2271 = 8'h97 == r_count_10_io_out ? io_r_151_b : _GEN_2270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2272 = 8'h98 == r_count_10_io_out ? io_r_152_b : _GEN_2271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2273 = 8'h99 == r_count_10_io_out ? io_r_153_b : _GEN_2272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2274 = 8'h9a == r_count_10_io_out ? io_r_154_b : _GEN_2273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2275 = 8'h9b == r_count_10_io_out ? io_r_155_b : _GEN_2274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2276 = 8'h9c == r_count_10_io_out ? io_r_156_b : _GEN_2275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2277 = 8'h9d == r_count_10_io_out ? io_r_157_b : _GEN_2276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2278 = 8'h9e == r_count_10_io_out ? io_r_158_b : _GEN_2277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2279 = 8'h9f == r_count_10_io_out ? io_r_159_b : _GEN_2278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2280 = 8'ha0 == r_count_10_io_out ? io_r_160_b : _GEN_2279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2281 = 8'ha1 == r_count_10_io_out ? io_r_161_b : _GEN_2280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2282 = 8'ha2 == r_count_10_io_out ? io_r_162_b : _GEN_2281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2283 = 8'ha3 == r_count_10_io_out ? io_r_163_b : _GEN_2282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2284 = 8'ha4 == r_count_10_io_out ? io_r_164_b : _GEN_2283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2285 = 8'ha5 == r_count_10_io_out ? io_r_165_b : _GEN_2284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2286 = 8'ha6 == r_count_10_io_out ? io_r_166_b : _GEN_2285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2287 = 8'ha7 == r_count_10_io_out ? io_r_167_b : _GEN_2286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2288 = 8'ha8 == r_count_10_io_out ? io_r_168_b : _GEN_2287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2289 = 8'ha9 == r_count_10_io_out ? io_r_169_b : _GEN_2288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2290 = 8'haa == r_count_10_io_out ? io_r_170_b : _GEN_2289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2291 = 8'hab == r_count_10_io_out ? io_r_171_b : _GEN_2290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2292 = 8'hac == r_count_10_io_out ? io_r_172_b : _GEN_2291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2293 = 8'had == r_count_10_io_out ? io_r_173_b : _GEN_2292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2294 = 8'hae == r_count_10_io_out ? io_r_174_b : _GEN_2293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2295 = 8'haf == r_count_10_io_out ? io_r_175_b : _GEN_2294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2296 = 8'hb0 == r_count_10_io_out ? io_r_176_b : _GEN_2295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2297 = 8'hb1 == r_count_10_io_out ? io_r_177_b : _GEN_2296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2298 = 8'hb2 == r_count_10_io_out ? io_r_178_b : _GEN_2297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2299 = 8'hb3 == r_count_10_io_out ? io_r_179_b : _GEN_2298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2300 = 8'hb4 == r_count_10_io_out ? io_r_180_b : _GEN_2299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2301 = 8'hb5 == r_count_10_io_out ? io_r_181_b : _GEN_2300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2302 = 8'hb6 == r_count_10_io_out ? io_r_182_b : _GEN_2301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2303 = 8'hb7 == r_count_10_io_out ? io_r_183_b : _GEN_2302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2304 = 8'hb8 == r_count_10_io_out ? io_r_184_b : _GEN_2303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2305 = 8'hb9 == r_count_10_io_out ? io_r_185_b : _GEN_2304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2306 = 8'hba == r_count_10_io_out ? io_r_186_b : _GEN_2305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2307 = 8'hbb == r_count_10_io_out ? io_r_187_b : _GEN_2306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2308 = 8'hbc == r_count_10_io_out ? io_r_188_b : _GEN_2307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2309 = 8'hbd == r_count_10_io_out ? io_r_189_b : _GEN_2308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2310 = 8'hbe == r_count_10_io_out ? io_r_190_b : _GEN_2309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2311 = 8'hbf == r_count_10_io_out ? io_r_191_b : _GEN_2310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2312 = 8'hc0 == r_count_10_io_out ? io_r_192_b : _GEN_2311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2313 = 8'hc1 == r_count_10_io_out ? io_r_193_b : _GEN_2312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2314 = 8'hc2 == r_count_10_io_out ? io_r_194_b : _GEN_2313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2315 = 8'hc3 == r_count_10_io_out ? io_r_195_b : _GEN_2314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2316 = 8'hc4 == r_count_10_io_out ? io_r_196_b : _GEN_2315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2317 = 8'hc5 == r_count_10_io_out ? io_r_197_b : _GEN_2316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2318 = 8'hc6 == r_count_10_io_out ? io_r_198_b : _GEN_2317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2321 = 8'h1 == r_count_11_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2322 = 8'h2 == r_count_11_io_out ? io_r_2_b : _GEN_2321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2323 = 8'h3 == r_count_11_io_out ? io_r_3_b : _GEN_2322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2324 = 8'h4 == r_count_11_io_out ? io_r_4_b : _GEN_2323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2325 = 8'h5 == r_count_11_io_out ? io_r_5_b : _GEN_2324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2326 = 8'h6 == r_count_11_io_out ? io_r_6_b : _GEN_2325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2327 = 8'h7 == r_count_11_io_out ? io_r_7_b : _GEN_2326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2328 = 8'h8 == r_count_11_io_out ? io_r_8_b : _GEN_2327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2329 = 8'h9 == r_count_11_io_out ? io_r_9_b : _GEN_2328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2330 = 8'ha == r_count_11_io_out ? io_r_10_b : _GEN_2329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2331 = 8'hb == r_count_11_io_out ? io_r_11_b : _GEN_2330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2332 = 8'hc == r_count_11_io_out ? io_r_12_b : _GEN_2331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2333 = 8'hd == r_count_11_io_out ? io_r_13_b : _GEN_2332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2334 = 8'he == r_count_11_io_out ? io_r_14_b : _GEN_2333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2335 = 8'hf == r_count_11_io_out ? io_r_15_b : _GEN_2334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2336 = 8'h10 == r_count_11_io_out ? io_r_16_b : _GEN_2335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2337 = 8'h11 == r_count_11_io_out ? io_r_17_b : _GEN_2336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2338 = 8'h12 == r_count_11_io_out ? io_r_18_b : _GEN_2337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2339 = 8'h13 == r_count_11_io_out ? io_r_19_b : _GEN_2338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2340 = 8'h14 == r_count_11_io_out ? io_r_20_b : _GEN_2339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2341 = 8'h15 == r_count_11_io_out ? io_r_21_b : _GEN_2340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2342 = 8'h16 == r_count_11_io_out ? io_r_22_b : _GEN_2341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2343 = 8'h17 == r_count_11_io_out ? io_r_23_b : _GEN_2342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2344 = 8'h18 == r_count_11_io_out ? io_r_24_b : _GEN_2343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2345 = 8'h19 == r_count_11_io_out ? io_r_25_b : _GEN_2344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2346 = 8'h1a == r_count_11_io_out ? io_r_26_b : _GEN_2345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2347 = 8'h1b == r_count_11_io_out ? io_r_27_b : _GEN_2346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2348 = 8'h1c == r_count_11_io_out ? io_r_28_b : _GEN_2347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2349 = 8'h1d == r_count_11_io_out ? io_r_29_b : _GEN_2348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2350 = 8'h1e == r_count_11_io_out ? io_r_30_b : _GEN_2349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2351 = 8'h1f == r_count_11_io_out ? io_r_31_b : _GEN_2350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2352 = 8'h20 == r_count_11_io_out ? io_r_32_b : _GEN_2351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2353 = 8'h21 == r_count_11_io_out ? io_r_33_b : _GEN_2352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2354 = 8'h22 == r_count_11_io_out ? io_r_34_b : _GEN_2353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2355 = 8'h23 == r_count_11_io_out ? io_r_35_b : _GEN_2354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2356 = 8'h24 == r_count_11_io_out ? io_r_36_b : _GEN_2355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2357 = 8'h25 == r_count_11_io_out ? io_r_37_b : _GEN_2356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2358 = 8'h26 == r_count_11_io_out ? io_r_38_b : _GEN_2357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2359 = 8'h27 == r_count_11_io_out ? io_r_39_b : _GEN_2358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2360 = 8'h28 == r_count_11_io_out ? io_r_40_b : _GEN_2359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2361 = 8'h29 == r_count_11_io_out ? io_r_41_b : _GEN_2360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2362 = 8'h2a == r_count_11_io_out ? io_r_42_b : _GEN_2361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2363 = 8'h2b == r_count_11_io_out ? io_r_43_b : _GEN_2362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2364 = 8'h2c == r_count_11_io_out ? io_r_44_b : _GEN_2363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2365 = 8'h2d == r_count_11_io_out ? io_r_45_b : _GEN_2364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2366 = 8'h2e == r_count_11_io_out ? io_r_46_b : _GEN_2365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2367 = 8'h2f == r_count_11_io_out ? io_r_47_b : _GEN_2366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2368 = 8'h30 == r_count_11_io_out ? io_r_48_b : _GEN_2367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2369 = 8'h31 == r_count_11_io_out ? io_r_49_b : _GEN_2368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2370 = 8'h32 == r_count_11_io_out ? io_r_50_b : _GEN_2369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2371 = 8'h33 == r_count_11_io_out ? io_r_51_b : _GEN_2370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2372 = 8'h34 == r_count_11_io_out ? io_r_52_b : _GEN_2371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2373 = 8'h35 == r_count_11_io_out ? io_r_53_b : _GEN_2372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2374 = 8'h36 == r_count_11_io_out ? io_r_54_b : _GEN_2373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2375 = 8'h37 == r_count_11_io_out ? io_r_55_b : _GEN_2374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2376 = 8'h38 == r_count_11_io_out ? io_r_56_b : _GEN_2375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2377 = 8'h39 == r_count_11_io_out ? io_r_57_b : _GEN_2376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2378 = 8'h3a == r_count_11_io_out ? io_r_58_b : _GEN_2377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2379 = 8'h3b == r_count_11_io_out ? io_r_59_b : _GEN_2378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2380 = 8'h3c == r_count_11_io_out ? io_r_60_b : _GEN_2379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2381 = 8'h3d == r_count_11_io_out ? io_r_61_b : _GEN_2380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2382 = 8'h3e == r_count_11_io_out ? io_r_62_b : _GEN_2381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2383 = 8'h3f == r_count_11_io_out ? io_r_63_b : _GEN_2382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2384 = 8'h40 == r_count_11_io_out ? io_r_64_b : _GEN_2383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2385 = 8'h41 == r_count_11_io_out ? io_r_65_b : _GEN_2384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2386 = 8'h42 == r_count_11_io_out ? io_r_66_b : _GEN_2385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2387 = 8'h43 == r_count_11_io_out ? io_r_67_b : _GEN_2386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2388 = 8'h44 == r_count_11_io_out ? io_r_68_b : _GEN_2387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2389 = 8'h45 == r_count_11_io_out ? io_r_69_b : _GEN_2388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2390 = 8'h46 == r_count_11_io_out ? io_r_70_b : _GEN_2389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2391 = 8'h47 == r_count_11_io_out ? io_r_71_b : _GEN_2390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2392 = 8'h48 == r_count_11_io_out ? io_r_72_b : _GEN_2391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2393 = 8'h49 == r_count_11_io_out ? io_r_73_b : _GEN_2392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2394 = 8'h4a == r_count_11_io_out ? io_r_74_b : _GEN_2393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2395 = 8'h4b == r_count_11_io_out ? io_r_75_b : _GEN_2394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2396 = 8'h4c == r_count_11_io_out ? io_r_76_b : _GEN_2395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2397 = 8'h4d == r_count_11_io_out ? io_r_77_b : _GEN_2396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2398 = 8'h4e == r_count_11_io_out ? io_r_78_b : _GEN_2397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2399 = 8'h4f == r_count_11_io_out ? io_r_79_b : _GEN_2398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2400 = 8'h50 == r_count_11_io_out ? io_r_80_b : _GEN_2399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2401 = 8'h51 == r_count_11_io_out ? io_r_81_b : _GEN_2400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2402 = 8'h52 == r_count_11_io_out ? io_r_82_b : _GEN_2401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2403 = 8'h53 == r_count_11_io_out ? io_r_83_b : _GEN_2402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2404 = 8'h54 == r_count_11_io_out ? io_r_84_b : _GEN_2403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2405 = 8'h55 == r_count_11_io_out ? io_r_85_b : _GEN_2404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2406 = 8'h56 == r_count_11_io_out ? io_r_86_b : _GEN_2405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2407 = 8'h57 == r_count_11_io_out ? io_r_87_b : _GEN_2406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2408 = 8'h58 == r_count_11_io_out ? io_r_88_b : _GEN_2407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2409 = 8'h59 == r_count_11_io_out ? io_r_89_b : _GEN_2408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2410 = 8'h5a == r_count_11_io_out ? io_r_90_b : _GEN_2409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2411 = 8'h5b == r_count_11_io_out ? io_r_91_b : _GEN_2410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2412 = 8'h5c == r_count_11_io_out ? io_r_92_b : _GEN_2411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2413 = 8'h5d == r_count_11_io_out ? io_r_93_b : _GEN_2412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2414 = 8'h5e == r_count_11_io_out ? io_r_94_b : _GEN_2413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2415 = 8'h5f == r_count_11_io_out ? io_r_95_b : _GEN_2414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2416 = 8'h60 == r_count_11_io_out ? io_r_96_b : _GEN_2415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2417 = 8'h61 == r_count_11_io_out ? io_r_97_b : _GEN_2416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2418 = 8'h62 == r_count_11_io_out ? io_r_98_b : _GEN_2417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2419 = 8'h63 == r_count_11_io_out ? io_r_99_b : _GEN_2418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2420 = 8'h64 == r_count_11_io_out ? io_r_100_b : _GEN_2419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2421 = 8'h65 == r_count_11_io_out ? io_r_101_b : _GEN_2420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2422 = 8'h66 == r_count_11_io_out ? io_r_102_b : _GEN_2421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2423 = 8'h67 == r_count_11_io_out ? io_r_103_b : _GEN_2422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2424 = 8'h68 == r_count_11_io_out ? io_r_104_b : _GEN_2423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2425 = 8'h69 == r_count_11_io_out ? io_r_105_b : _GEN_2424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2426 = 8'h6a == r_count_11_io_out ? io_r_106_b : _GEN_2425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2427 = 8'h6b == r_count_11_io_out ? io_r_107_b : _GEN_2426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2428 = 8'h6c == r_count_11_io_out ? io_r_108_b : _GEN_2427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2429 = 8'h6d == r_count_11_io_out ? io_r_109_b : _GEN_2428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2430 = 8'h6e == r_count_11_io_out ? io_r_110_b : _GEN_2429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2431 = 8'h6f == r_count_11_io_out ? io_r_111_b : _GEN_2430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2432 = 8'h70 == r_count_11_io_out ? io_r_112_b : _GEN_2431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2433 = 8'h71 == r_count_11_io_out ? io_r_113_b : _GEN_2432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2434 = 8'h72 == r_count_11_io_out ? io_r_114_b : _GEN_2433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2435 = 8'h73 == r_count_11_io_out ? io_r_115_b : _GEN_2434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2436 = 8'h74 == r_count_11_io_out ? io_r_116_b : _GEN_2435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2437 = 8'h75 == r_count_11_io_out ? io_r_117_b : _GEN_2436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2438 = 8'h76 == r_count_11_io_out ? io_r_118_b : _GEN_2437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2439 = 8'h77 == r_count_11_io_out ? io_r_119_b : _GEN_2438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2440 = 8'h78 == r_count_11_io_out ? io_r_120_b : _GEN_2439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2441 = 8'h79 == r_count_11_io_out ? io_r_121_b : _GEN_2440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2442 = 8'h7a == r_count_11_io_out ? io_r_122_b : _GEN_2441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2443 = 8'h7b == r_count_11_io_out ? io_r_123_b : _GEN_2442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2444 = 8'h7c == r_count_11_io_out ? io_r_124_b : _GEN_2443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2445 = 8'h7d == r_count_11_io_out ? io_r_125_b : _GEN_2444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2446 = 8'h7e == r_count_11_io_out ? io_r_126_b : _GEN_2445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2447 = 8'h7f == r_count_11_io_out ? io_r_127_b : _GEN_2446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2448 = 8'h80 == r_count_11_io_out ? io_r_128_b : _GEN_2447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2449 = 8'h81 == r_count_11_io_out ? io_r_129_b : _GEN_2448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2450 = 8'h82 == r_count_11_io_out ? io_r_130_b : _GEN_2449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2451 = 8'h83 == r_count_11_io_out ? io_r_131_b : _GEN_2450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2452 = 8'h84 == r_count_11_io_out ? io_r_132_b : _GEN_2451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2453 = 8'h85 == r_count_11_io_out ? io_r_133_b : _GEN_2452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2454 = 8'h86 == r_count_11_io_out ? io_r_134_b : _GEN_2453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2455 = 8'h87 == r_count_11_io_out ? io_r_135_b : _GEN_2454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2456 = 8'h88 == r_count_11_io_out ? io_r_136_b : _GEN_2455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2457 = 8'h89 == r_count_11_io_out ? io_r_137_b : _GEN_2456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2458 = 8'h8a == r_count_11_io_out ? io_r_138_b : _GEN_2457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2459 = 8'h8b == r_count_11_io_out ? io_r_139_b : _GEN_2458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2460 = 8'h8c == r_count_11_io_out ? io_r_140_b : _GEN_2459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2461 = 8'h8d == r_count_11_io_out ? io_r_141_b : _GEN_2460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2462 = 8'h8e == r_count_11_io_out ? io_r_142_b : _GEN_2461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2463 = 8'h8f == r_count_11_io_out ? io_r_143_b : _GEN_2462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2464 = 8'h90 == r_count_11_io_out ? io_r_144_b : _GEN_2463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2465 = 8'h91 == r_count_11_io_out ? io_r_145_b : _GEN_2464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2466 = 8'h92 == r_count_11_io_out ? io_r_146_b : _GEN_2465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2467 = 8'h93 == r_count_11_io_out ? io_r_147_b : _GEN_2466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2468 = 8'h94 == r_count_11_io_out ? io_r_148_b : _GEN_2467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2469 = 8'h95 == r_count_11_io_out ? io_r_149_b : _GEN_2468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2470 = 8'h96 == r_count_11_io_out ? io_r_150_b : _GEN_2469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2471 = 8'h97 == r_count_11_io_out ? io_r_151_b : _GEN_2470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2472 = 8'h98 == r_count_11_io_out ? io_r_152_b : _GEN_2471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2473 = 8'h99 == r_count_11_io_out ? io_r_153_b : _GEN_2472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2474 = 8'h9a == r_count_11_io_out ? io_r_154_b : _GEN_2473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2475 = 8'h9b == r_count_11_io_out ? io_r_155_b : _GEN_2474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2476 = 8'h9c == r_count_11_io_out ? io_r_156_b : _GEN_2475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2477 = 8'h9d == r_count_11_io_out ? io_r_157_b : _GEN_2476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2478 = 8'h9e == r_count_11_io_out ? io_r_158_b : _GEN_2477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2479 = 8'h9f == r_count_11_io_out ? io_r_159_b : _GEN_2478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2480 = 8'ha0 == r_count_11_io_out ? io_r_160_b : _GEN_2479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2481 = 8'ha1 == r_count_11_io_out ? io_r_161_b : _GEN_2480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2482 = 8'ha2 == r_count_11_io_out ? io_r_162_b : _GEN_2481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2483 = 8'ha3 == r_count_11_io_out ? io_r_163_b : _GEN_2482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2484 = 8'ha4 == r_count_11_io_out ? io_r_164_b : _GEN_2483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2485 = 8'ha5 == r_count_11_io_out ? io_r_165_b : _GEN_2484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2486 = 8'ha6 == r_count_11_io_out ? io_r_166_b : _GEN_2485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2487 = 8'ha7 == r_count_11_io_out ? io_r_167_b : _GEN_2486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2488 = 8'ha8 == r_count_11_io_out ? io_r_168_b : _GEN_2487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2489 = 8'ha9 == r_count_11_io_out ? io_r_169_b : _GEN_2488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2490 = 8'haa == r_count_11_io_out ? io_r_170_b : _GEN_2489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2491 = 8'hab == r_count_11_io_out ? io_r_171_b : _GEN_2490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2492 = 8'hac == r_count_11_io_out ? io_r_172_b : _GEN_2491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2493 = 8'had == r_count_11_io_out ? io_r_173_b : _GEN_2492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2494 = 8'hae == r_count_11_io_out ? io_r_174_b : _GEN_2493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2495 = 8'haf == r_count_11_io_out ? io_r_175_b : _GEN_2494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2496 = 8'hb0 == r_count_11_io_out ? io_r_176_b : _GEN_2495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2497 = 8'hb1 == r_count_11_io_out ? io_r_177_b : _GEN_2496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2498 = 8'hb2 == r_count_11_io_out ? io_r_178_b : _GEN_2497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2499 = 8'hb3 == r_count_11_io_out ? io_r_179_b : _GEN_2498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2500 = 8'hb4 == r_count_11_io_out ? io_r_180_b : _GEN_2499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2501 = 8'hb5 == r_count_11_io_out ? io_r_181_b : _GEN_2500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2502 = 8'hb6 == r_count_11_io_out ? io_r_182_b : _GEN_2501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2503 = 8'hb7 == r_count_11_io_out ? io_r_183_b : _GEN_2502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2504 = 8'hb8 == r_count_11_io_out ? io_r_184_b : _GEN_2503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2505 = 8'hb9 == r_count_11_io_out ? io_r_185_b : _GEN_2504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2506 = 8'hba == r_count_11_io_out ? io_r_186_b : _GEN_2505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2507 = 8'hbb == r_count_11_io_out ? io_r_187_b : _GEN_2506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2508 = 8'hbc == r_count_11_io_out ? io_r_188_b : _GEN_2507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2509 = 8'hbd == r_count_11_io_out ? io_r_189_b : _GEN_2508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2510 = 8'hbe == r_count_11_io_out ? io_r_190_b : _GEN_2509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2511 = 8'hbf == r_count_11_io_out ? io_r_191_b : _GEN_2510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2512 = 8'hc0 == r_count_11_io_out ? io_r_192_b : _GEN_2511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2513 = 8'hc1 == r_count_11_io_out ? io_r_193_b : _GEN_2512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2514 = 8'hc2 == r_count_11_io_out ? io_r_194_b : _GEN_2513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2515 = 8'hc3 == r_count_11_io_out ? io_r_195_b : _GEN_2514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2516 = 8'hc4 == r_count_11_io_out ? io_r_196_b : _GEN_2515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2517 = 8'hc5 == r_count_11_io_out ? io_r_197_b : _GEN_2516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2518 = 8'hc6 == r_count_11_io_out ? io_r_198_b : _GEN_2517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2521 = 8'h1 == r_count_12_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2522 = 8'h2 == r_count_12_io_out ? io_r_2_b : _GEN_2521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2523 = 8'h3 == r_count_12_io_out ? io_r_3_b : _GEN_2522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2524 = 8'h4 == r_count_12_io_out ? io_r_4_b : _GEN_2523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2525 = 8'h5 == r_count_12_io_out ? io_r_5_b : _GEN_2524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2526 = 8'h6 == r_count_12_io_out ? io_r_6_b : _GEN_2525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2527 = 8'h7 == r_count_12_io_out ? io_r_7_b : _GEN_2526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2528 = 8'h8 == r_count_12_io_out ? io_r_8_b : _GEN_2527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2529 = 8'h9 == r_count_12_io_out ? io_r_9_b : _GEN_2528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2530 = 8'ha == r_count_12_io_out ? io_r_10_b : _GEN_2529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2531 = 8'hb == r_count_12_io_out ? io_r_11_b : _GEN_2530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2532 = 8'hc == r_count_12_io_out ? io_r_12_b : _GEN_2531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2533 = 8'hd == r_count_12_io_out ? io_r_13_b : _GEN_2532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2534 = 8'he == r_count_12_io_out ? io_r_14_b : _GEN_2533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2535 = 8'hf == r_count_12_io_out ? io_r_15_b : _GEN_2534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2536 = 8'h10 == r_count_12_io_out ? io_r_16_b : _GEN_2535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2537 = 8'h11 == r_count_12_io_out ? io_r_17_b : _GEN_2536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2538 = 8'h12 == r_count_12_io_out ? io_r_18_b : _GEN_2537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2539 = 8'h13 == r_count_12_io_out ? io_r_19_b : _GEN_2538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2540 = 8'h14 == r_count_12_io_out ? io_r_20_b : _GEN_2539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2541 = 8'h15 == r_count_12_io_out ? io_r_21_b : _GEN_2540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2542 = 8'h16 == r_count_12_io_out ? io_r_22_b : _GEN_2541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2543 = 8'h17 == r_count_12_io_out ? io_r_23_b : _GEN_2542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2544 = 8'h18 == r_count_12_io_out ? io_r_24_b : _GEN_2543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2545 = 8'h19 == r_count_12_io_out ? io_r_25_b : _GEN_2544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2546 = 8'h1a == r_count_12_io_out ? io_r_26_b : _GEN_2545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2547 = 8'h1b == r_count_12_io_out ? io_r_27_b : _GEN_2546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2548 = 8'h1c == r_count_12_io_out ? io_r_28_b : _GEN_2547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2549 = 8'h1d == r_count_12_io_out ? io_r_29_b : _GEN_2548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2550 = 8'h1e == r_count_12_io_out ? io_r_30_b : _GEN_2549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2551 = 8'h1f == r_count_12_io_out ? io_r_31_b : _GEN_2550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2552 = 8'h20 == r_count_12_io_out ? io_r_32_b : _GEN_2551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2553 = 8'h21 == r_count_12_io_out ? io_r_33_b : _GEN_2552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2554 = 8'h22 == r_count_12_io_out ? io_r_34_b : _GEN_2553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2555 = 8'h23 == r_count_12_io_out ? io_r_35_b : _GEN_2554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2556 = 8'h24 == r_count_12_io_out ? io_r_36_b : _GEN_2555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2557 = 8'h25 == r_count_12_io_out ? io_r_37_b : _GEN_2556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2558 = 8'h26 == r_count_12_io_out ? io_r_38_b : _GEN_2557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2559 = 8'h27 == r_count_12_io_out ? io_r_39_b : _GEN_2558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2560 = 8'h28 == r_count_12_io_out ? io_r_40_b : _GEN_2559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2561 = 8'h29 == r_count_12_io_out ? io_r_41_b : _GEN_2560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2562 = 8'h2a == r_count_12_io_out ? io_r_42_b : _GEN_2561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2563 = 8'h2b == r_count_12_io_out ? io_r_43_b : _GEN_2562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2564 = 8'h2c == r_count_12_io_out ? io_r_44_b : _GEN_2563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2565 = 8'h2d == r_count_12_io_out ? io_r_45_b : _GEN_2564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2566 = 8'h2e == r_count_12_io_out ? io_r_46_b : _GEN_2565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2567 = 8'h2f == r_count_12_io_out ? io_r_47_b : _GEN_2566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2568 = 8'h30 == r_count_12_io_out ? io_r_48_b : _GEN_2567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2569 = 8'h31 == r_count_12_io_out ? io_r_49_b : _GEN_2568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2570 = 8'h32 == r_count_12_io_out ? io_r_50_b : _GEN_2569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2571 = 8'h33 == r_count_12_io_out ? io_r_51_b : _GEN_2570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2572 = 8'h34 == r_count_12_io_out ? io_r_52_b : _GEN_2571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2573 = 8'h35 == r_count_12_io_out ? io_r_53_b : _GEN_2572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2574 = 8'h36 == r_count_12_io_out ? io_r_54_b : _GEN_2573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2575 = 8'h37 == r_count_12_io_out ? io_r_55_b : _GEN_2574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2576 = 8'h38 == r_count_12_io_out ? io_r_56_b : _GEN_2575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2577 = 8'h39 == r_count_12_io_out ? io_r_57_b : _GEN_2576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2578 = 8'h3a == r_count_12_io_out ? io_r_58_b : _GEN_2577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2579 = 8'h3b == r_count_12_io_out ? io_r_59_b : _GEN_2578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2580 = 8'h3c == r_count_12_io_out ? io_r_60_b : _GEN_2579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2581 = 8'h3d == r_count_12_io_out ? io_r_61_b : _GEN_2580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2582 = 8'h3e == r_count_12_io_out ? io_r_62_b : _GEN_2581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2583 = 8'h3f == r_count_12_io_out ? io_r_63_b : _GEN_2582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2584 = 8'h40 == r_count_12_io_out ? io_r_64_b : _GEN_2583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2585 = 8'h41 == r_count_12_io_out ? io_r_65_b : _GEN_2584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2586 = 8'h42 == r_count_12_io_out ? io_r_66_b : _GEN_2585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2587 = 8'h43 == r_count_12_io_out ? io_r_67_b : _GEN_2586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2588 = 8'h44 == r_count_12_io_out ? io_r_68_b : _GEN_2587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2589 = 8'h45 == r_count_12_io_out ? io_r_69_b : _GEN_2588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2590 = 8'h46 == r_count_12_io_out ? io_r_70_b : _GEN_2589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2591 = 8'h47 == r_count_12_io_out ? io_r_71_b : _GEN_2590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2592 = 8'h48 == r_count_12_io_out ? io_r_72_b : _GEN_2591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2593 = 8'h49 == r_count_12_io_out ? io_r_73_b : _GEN_2592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2594 = 8'h4a == r_count_12_io_out ? io_r_74_b : _GEN_2593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2595 = 8'h4b == r_count_12_io_out ? io_r_75_b : _GEN_2594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2596 = 8'h4c == r_count_12_io_out ? io_r_76_b : _GEN_2595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2597 = 8'h4d == r_count_12_io_out ? io_r_77_b : _GEN_2596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2598 = 8'h4e == r_count_12_io_out ? io_r_78_b : _GEN_2597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2599 = 8'h4f == r_count_12_io_out ? io_r_79_b : _GEN_2598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2600 = 8'h50 == r_count_12_io_out ? io_r_80_b : _GEN_2599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2601 = 8'h51 == r_count_12_io_out ? io_r_81_b : _GEN_2600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2602 = 8'h52 == r_count_12_io_out ? io_r_82_b : _GEN_2601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2603 = 8'h53 == r_count_12_io_out ? io_r_83_b : _GEN_2602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2604 = 8'h54 == r_count_12_io_out ? io_r_84_b : _GEN_2603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2605 = 8'h55 == r_count_12_io_out ? io_r_85_b : _GEN_2604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2606 = 8'h56 == r_count_12_io_out ? io_r_86_b : _GEN_2605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2607 = 8'h57 == r_count_12_io_out ? io_r_87_b : _GEN_2606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2608 = 8'h58 == r_count_12_io_out ? io_r_88_b : _GEN_2607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2609 = 8'h59 == r_count_12_io_out ? io_r_89_b : _GEN_2608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2610 = 8'h5a == r_count_12_io_out ? io_r_90_b : _GEN_2609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2611 = 8'h5b == r_count_12_io_out ? io_r_91_b : _GEN_2610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2612 = 8'h5c == r_count_12_io_out ? io_r_92_b : _GEN_2611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2613 = 8'h5d == r_count_12_io_out ? io_r_93_b : _GEN_2612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2614 = 8'h5e == r_count_12_io_out ? io_r_94_b : _GEN_2613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2615 = 8'h5f == r_count_12_io_out ? io_r_95_b : _GEN_2614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2616 = 8'h60 == r_count_12_io_out ? io_r_96_b : _GEN_2615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2617 = 8'h61 == r_count_12_io_out ? io_r_97_b : _GEN_2616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2618 = 8'h62 == r_count_12_io_out ? io_r_98_b : _GEN_2617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2619 = 8'h63 == r_count_12_io_out ? io_r_99_b : _GEN_2618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2620 = 8'h64 == r_count_12_io_out ? io_r_100_b : _GEN_2619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2621 = 8'h65 == r_count_12_io_out ? io_r_101_b : _GEN_2620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2622 = 8'h66 == r_count_12_io_out ? io_r_102_b : _GEN_2621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2623 = 8'h67 == r_count_12_io_out ? io_r_103_b : _GEN_2622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2624 = 8'h68 == r_count_12_io_out ? io_r_104_b : _GEN_2623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2625 = 8'h69 == r_count_12_io_out ? io_r_105_b : _GEN_2624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2626 = 8'h6a == r_count_12_io_out ? io_r_106_b : _GEN_2625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2627 = 8'h6b == r_count_12_io_out ? io_r_107_b : _GEN_2626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2628 = 8'h6c == r_count_12_io_out ? io_r_108_b : _GEN_2627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2629 = 8'h6d == r_count_12_io_out ? io_r_109_b : _GEN_2628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2630 = 8'h6e == r_count_12_io_out ? io_r_110_b : _GEN_2629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2631 = 8'h6f == r_count_12_io_out ? io_r_111_b : _GEN_2630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2632 = 8'h70 == r_count_12_io_out ? io_r_112_b : _GEN_2631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2633 = 8'h71 == r_count_12_io_out ? io_r_113_b : _GEN_2632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2634 = 8'h72 == r_count_12_io_out ? io_r_114_b : _GEN_2633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2635 = 8'h73 == r_count_12_io_out ? io_r_115_b : _GEN_2634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2636 = 8'h74 == r_count_12_io_out ? io_r_116_b : _GEN_2635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2637 = 8'h75 == r_count_12_io_out ? io_r_117_b : _GEN_2636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2638 = 8'h76 == r_count_12_io_out ? io_r_118_b : _GEN_2637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2639 = 8'h77 == r_count_12_io_out ? io_r_119_b : _GEN_2638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2640 = 8'h78 == r_count_12_io_out ? io_r_120_b : _GEN_2639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2641 = 8'h79 == r_count_12_io_out ? io_r_121_b : _GEN_2640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2642 = 8'h7a == r_count_12_io_out ? io_r_122_b : _GEN_2641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2643 = 8'h7b == r_count_12_io_out ? io_r_123_b : _GEN_2642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2644 = 8'h7c == r_count_12_io_out ? io_r_124_b : _GEN_2643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2645 = 8'h7d == r_count_12_io_out ? io_r_125_b : _GEN_2644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2646 = 8'h7e == r_count_12_io_out ? io_r_126_b : _GEN_2645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2647 = 8'h7f == r_count_12_io_out ? io_r_127_b : _GEN_2646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2648 = 8'h80 == r_count_12_io_out ? io_r_128_b : _GEN_2647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2649 = 8'h81 == r_count_12_io_out ? io_r_129_b : _GEN_2648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2650 = 8'h82 == r_count_12_io_out ? io_r_130_b : _GEN_2649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2651 = 8'h83 == r_count_12_io_out ? io_r_131_b : _GEN_2650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2652 = 8'h84 == r_count_12_io_out ? io_r_132_b : _GEN_2651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2653 = 8'h85 == r_count_12_io_out ? io_r_133_b : _GEN_2652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2654 = 8'h86 == r_count_12_io_out ? io_r_134_b : _GEN_2653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2655 = 8'h87 == r_count_12_io_out ? io_r_135_b : _GEN_2654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2656 = 8'h88 == r_count_12_io_out ? io_r_136_b : _GEN_2655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2657 = 8'h89 == r_count_12_io_out ? io_r_137_b : _GEN_2656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2658 = 8'h8a == r_count_12_io_out ? io_r_138_b : _GEN_2657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2659 = 8'h8b == r_count_12_io_out ? io_r_139_b : _GEN_2658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2660 = 8'h8c == r_count_12_io_out ? io_r_140_b : _GEN_2659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2661 = 8'h8d == r_count_12_io_out ? io_r_141_b : _GEN_2660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2662 = 8'h8e == r_count_12_io_out ? io_r_142_b : _GEN_2661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2663 = 8'h8f == r_count_12_io_out ? io_r_143_b : _GEN_2662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2664 = 8'h90 == r_count_12_io_out ? io_r_144_b : _GEN_2663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2665 = 8'h91 == r_count_12_io_out ? io_r_145_b : _GEN_2664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2666 = 8'h92 == r_count_12_io_out ? io_r_146_b : _GEN_2665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2667 = 8'h93 == r_count_12_io_out ? io_r_147_b : _GEN_2666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2668 = 8'h94 == r_count_12_io_out ? io_r_148_b : _GEN_2667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2669 = 8'h95 == r_count_12_io_out ? io_r_149_b : _GEN_2668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2670 = 8'h96 == r_count_12_io_out ? io_r_150_b : _GEN_2669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2671 = 8'h97 == r_count_12_io_out ? io_r_151_b : _GEN_2670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2672 = 8'h98 == r_count_12_io_out ? io_r_152_b : _GEN_2671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2673 = 8'h99 == r_count_12_io_out ? io_r_153_b : _GEN_2672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2674 = 8'h9a == r_count_12_io_out ? io_r_154_b : _GEN_2673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2675 = 8'h9b == r_count_12_io_out ? io_r_155_b : _GEN_2674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2676 = 8'h9c == r_count_12_io_out ? io_r_156_b : _GEN_2675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2677 = 8'h9d == r_count_12_io_out ? io_r_157_b : _GEN_2676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2678 = 8'h9e == r_count_12_io_out ? io_r_158_b : _GEN_2677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2679 = 8'h9f == r_count_12_io_out ? io_r_159_b : _GEN_2678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2680 = 8'ha0 == r_count_12_io_out ? io_r_160_b : _GEN_2679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2681 = 8'ha1 == r_count_12_io_out ? io_r_161_b : _GEN_2680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2682 = 8'ha2 == r_count_12_io_out ? io_r_162_b : _GEN_2681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2683 = 8'ha3 == r_count_12_io_out ? io_r_163_b : _GEN_2682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2684 = 8'ha4 == r_count_12_io_out ? io_r_164_b : _GEN_2683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2685 = 8'ha5 == r_count_12_io_out ? io_r_165_b : _GEN_2684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2686 = 8'ha6 == r_count_12_io_out ? io_r_166_b : _GEN_2685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2687 = 8'ha7 == r_count_12_io_out ? io_r_167_b : _GEN_2686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2688 = 8'ha8 == r_count_12_io_out ? io_r_168_b : _GEN_2687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2689 = 8'ha9 == r_count_12_io_out ? io_r_169_b : _GEN_2688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2690 = 8'haa == r_count_12_io_out ? io_r_170_b : _GEN_2689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2691 = 8'hab == r_count_12_io_out ? io_r_171_b : _GEN_2690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2692 = 8'hac == r_count_12_io_out ? io_r_172_b : _GEN_2691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2693 = 8'had == r_count_12_io_out ? io_r_173_b : _GEN_2692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2694 = 8'hae == r_count_12_io_out ? io_r_174_b : _GEN_2693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2695 = 8'haf == r_count_12_io_out ? io_r_175_b : _GEN_2694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2696 = 8'hb0 == r_count_12_io_out ? io_r_176_b : _GEN_2695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2697 = 8'hb1 == r_count_12_io_out ? io_r_177_b : _GEN_2696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2698 = 8'hb2 == r_count_12_io_out ? io_r_178_b : _GEN_2697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2699 = 8'hb3 == r_count_12_io_out ? io_r_179_b : _GEN_2698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2700 = 8'hb4 == r_count_12_io_out ? io_r_180_b : _GEN_2699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2701 = 8'hb5 == r_count_12_io_out ? io_r_181_b : _GEN_2700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2702 = 8'hb6 == r_count_12_io_out ? io_r_182_b : _GEN_2701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2703 = 8'hb7 == r_count_12_io_out ? io_r_183_b : _GEN_2702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2704 = 8'hb8 == r_count_12_io_out ? io_r_184_b : _GEN_2703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2705 = 8'hb9 == r_count_12_io_out ? io_r_185_b : _GEN_2704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2706 = 8'hba == r_count_12_io_out ? io_r_186_b : _GEN_2705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2707 = 8'hbb == r_count_12_io_out ? io_r_187_b : _GEN_2706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2708 = 8'hbc == r_count_12_io_out ? io_r_188_b : _GEN_2707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2709 = 8'hbd == r_count_12_io_out ? io_r_189_b : _GEN_2708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2710 = 8'hbe == r_count_12_io_out ? io_r_190_b : _GEN_2709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2711 = 8'hbf == r_count_12_io_out ? io_r_191_b : _GEN_2710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2712 = 8'hc0 == r_count_12_io_out ? io_r_192_b : _GEN_2711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2713 = 8'hc1 == r_count_12_io_out ? io_r_193_b : _GEN_2712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2714 = 8'hc2 == r_count_12_io_out ? io_r_194_b : _GEN_2713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2715 = 8'hc3 == r_count_12_io_out ? io_r_195_b : _GEN_2714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2716 = 8'hc4 == r_count_12_io_out ? io_r_196_b : _GEN_2715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2717 = 8'hc5 == r_count_12_io_out ? io_r_197_b : _GEN_2716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2718 = 8'hc6 == r_count_12_io_out ? io_r_198_b : _GEN_2717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2721 = 8'h1 == r_count_13_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2722 = 8'h2 == r_count_13_io_out ? io_r_2_b : _GEN_2721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2723 = 8'h3 == r_count_13_io_out ? io_r_3_b : _GEN_2722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2724 = 8'h4 == r_count_13_io_out ? io_r_4_b : _GEN_2723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2725 = 8'h5 == r_count_13_io_out ? io_r_5_b : _GEN_2724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2726 = 8'h6 == r_count_13_io_out ? io_r_6_b : _GEN_2725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2727 = 8'h7 == r_count_13_io_out ? io_r_7_b : _GEN_2726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2728 = 8'h8 == r_count_13_io_out ? io_r_8_b : _GEN_2727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2729 = 8'h9 == r_count_13_io_out ? io_r_9_b : _GEN_2728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2730 = 8'ha == r_count_13_io_out ? io_r_10_b : _GEN_2729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2731 = 8'hb == r_count_13_io_out ? io_r_11_b : _GEN_2730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2732 = 8'hc == r_count_13_io_out ? io_r_12_b : _GEN_2731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2733 = 8'hd == r_count_13_io_out ? io_r_13_b : _GEN_2732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2734 = 8'he == r_count_13_io_out ? io_r_14_b : _GEN_2733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2735 = 8'hf == r_count_13_io_out ? io_r_15_b : _GEN_2734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2736 = 8'h10 == r_count_13_io_out ? io_r_16_b : _GEN_2735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2737 = 8'h11 == r_count_13_io_out ? io_r_17_b : _GEN_2736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2738 = 8'h12 == r_count_13_io_out ? io_r_18_b : _GEN_2737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2739 = 8'h13 == r_count_13_io_out ? io_r_19_b : _GEN_2738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2740 = 8'h14 == r_count_13_io_out ? io_r_20_b : _GEN_2739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2741 = 8'h15 == r_count_13_io_out ? io_r_21_b : _GEN_2740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2742 = 8'h16 == r_count_13_io_out ? io_r_22_b : _GEN_2741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2743 = 8'h17 == r_count_13_io_out ? io_r_23_b : _GEN_2742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2744 = 8'h18 == r_count_13_io_out ? io_r_24_b : _GEN_2743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2745 = 8'h19 == r_count_13_io_out ? io_r_25_b : _GEN_2744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2746 = 8'h1a == r_count_13_io_out ? io_r_26_b : _GEN_2745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2747 = 8'h1b == r_count_13_io_out ? io_r_27_b : _GEN_2746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2748 = 8'h1c == r_count_13_io_out ? io_r_28_b : _GEN_2747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2749 = 8'h1d == r_count_13_io_out ? io_r_29_b : _GEN_2748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2750 = 8'h1e == r_count_13_io_out ? io_r_30_b : _GEN_2749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2751 = 8'h1f == r_count_13_io_out ? io_r_31_b : _GEN_2750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2752 = 8'h20 == r_count_13_io_out ? io_r_32_b : _GEN_2751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2753 = 8'h21 == r_count_13_io_out ? io_r_33_b : _GEN_2752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2754 = 8'h22 == r_count_13_io_out ? io_r_34_b : _GEN_2753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2755 = 8'h23 == r_count_13_io_out ? io_r_35_b : _GEN_2754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2756 = 8'h24 == r_count_13_io_out ? io_r_36_b : _GEN_2755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2757 = 8'h25 == r_count_13_io_out ? io_r_37_b : _GEN_2756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2758 = 8'h26 == r_count_13_io_out ? io_r_38_b : _GEN_2757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2759 = 8'h27 == r_count_13_io_out ? io_r_39_b : _GEN_2758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2760 = 8'h28 == r_count_13_io_out ? io_r_40_b : _GEN_2759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2761 = 8'h29 == r_count_13_io_out ? io_r_41_b : _GEN_2760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2762 = 8'h2a == r_count_13_io_out ? io_r_42_b : _GEN_2761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2763 = 8'h2b == r_count_13_io_out ? io_r_43_b : _GEN_2762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2764 = 8'h2c == r_count_13_io_out ? io_r_44_b : _GEN_2763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2765 = 8'h2d == r_count_13_io_out ? io_r_45_b : _GEN_2764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2766 = 8'h2e == r_count_13_io_out ? io_r_46_b : _GEN_2765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2767 = 8'h2f == r_count_13_io_out ? io_r_47_b : _GEN_2766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2768 = 8'h30 == r_count_13_io_out ? io_r_48_b : _GEN_2767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2769 = 8'h31 == r_count_13_io_out ? io_r_49_b : _GEN_2768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2770 = 8'h32 == r_count_13_io_out ? io_r_50_b : _GEN_2769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2771 = 8'h33 == r_count_13_io_out ? io_r_51_b : _GEN_2770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2772 = 8'h34 == r_count_13_io_out ? io_r_52_b : _GEN_2771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2773 = 8'h35 == r_count_13_io_out ? io_r_53_b : _GEN_2772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2774 = 8'h36 == r_count_13_io_out ? io_r_54_b : _GEN_2773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2775 = 8'h37 == r_count_13_io_out ? io_r_55_b : _GEN_2774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2776 = 8'h38 == r_count_13_io_out ? io_r_56_b : _GEN_2775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2777 = 8'h39 == r_count_13_io_out ? io_r_57_b : _GEN_2776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2778 = 8'h3a == r_count_13_io_out ? io_r_58_b : _GEN_2777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2779 = 8'h3b == r_count_13_io_out ? io_r_59_b : _GEN_2778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2780 = 8'h3c == r_count_13_io_out ? io_r_60_b : _GEN_2779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2781 = 8'h3d == r_count_13_io_out ? io_r_61_b : _GEN_2780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2782 = 8'h3e == r_count_13_io_out ? io_r_62_b : _GEN_2781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2783 = 8'h3f == r_count_13_io_out ? io_r_63_b : _GEN_2782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2784 = 8'h40 == r_count_13_io_out ? io_r_64_b : _GEN_2783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2785 = 8'h41 == r_count_13_io_out ? io_r_65_b : _GEN_2784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2786 = 8'h42 == r_count_13_io_out ? io_r_66_b : _GEN_2785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2787 = 8'h43 == r_count_13_io_out ? io_r_67_b : _GEN_2786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2788 = 8'h44 == r_count_13_io_out ? io_r_68_b : _GEN_2787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2789 = 8'h45 == r_count_13_io_out ? io_r_69_b : _GEN_2788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2790 = 8'h46 == r_count_13_io_out ? io_r_70_b : _GEN_2789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2791 = 8'h47 == r_count_13_io_out ? io_r_71_b : _GEN_2790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2792 = 8'h48 == r_count_13_io_out ? io_r_72_b : _GEN_2791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2793 = 8'h49 == r_count_13_io_out ? io_r_73_b : _GEN_2792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2794 = 8'h4a == r_count_13_io_out ? io_r_74_b : _GEN_2793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2795 = 8'h4b == r_count_13_io_out ? io_r_75_b : _GEN_2794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2796 = 8'h4c == r_count_13_io_out ? io_r_76_b : _GEN_2795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2797 = 8'h4d == r_count_13_io_out ? io_r_77_b : _GEN_2796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2798 = 8'h4e == r_count_13_io_out ? io_r_78_b : _GEN_2797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2799 = 8'h4f == r_count_13_io_out ? io_r_79_b : _GEN_2798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2800 = 8'h50 == r_count_13_io_out ? io_r_80_b : _GEN_2799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2801 = 8'h51 == r_count_13_io_out ? io_r_81_b : _GEN_2800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2802 = 8'h52 == r_count_13_io_out ? io_r_82_b : _GEN_2801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2803 = 8'h53 == r_count_13_io_out ? io_r_83_b : _GEN_2802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2804 = 8'h54 == r_count_13_io_out ? io_r_84_b : _GEN_2803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2805 = 8'h55 == r_count_13_io_out ? io_r_85_b : _GEN_2804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2806 = 8'h56 == r_count_13_io_out ? io_r_86_b : _GEN_2805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2807 = 8'h57 == r_count_13_io_out ? io_r_87_b : _GEN_2806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2808 = 8'h58 == r_count_13_io_out ? io_r_88_b : _GEN_2807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2809 = 8'h59 == r_count_13_io_out ? io_r_89_b : _GEN_2808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2810 = 8'h5a == r_count_13_io_out ? io_r_90_b : _GEN_2809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2811 = 8'h5b == r_count_13_io_out ? io_r_91_b : _GEN_2810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2812 = 8'h5c == r_count_13_io_out ? io_r_92_b : _GEN_2811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2813 = 8'h5d == r_count_13_io_out ? io_r_93_b : _GEN_2812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2814 = 8'h5e == r_count_13_io_out ? io_r_94_b : _GEN_2813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2815 = 8'h5f == r_count_13_io_out ? io_r_95_b : _GEN_2814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2816 = 8'h60 == r_count_13_io_out ? io_r_96_b : _GEN_2815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2817 = 8'h61 == r_count_13_io_out ? io_r_97_b : _GEN_2816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2818 = 8'h62 == r_count_13_io_out ? io_r_98_b : _GEN_2817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2819 = 8'h63 == r_count_13_io_out ? io_r_99_b : _GEN_2818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2820 = 8'h64 == r_count_13_io_out ? io_r_100_b : _GEN_2819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2821 = 8'h65 == r_count_13_io_out ? io_r_101_b : _GEN_2820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2822 = 8'h66 == r_count_13_io_out ? io_r_102_b : _GEN_2821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2823 = 8'h67 == r_count_13_io_out ? io_r_103_b : _GEN_2822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2824 = 8'h68 == r_count_13_io_out ? io_r_104_b : _GEN_2823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2825 = 8'h69 == r_count_13_io_out ? io_r_105_b : _GEN_2824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2826 = 8'h6a == r_count_13_io_out ? io_r_106_b : _GEN_2825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2827 = 8'h6b == r_count_13_io_out ? io_r_107_b : _GEN_2826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2828 = 8'h6c == r_count_13_io_out ? io_r_108_b : _GEN_2827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2829 = 8'h6d == r_count_13_io_out ? io_r_109_b : _GEN_2828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2830 = 8'h6e == r_count_13_io_out ? io_r_110_b : _GEN_2829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2831 = 8'h6f == r_count_13_io_out ? io_r_111_b : _GEN_2830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2832 = 8'h70 == r_count_13_io_out ? io_r_112_b : _GEN_2831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2833 = 8'h71 == r_count_13_io_out ? io_r_113_b : _GEN_2832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2834 = 8'h72 == r_count_13_io_out ? io_r_114_b : _GEN_2833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2835 = 8'h73 == r_count_13_io_out ? io_r_115_b : _GEN_2834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2836 = 8'h74 == r_count_13_io_out ? io_r_116_b : _GEN_2835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2837 = 8'h75 == r_count_13_io_out ? io_r_117_b : _GEN_2836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2838 = 8'h76 == r_count_13_io_out ? io_r_118_b : _GEN_2837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2839 = 8'h77 == r_count_13_io_out ? io_r_119_b : _GEN_2838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2840 = 8'h78 == r_count_13_io_out ? io_r_120_b : _GEN_2839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2841 = 8'h79 == r_count_13_io_out ? io_r_121_b : _GEN_2840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2842 = 8'h7a == r_count_13_io_out ? io_r_122_b : _GEN_2841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2843 = 8'h7b == r_count_13_io_out ? io_r_123_b : _GEN_2842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2844 = 8'h7c == r_count_13_io_out ? io_r_124_b : _GEN_2843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2845 = 8'h7d == r_count_13_io_out ? io_r_125_b : _GEN_2844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2846 = 8'h7e == r_count_13_io_out ? io_r_126_b : _GEN_2845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2847 = 8'h7f == r_count_13_io_out ? io_r_127_b : _GEN_2846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2848 = 8'h80 == r_count_13_io_out ? io_r_128_b : _GEN_2847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2849 = 8'h81 == r_count_13_io_out ? io_r_129_b : _GEN_2848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2850 = 8'h82 == r_count_13_io_out ? io_r_130_b : _GEN_2849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2851 = 8'h83 == r_count_13_io_out ? io_r_131_b : _GEN_2850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2852 = 8'h84 == r_count_13_io_out ? io_r_132_b : _GEN_2851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2853 = 8'h85 == r_count_13_io_out ? io_r_133_b : _GEN_2852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2854 = 8'h86 == r_count_13_io_out ? io_r_134_b : _GEN_2853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2855 = 8'h87 == r_count_13_io_out ? io_r_135_b : _GEN_2854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2856 = 8'h88 == r_count_13_io_out ? io_r_136_b : _GEN_2855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2857 = 8'h89 == r_count_13_io_out ? io_r_137_b : _GEN_2856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2858 = 8'h8a == r_count_13_io_out ? io_r_138_b : _GEN_2857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2859 = 8'h8b == r_count_13_io_out ? io_r_139_b : _GEN_2858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2860 = 8'h8c == r_count_13_io_out ? io_r_140_b : _GEN_2859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2861 = 8'h8d == r_count_13_io_out ? io_r_141_b : _GEN_2860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2862 = 8'h8e == r_count_13_io_out ? io_r_142_b : _GEN_2861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2863 = 8'h8f == r_count_13_io_out ? io_r_143_b : _GEN_2862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2864 = 8'h90 == r_count_13_io_out ? io_r_144_b : _GEN_2863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2865 = 8'h91 == r_count_13_io_out ? io_r_145_b : _GEN_2864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2866 = 8'h92 == r_count_13_io_out ? io_r_146_b : _GEN_2865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2867 = 8'h93 == r_count_13_io_out ? io_r_147_b : _GEN_2866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2868 = 8'h94 == r_count_13_io_out ? io_r_148_b : _GEN_2867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2869 = 8'h95 == r_count_13_io_out ? io_r_149_b : _GEN_2868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2870 = 8'h96 == r_count_13_io_out ? io_r_150_b : _GEN_2869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2871 = 8'h97 == r_count_13_io_out ? io_r_151_b : _GEN_2870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2872 = 8'h98 == r_count_13_io_out ? io_r_152_b : _GEN_2871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2873 = 8'h99 == r_count_13_io_out ? io_r_153_b : _GEN_2872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2874 = 8'h9a == r_count_13_io_out ? io_r_154_b : _GEN_2873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2875 = 8'h9b == r_count_13_io_out ? io_r_155_b : _GEN_2874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2876 = 8'h9c == r_count_13_io_out ? io_r_156_b : _GEN_2875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2877 = 8'h9d == r_count_13_io_out ? io_r_157_b : _GEN_2876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2878 = 8'h9e == r_count_13_io_out ? io_r_158_b : _GEN_2877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2879 = 8'h9f == r_count_13_io_out ? io_r_159_b : _GEN_2878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2880 = 8'ha0 == r_count_13_io_out ? io_r_160_b : _GEN_2879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2881 = 8'ha1 == r_count_13_io_out ? io_r_161_b : _GEN_2880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2882 = 8'ha2 == r_count_13_io_out ? io_r_162_b : _GEN_2881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2883 = 8'ha3 == r_count_13_io_out ? io_r_163_b : _GEN_2882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2884 = 8'ha4 == r_count_13_io_out ? io_r_164_b : _GEN_2883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2885 = 8'ha5 == r_count_13_io_out ? io_r_165_b : _GEN_2884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2886 = 8'ha6 == r_count_13_io_out ? io_r_166_b : _GEN_2885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2887 = 8'ha7 == r_count_13_io_out ? io_r_167_b : _GEN_2886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2888 = 8'ha8 == r_count_13_io_out ? io_r_168_b : _GEN_2887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2889 = 8'ha9 == r_count_13_io_out ? io_r_169_b : _GEN_2888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2890 = 8'haa == r_count_13_io_out ? io_r_170_b : _GEN_2889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2891 = 8'hab == r_count_13_io_out ? io_r_171_b : _GEN_2890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2892 = 8'hac == r_count_13_io_out ? io_r_172_b : _GEN_2891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2893 = 8'had == r_count_13_io_out ? io_r_173_b : _GEN_2892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2894 = 8'hae == r_count_13_io_out ? io_r_174_b : _GEN_2893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2895 = 8'haf == r_count_13_io_out ? io_r_175_b : _GEN_2894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2896 = 8'hb0 == r_count_13_io_out ? io_r_176_b : _GEN_2895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2897 = 8'hb1 == r_count_13_io_out ? io_r_177_b : _GEN_2896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2898 = 8'hb2 == r_count_13_io_out ? io_r_178_b : _GEN_2897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2899 = 8'hb3 == r_count_13_io_out ? io_r_179_b : _GEN_2898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2900 = 8'hb4 == r_count_13_io_out ? io_r_180_b : _GEN_2899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2901 = 8'hb5 == r_count_13_io_out ? io_r_181_b : _GEN_2900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2902 = 8'hb6 == r_count_13_io_out ? io_r_182_b : _GEN_2901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2903 = 8'hb7 == r_count_13_io_out ? io_r_183_b : _GEN_2902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2904 = 8'hb8 == r_count_13_io_out ? io_r_184_b : _GEN_2903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2905 = 8'hb9 == r_count_13_io_out ? io_r_185_b : _GEN_2904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2906 = 8'hba == r_count_13_io_out ? io_r_186_b : _GEN_2905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2907 = 8'hbb == r_count_13_io_out ? io_r_187_b : _GEN_2906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2908 = 8'hbc == r_count_13_io_out ? io_r_188_b : _GEN_2907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2909 = 8'hbd == r_count_13_io_out ? io_r_189_b : _GEN_2908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2910 = 8'hbe == r_count_13_io_out ? io_r_190_b : _GEN_2909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2911 = 8'hbf == r_count_13_io_out ? io_r_191_b : _GEN_2910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2912 = 8'hc0 == r_count_13_io_out ? io_r_192_b : _GEN_2911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2913 = 8'hc1 == r_count_13_io_out ? io_r_193_b : _GEN_2912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2914 = 8'hc2 == r_count_13_io_out ? io_r_194_b : _GEN_2913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2915 = 8'hc3 == r_count_13_io_out ? io_r_195_b : _GEN_2914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2916 = 8'hc4 == r_count_13_io_out ? io_r_196_b : _GEN_2915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2917 = 8'hc5 == r_count_13_io_out ? io_r_197_b : _GEN_2916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2918 = 8'hc6 == r_count_13_io_out ? io_r_198_b : _GEN_2917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2921 = 8'h1 == r_count_14_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2922 = 8'h2 == r_count_14_io_out ? io_r_2_b : _GEN_2921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2923 = 8'h3 == r_count_14_io_out ? io_r_3_b : _GEN_2922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2924 = 8'h4 == r_count_14_io_out ? io_r_4_b : _GEN_2923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2925 = 8'h5 == r_count_14_io_out ? io_r_5_b : _GEN_2924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2926 = 8'h6 == r_count_14_io_out ? io_r_6_b : _GEN_2925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2927 = 8'h7 == r_count_14_io_out ? io_r_7_b : _GEN_2926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2928 = 8'h8 == r_count_14_io_out ? io_r_8_b : _GEN_2927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2929 = 8'h9 == r_count_14_io_out ? io_r_9_b : _GEN_2928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2930 = 8'ha == r_count_14_io_out ? io_r_10_b : _GEN_2929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2931 = 8'hb == r_count_14_io_out ? io_r_11_b : _GEN_2930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2932 = 8'hc == r_count_14_io_out ? io_r_12_b : _GEN_2931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2933 = 8'hd == r_count_14_io_out ? io_r_13_b : _GEN_2932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2934 = 8'he == r_count_14_io_out ? io_r_14_b : _GEN_2933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2935 = 8'hf == r_count_14_io_out ? io_r_15_b : _GEN_2934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2936 = 8'h10 == r_count_14_io_out ? io_r_16_b : _GEN_2935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2937 = 8'h11 == r_count_14_io_out ? io_r_17_b : _GEN_2936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2938 = 8'h12 == r_count_14_io_out ? io_r_18_b : _GEN_2937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2939 = 8'h13 == r_count_14_io_out ? io_r_19_b : _GEN_2938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2940 = 8'h14 == r_count_14_io_out ? io_r_20_b : _GEN_2939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2941 = 8'h15 == r_count_14_io_out ? io_r_21_b : _GEN_2940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2942 = 8'h16 == r_count_14_io_out ? io_r_22_b : _GEN_2941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2943 = 8'h17 == r_count_14_io_out ? io_r_23_b : _GEN_2942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2944 = 8'h18 == r_count_14_io_out ? io_r_24_b : _GEN_2943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2945 = 8'h19 == r_count_14_io_out ? io_r_25_b : _GEN_2944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2946 = 8'h1a == r_count_14_io_out ? io_r_26_b : _GEN_2945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2947 = 8'h1b == r_count_14_io_out ? io_r_27_b : _GEN_2946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2948 = 8'h1c == r_count_14_io_out ? io_r_28_b : _GEN_2947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2949 = 8'h1d == r_count_14_io_out ? io_r_29_b : _GEN_2948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2950 = 8'h1e == r_count_14_io_out ? io_r_30_b : _GEN_2949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2951 = 8'h1f == r_count_14_io_out ? io_r_31_b : _GEN_2950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2952 = 8'h20 == r_count_14_io_out ? io_r_32_b : _GEN_2951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2953 = 8'h21 == r_count_14_io_out ? io_r_33_b : _GEN_2952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2954 = 8'h22 == r_count_14_io_out ? io_r_34_b : _GEN_2953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2955 = 8'h23 == r_count_14_io_out ? io_r_35_b : _GEN_2954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2956 = 8'h24 == r_count_14_io_out ? io_r_36_b : _GEN_2955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2957 = 8'h25 == r_count_14_io_out ? io_r_37_b : _GEN_2956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2958 = 8'h26 == r_count_14_io_out ? io_r_38_b : _GEN_2957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2959 = 8'h27 == r_count_14_io_out ? io_r_39_b : _GEN_2958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2960 = 8'h28 == r_count_14_io_out ? io_r_40_b : _GEN_2959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2961 = 8'h29 == r_count_14_io_out ? io_r_41_b : _GEN_2960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2962 = 8'h2a == r_count_14_io_out ? io_r_42_b : _GEN_2961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2963 = 8'h2b == r_count_14_io_out ? io_r_43_b : _GEN_2962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2964 = 8'h2c == r_count_14_io_out ? io_r_44_b : _GEN_2963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2965 = 8'h2d == r_count_14_io_out ? io_r_45_b : _GEN_2964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2966 = 8'h2e == r_count_14_io_out ? io_r_46_b : _GEN_2965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2967 = 8'h2f == r_count_14_io_out ? io_r_47_b : _GEN_2966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2968 = 8'h30 == r_count_14_io_out ? io_r_48_b : _GEN_2967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2969 = 8'h31 == r_count_14_io_out ? io_r_49_b : _GEN_2968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2970 = 8'h32 == r_count_14_io_out ? io_r_50_b : _GEN_2969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2971 = 8'h33 == r_count_14_io_out ? io_r_51_b : _GEN_2970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2972 = 8'h34 == r_count_14_io_out ? io_r_52_b : _GEN_2971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2973 = 8'h35 == r_count_14_io_out ? io_r_53_b : _GEN_2972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2974 = 8'h36 == r_count_14_io_out ? io_r_54_b : _GEN_2973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2975 = 8'h37 == r_count_14_io_out ? io_r_55_b : _GEN_2974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2976 = 8'h38 == r_count_14_io_out ? io_r_56_b : _GEN_2975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2977 = 8'h39 == r_count_14_io_out ? io_r_57_b : _GEN_2976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2978 = 8'h3a == r_count_14_io_out ? io_r_58_b : _GEN_2977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2979 = 8'h3b == r_count_14_io_out ? io_r_59_b : _GEN_2978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2980 = 8'h3c == r_count_14_io_out ? io_r_60_b : _GEN_2979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2981 = 8'h3d == r_count_14_io_out ? io_r_61_b : _GEN_2980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2982 = 8'h3e == r_count_14_io_out ? io_r_62_b : _GEN_2981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2983 = 8'h3f == r_count_14_io_out ? io_r_63_b : _GEN_2982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2984 = 8'h40 == r_count_14_io_out ? io_r_64_b : _GEN_2983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2985 = 8'h41 == r_count_14_io_out ? io_r_65_b : _GEN_2984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2986 = 8'h42 == r_count_14_io_out ? io_r_66_b : _GEN_2985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2987 = 8'h43 == r_count_14_io_out ? io_r_67_b : _GEN_2986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2988 = 8'h44 == r_count_14_io_out ? io_r_68_b : _GEN_2987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2989 = 8'h45 == r_count_14_io_out ? io_r_69_b : _GEN_2988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2990 = 8'h46 == r_count_14_io_out ? io_r_70_b : _GEN_2989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2991 = 8'h47 == r_count_14_io_out ? io_r_71_b : _GEN_2990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2992 = 8'h48 == r_count_14_io_out ? io_r_72_b : _GEN_2991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2993 = 8'h49 == r_count_14_io_out ? io_r_73_b : _GEN_2992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2994 = 8'h4a == r_count_14_io_out ? io_r_74_b : _GEN_2993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2995 = 8'h4b == r_count_14_io_out ? io_r_75_b : _GEN_2994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2996 = 8'h4c == r_count_14_io_out ? io_r_76_b : _GEN_2995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2997 = 8'h4d == r_count_14_io_out ? io_r_77_b : _GEN_2996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2998 = 8'h4e == r_count_14_io_out ? io_r_78_b : _GEN_2997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2999 = 8'h4f == r_count_14_io_out ? io_r_79_b : _GEN_2998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3000 = 8'h50 == r_count_14_io_out ? io_r_80_b : _GEN_2999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3001 = 8'h51 == r_count_14_io_out ? io_r_81_b : _GEN_3000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3002 = 8'h52 == r_count_14_io_out ? io_r_82_b : _GEN_3001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3003 = 8'h53 == r_count_14_io_out ? io_r_83_b : _GEN_3002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3004 = 8'h54 == r_count_14_io_out ? io_r_84_b : _GEN_3003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3005 = 8'h55 == r_count_14_io_out ? io_r_85_b : _GEN_3004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3006 = 8'h56 == r_count_14_io_out ? io_r_86_b : _GEN_3005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3007 = 8'h57 == r_count_14_io_out ? io_r_87_b : _GEN_3006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3008 = 8'h58 == r_count_14_io_out ? io_r_88_b : _GEN_3007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3009 = 8'h59 == r_count_14_io_out ? io_r_89_b : _GEN_3008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3010 = 8'h5a == r_count_14_io_out ? io_r_90_b : _GEN_3009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3011 = 8'h5b == r_count_14_io_out ? io_r_91_b : _GEN_3010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3012 = 8'h5c == r_count_14_io_out ? io_r_92_b : _GEN_3011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3013 = 8'h5d == r_count_14_io_out ? io_r_93_b : _GEN_3012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3014 = 8'h5e == r_count_14_io_out ? io_r_94_b : _GEN_3013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3015 = 8'h5f == r_count_14_io_out ? io_r_95_b : _GEN_3014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3016 = 8'h60 == r_count_14_io_out ? io_r_96_b : _GEN_3015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3017 = 8'h61 == r_count_14_io_out ? io_r_97_b : _GEN_3016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3018 = 8'h62 == r_count_14_io_out ? io_r_98_b : _GEN_3017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3019 = 8'h63 == r_count_14_io_out ? io_r_99_b : _GEN_3018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3020 = 8'h64 == r_count_14_io_out ? io_r_100_b : _GEN_3019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3021 = 8'h65 == r_count_14_io_out ? io_r_101_b : _GEN_3020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3022 = 8'h66 == r_count_14_io_out ? io_r_102_b : _GEN_3021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3023 = 8'h67 == r_count_14_io_out ? io_r_103_b : _GEN_3022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3024 = 8'h68 == r_count_14_io_out ? io_r_104_b : _GEN_3023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3025 = 8'h69 == r_count_14_io_out ? io_r_105_b : _GEN_3024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3026 = 8'h6a == r_count_14_io_out ? io_r_106_b : _GEN_3025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3027 = 8'h6b == r_count_14_io_out ? io_r_107_b : _GEN_3026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3028 = 8'h6c == r_count_14_io_out ? io_r_108_b : _GEN_3027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3029 = 8'h6d == r_count_14_io_out ? io_r_109_b : _GEN_3028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3030 = 8'h6e == r_count_14_io_out ? io_r_110_b : _GEN_3029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3031 = 8'h6f == r_count_14_io_out ? io_r_111_b : _GEN_3030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3032 = 8'h70 == r_count_14_io_out ? io_r_112_b : _GEN_3031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3033 = 8'h71 == r_count_14_io_out ? io_r_113_b : _GEN_3032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3034 = 8'h72 == r_count_14_io_out ? io_r_114_b : _GEN_3033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3035 = 8'h73 == r_count_14_io_out ? io_r_115_b : _GEN_3034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3036 = 8'h74 == r_count_14_io_out ? io_r_116_b : _GEN_3035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3037 = 8'h75 == r_count_14_io_out ? io_r_117_b : _GEN_3036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3038 = 8'h76 == r_count_14_io_out ? io_r_118_b : _GEN_3037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3039 = 8'h77 == r_count_14_io_out ? io_r_119_b : _GEN_3038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3040 = 8'h78 == r_count_14_io_out ? io_r_120_b : _GEN_3039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3041 = 8'h79 == r_count_14_io_out ? io_r_121_b : _GEN_3040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3042 = 8'h7a == r_count_14_io_out ? io_r_122_b : _GEN_3041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3043 = 8'h7b == r_count_14_io_out ? io_r_123_b : _GEN_3042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3044 = 8'h7c == r_count_14_io_out ? io_r_124_b : _GEN_3043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3045 = 8'h7d == r_count_14_io_out ? io_r_125_b : _GEN_3044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3046 = 8'h7e == r_count_14_io_out ? io_r_126_b : _GEN_3045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3047 = 8'h7f == r_count_14_io_out ? io_r_127_b : _GEN_3046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3048 = 8'h80 == r_count_14_io_out ? io_r_128_b : _GEN_3047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3049 = 8'h81 == r_count_14_io_out ? io_r_129_b : _GEN_3048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3050 = 8'h82 == r_count_14_io_out ? io_r_130_b : _GEN_3049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3051 = 8'h83 == r_count_14_io_out ? io_r_131_b : _GEN_3050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3052 = 8'h84 == r_count_14_io_out ? io_r_132_b : _GEN_3051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3053 = 8'h85 == r_count_14_io_out ? io_r_133_b : _GEN_3052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3054 = 8'h86 == r_count_14_io_out ? io_r_134_b : _GEN_3053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3055 = 8'h87 == r_count_14_io_out ? io_r_135_b : _GEN_3054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3056 = 8'h88 == r_count_14_io_out ? io_r_136_b : _GEN_3055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3057 = 8'h89 == r_count_14_io_out ? io_r_137_b : _GEN_3056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3058 = 8'h8a == r_count_14_io_out ? io_r_138_b : _GEN_3057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3059 = 8'h8b == r_count_14_io_out ? io_r_139_b : _GEN_3058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3060 = 8'h8c == r_count_14_io_out ? io_r_140_b : _GEN_3059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3061 = 8'h8d == r_count_14_io_out ? io_r_141_b : _GEN_3060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3062 = 8'h8e == r_count_14_io_out ? io_r_142_b : _GEN_3061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3063 = 8'h8f == r_count_14_io_out ? io_r_143_b : _GEN_3062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3064 = 8'h90 == r_count_14_io_out ? io_r_144_b : _GEN_3063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3065 = 8'h91 == r_count_14_io_out ? io_r_145_b : _GEN_3064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3066 = 8'h92 == r_count_14_io_out ? io_r_146_b : _GEN_3065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3067 = 8'h93 == r_count_14_io_out ? io_r_147_b : _GEN_3066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3068 = 8'h94 == r_count_14_io_out ? io_r_148_b : _GEN_3067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3069 = 8'h95 == r_count_14_io_out ? io_r_149_b : _GEN_3068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3070 = 8'h96 == r_count_14_io_out ? io_r_150_b : _GEN_3069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3071 = 8'h97 == r_count_14_io_out ? io_r_151_b : _GEN_3070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3072 = 8'h98 == r_count_14_io_out ? io_r_152_b : _GEN_3071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3073 = 8'h99 == r_count_14_io_out ? io_r_153_b : _GEN_3072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3074 = 8'h9a == r_count_14_io_out ? io_r_154_b : _GEN_3073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3075 = 8'h9b == r_count_14_io_out ? io_r_155_b : _GEN_3074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3076 = 8'h9c == r_count_14_io_out ? io_r_156_b : _GEN_3075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3077 = 8'h9d == r_count_14_io_out ? io_r_157_b : _GEN_3076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3078 = 8'h9e == r_count_14_io_out ? io_r_158_b : _GEN_3077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3079 = 8'h9f == r_count_14_io_out ? io_r_159_b : _GEN_3078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3080 = 8'ha0 == r_count_14_io_out ? io_r_160_b : _GEN_3079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3081 = 8'ha1 == r_count_14_io_out ? io_r_161_b : _GEN_3080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3082 = 8'ha2 == r_count_14_io_out ? io_r_162_b : _GEN_3081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3083 = 8'ha3 == r_count_14_io_out ? io_r_163_b : _GEN_3082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3084 = 8'ha4 == r_count_14_io_out ? io_r_164_b : _GEN_3083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3085 = 8'ha5 == r_count_14_io_out ? io_r_165_b : _GEN_3084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3086 = 8'ha6 == r_count_14_io_out ? io_r_166_b : _GEN_3085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3087 = 8'ha7 == r_count_14_io_out ? io_r_167_b : _GEN_3086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3088 = 8'ha8 == r_count_14_io_out ? io_r_168_b : _GEN_3087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3089 = 8'ha9 == r_count_14_io_out ? io_r_169_b : _GEN_3088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3090 = 8'haa == r_count_14_io_out ? io_r_170_b : _GEN_3089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3091 = 8'hab == r_count_14_io_out ? io_r_171_b : _GEN_3090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3092 = 8'hac == r_count_14_io_out ? io_r_172_b : _GEN_3091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3093 = 8'had == r_count_14_io_out ? io_r_173_b : _GEN_3092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3094 = 8'hae == r_count_14_io_out ? io_r_174_b : _GEN_3093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3095 = 8'haf == r_count_14_io_out ? io_r_175_b : _GEN_3094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3096 = 8'hb0 == r_count_14_io_out ? io_r_176_b : _GEN_3095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3097 = 8'hb1 == r_count_14_io_out ? io_r_177_b : _GEN_3096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3098 = 8'hb2 == r_count_14_io_out ? io_r_178_b : _GEN_3097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3099 = 8'hb3 == r_count_14_io_out ? io_r_179_b : _GEN_3098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3100 = 8'hb4 == r_count_14_io_out ? io_r_180_b : _GEN_3099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3101 = 8'hb5 == r_count_14_io_out ? io_r_181_b : _GEN_3100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3102 = 8'hb6 == r_count_14_io_out ? io_r_182_b : _GEN_3101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3103 = 8'hb7 == r_count_14_io_out ? io_r_183_b : _GEN_3102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3104 = 8'hb8 == r_count_14_io_out ? io_r_184_b : _GEN_3103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3105 = 8'hb9 == r_count_14_io_out ? io_r_185_b : _GEN_3104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3106 = 8'hba == r_count_14_io_out ? io_r_186_b : _GEN_3105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3107 = 8'hbb == r_count_14_io_out ? io_r_187_b : _GEN_3106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3108 = 8'hbc == r_count_14_io_out ? io_r_188_b : _GEN_3107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3109 = 8'hbd == r_count_14_io_out ? io_r_189_b : _GEN_3108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3110 = 8'hbe == r_count_14_io_out ? io_r_190_b : _GEN_3109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3111 = 8'hbf == r_count_14_io_out ? io_r_191_b : _GEN_3110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3112 = 8'hc0 == r_count_14_io_out ? io_r_192_b : _GEN_3111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3113 = 8'hc1 == r_count_14_io_out ? io_r_193_b : _GEN_3112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3114 = 8'hc2 == r_count_14_io_out ? io_r_194_b : _GEN_3113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3115 = 8'hc3 == r_count_14_io_out ? io_r_195_b : _GEN_3114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3116 = 8'hc4 == r_count_14_io_out ? io_r_196_b : _GEN_3115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3117 = 8'hc5 == r_count_14_io_out ? io_r_197_b : _GEN_3116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3118 = 8'hc6 == r_count_14_io_out ? io_r_198_b : _GEN_3117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3121 = 8'h1 == r_count_15_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3122 = 8'h2 == r_count_15_io_out ? io_r_2_b : _GEN_3121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3123 = 8'h3 == r_count_15_io_out ? io_r_3_b : _GEN_3122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3124 = 8'h4 == r_count_15_io_out ? io_r_4_b : _GEN_3123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3125 = 8'h5 == r_count_15_io_out ? io_r_5_b : _GEN_3124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3126 = 8'h6 == r_count_15_io_out ? io_r_6_b : _GEN_3125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3127 = 8'h7 == r_count_15_io_out ? io_r_7_b : _GEN_3126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3128 = 8'h8 == r_count_15_io_out ? io_r_8_b : _GEN_3127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3129 = 8'h9 == r_count_15_io_out ? io_r_9_b : _GEN_3128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3130 = 8'ha == r_count_15_io_out ? io_r_10_b : _GEN_3129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3131 = 8'hb == r_count_15_io_out ? io_r_11_b : _GEN_3130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3132 = 8'hc == r_count_15_io_out ? io_r_12_b : _GEN_3131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3133 = 8'hd == r_count_15_io_out ? io_r_13_b : _GEN_3132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3134 = 8'he == r_count_15_io_out ? io_r_14_b : _GEN_3133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3135 = 8'hf == r_count_15_io_out ? io_r_15_b : _GEN_3134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3136 = 8'h10 == r_count_15_io_out ? io_r_16_b : _GEN_3135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3137 = 8'h11 == r_count_15_io_out ? io_r_17_b : _GEN_3136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3138 = 8'h12 == r_count_15_io_out ? io_r_18_b : _GEN_3137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3139 = 8'h13 == r_count_15_io_out ? io_r_19_b : _GEN_3138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3140 = 8'h14 == r_count_15_io_out ? io_r_20_b : _GEN_3139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3141 = 8'h15 == r_count_15_io_out ? io_r_21_b : _GEN_3140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3142 = 8'h16 == r_count_15_io_out ? io_r_22_b : _GEN_3141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3143 = 8'h17 == r_count_15_io_out ? io_r_23_b : _GEN_3142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3144 = 8'h18 == r_count_15_io_out ? io_r_24_b : _GEN_3143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3145 = 8'h19 == r_count_15_io_out ? io_r_25_b : _GEN_3144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3146 = 8'h1a == r_count_15_io_out ? io_r_26_b : _GEN_3145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3147 = 8'h1b == r_count_15_io_out ? io_r_27_b : _GEN_3146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3148 = 8'h1c == r_count_15_io_out ? io_r_28_b : _GEN_3147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3149 = 8'h1d == r_count_15_io_out ? io_r_29_b : _GEN_3148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3150 = 8'h1e == r_count_15_io_out ? io_r_30_b : _GEN_3149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3151 = 8'h1f == r_count_15_io_out ? io_r_31_b : _GEN_3150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3152 = 8'h20 == r_count_15_io_out ? io_r_32_b : _GEN_3151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3153 = 8'h21 == r_count_15_io_out ? io_r_33_b : _GEN_3152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3154 = 8'h22 == r_count_15_io_out ? io_r_34_b : _GEN_3153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3155 = 8'h23 == r_count_15_io_out ? io_r_35_b : _GEN_3154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3156 = 8'h24 == r_count_15_io_out ? io_r_36_b : _GEN_3155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3157 = 8'h25 == r_count_15_io_out ? io_r_37_b : _GEN_3156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3158 = 8'h26 == r_count_15_io_out ? io_r_38_b : _GEN_3157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3159 = 8'h27 == r_count_15_io_out ? io_r_39_b : _GEN_3158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3160 = 8'h28 == r_count_15_io_out ? io_r_40_b : _GEN_3159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3161 = 8'h29 == r_count_15_io_out ? io_r_41_b : _GEN_3160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3162 = 8'h2a == r_count_15_io_out ? io_r_42_b : _GEN_3161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3163 = 8'h2b == r_count_15_io_out ? io_r_43_b : _GEN_3162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3164 = 8'h2c == r_count_15_io_out ? io_r_44_b : _GEN_3163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3165 = 8'h2d == r_count_15_io_out ? io_r_45_b : _GEN_3164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3166 = 8'h2e == r_count_15_io_out ? io_r_46_b : _GEN_3165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3167 = 8'h2f == r_count_15_io_out ? io_r_47_b : _GEN_3166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3168 = 8'h30 == r_count_15_io_out ? io_r_48_b : _GEN_3167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3169 = 8'h31 == r_count_15_io_out ? io_r_49_b : _GEN_3168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3170 = 8'h32 == r_count_15_io_out ? io_r_50_b : _GEN_3169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3171 = 8'h33 == r_count_15_io_out ? io_r_51_b : _GEN_3170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3172 = 8'h34 == r_count_15_io_out ? io_r_52_b : _GEN_3171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3173 = 8'h35 == r_count_15_io_out ? io_r_53_b : _GEN_3172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3174 = 8'h36 == r_count_15_io_out ? io_r_54_b : _GEN_3173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3175 = 8'h37 == r_count_15_io_out ? io_r_55_b : _GEN_3174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3176 = 8'h38 == r_count_15_io_out ? io_r_56_b : _GEN_3175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3177 = 8'h39 == r_count_15_io_out ? io_r_57_b : _GEN_3176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3178 = 8'h3a == r_count_15_io_out ? io_r_58_b : _GEN_3177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3179 = 8'h3b == r_count_15_io_out ? io_r_59_b : _GEN_3178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3180 = 8'h3c == r_count_15_io_out ? io_r_60_b : _GEN_3179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3181 = 8'h3d == r_count_15_io_out ? io_r_61_b : _GEN_3180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3182 = 8'h3e == r_count_15_io_out ? io_r_62_b : _GEN_3181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3183 = 8'h3f == r_count_15_io_out ? io_r_63_b : _GEN_3182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3184 = 8'h40 == r_count_15_io_out ? io_r_64_b : _GEN_3183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3185 = 8'h41 == r_count_15_io_out ? io_r_65_b : _GEN_3184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3186 = 8'h42 == r_count_15_io_out ? io_r_66_b : _GEN_3185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3187 = 8'h43 == r_count_15_io_out ? io_r_67_b : _GEN_3186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3188 = 8'h44 == r_count_15_io_out ? io_r_68_b : _GEN_3187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3189 = 8'h45 == r_count_15_io_out ? io_r_69_b : _GEN_3188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3190 = 8'h46 == r_count_15_io_out ? io_r_70_b : _GEN_3189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3191 = 8'h47 == r_count_15_io_out ? io_r_71_b : _GEN_3190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3192 = 8'h48 == r_count_15_io_out ? io_r_72_b : _GEN_3191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3193 = 8'h49 == r_count_15_io_out ? io_r_73_b : _GEN_3192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3194 = 8'h4a == r_count_15_io_out ? io_r_74_b : _GEN_3193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3195 = 8'h4b == r_count_15_io_out ? io_r_75_b : _GEN_3194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3196 = 8'h4c == r_count_15_io_out ? io_r_76_b : _GEN_3195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3197 = 8'h4d == r_count_15_io_out ? io_r_77_b : _GEN_3196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3198 = 8'h4e == r_count_15_io_out ? io_r_78_b : _GEN_3197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3199 = 8'h4f == r_count_15_io_out ? io_r_79_b : _GEN_3198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3200 = 8'h50 == r_count_15_io_out ? io_r_80_b : _GEN_3199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3201 = 8'h51 == r_count_15_io_out ? io_r_81_b : _GEN_3200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3202 = 8'h52 == r_count_15_io_out ? io_r_82_b : _GEN_3201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3203 = 8'h53 == r_count_15_io_out ? io_r_83_b : _GEN_3202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3204 = 8'h54 == r_count_15_io_out ? io_r_84_b : _GEN_3203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3205 = 8'h55 == r_count_15_io_out ? io_r_85_b : _GEN_3204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3206 = 8'h56 == r_count_15_io_out ? io_r_86_b : _GEN_3205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3207 = 8'h57 == r_count_15_io_out ? io_r_87_b : _GEN_3206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3208 = 8'h58 == r_count_15_io_out ? io_r_88_b : _GEN_3207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3209 = 8'h59 == r_count_15_io_out ? io_r_89_b : _GEN_3208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3210 = 8'h5a == r_count_15_io_out ? io_r_90_b : _GEN_3209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3211 = 8'h5b == r_count_15_io_out ? io_r_91_b : _GEN_3210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3212 = 8'h5c == r_count_15_io_out ? io_r_92_b : _GEN_3211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3213 = 8'h5d == r_count_15_io_out ? io_r_93_b : _GEN_3212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3214 = 8'h5e == r_count_15_io_out ? io_r_94_b : _GEN_3213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3215 = 8'h5f == r_count_15_io_out ? io_r_95_b : _GEN_3214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3216 = 8'h60 == r_count_15_io_out ? io_r_96_b : _GEN_3215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3217 = 8'h61 == r_count_15_io_out ? io_r_97_b : _GEN_3216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3218 = 8'h62 == r_count_15_io_out ? io_r_98_b : _GEN_3217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3219 = 8'h63 == r_count_15_io_out ? io_r_99_b : _GEN_3218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3220 = 8'h64 == r_count_15_io_out ? io_r_100_b : _GEN_3219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3221 = 8'h65 == r_count_15_io_out ? io_r_101_b : _GEN_3220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3222 = 8'h66 == r_count_15_io_out ? io_r_102_b : _GEN_3221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3223 = 8'h67 == r_count_15_io_out ? io_r_103_b : _GEN_3222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3224 = 8'h68 == r_count_15_io_out ? io_r_104_b : _GEN_3223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3225 = 8'h69 == r_count_15_io_out ? io_r_105_b : _GEN_3224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3226 = 8'h6a == r_count_15_io_out ? io_r_106_b : _GEN_3225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3227 = 8'h6b == r_count_15_io_out ? io_r_107_b : _GEN_3226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3228 = 8'h6c == r_count_15_io_out ? io_r_108_b : _GEN_3227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3229 = 8'h6d == r_count_15_io_out ? io_r_109_b : _GEN_3228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3230 = 8'h6e == r_count_15_io_out ? io_r_110_b : _GEN_3229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3231 = 8'h6f == r_count_15_io_out ? io_r_111_b : _GEN_3230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3232 = 8'h70 == r_count_15_io_out ? io_r_112_b : _GEN_3231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3233 = 8'h71 == r_count_15_io_out ? io_r_113_b : _GEN_3232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3234 = 8'h72 == r_count_15_io_out ? io_r_114_b : _GEN_3233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3235 = 8'h73 == r_count_15_io_out ? io_r_115_b : _GEN_3234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3236 = 8'h74 == r_count_15_io_out ? io_r_116_b : _GEN_3235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3237 = 8'h75 == r_count_15_io_out ? io_r_117_b : _GEN_3236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3238 = 8'h76 == r_count_15_io_out ? io_r_118_b : _GEN_3237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3239 = 8'h77 == r_count_15_io_out ? io_r_119_b : _GEN_3238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3240 = 8'h78 == r_count_15_io_out ? io_r_120_b : _GEN_3239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3241 = 8'h79 == r_count_15_io_out ? io_r_121_b : _GEN_3240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3242 = 8'h7a == r_count_15_io_out ? io_r_122_b : _GEN_3241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3243 = 8'h7b == r_count_15_io_out ? io_r_123_b : _GEN_3242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3244 = 8'h7c == r_count_15_io_out ? io_r_124_b : _GEN_3243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3245 = 8'h7d == r_count_15_io_out ? io_r_125_b : _GEN_3244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3246 = 8'h7e == r_count_15_io_out ? io_r_126_b : _GEN_3245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3247 = 8'h7f == r_count_15_io_out ? io_r_127_b : _GEN_3246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3248 = 8'h80 == r_count_15_io_out ? io_r_128_b : _GEN_3247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3249 = 8'h81 == r_count_15_io_out ? io_r_129_b : _GEN_3248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3250 = 8'h82 == r_count_15_io_out ? io_r_130_b : _GEN_3249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3251 = 8'h83 == r_count_15_io_out ? io_r_131_b : _GEN_3250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3252 = 8'h84 == r_count_15_io_out ? io_r_132_b : _GEN_3251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3253 = 8'h85 == r_count_15_io_out ? io_r_133_b : _GEN_3252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3254 = 8'h86 == r_count_15_io_out ? io_r_134_b : _GEN_3253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3255 = 8'h87 == r_count_15_io_out ? io_r_135_b : _GEN_3254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3256 = 8'h88 == r_count_15_io_out ? io_r_136_b : _GEN_3255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3257 = 8'h89 == r_count_15_io_out ? io_r_137_b : _GEN_3256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3258 = 8'h8a == r_count_15_io_out ? io_r_138_b : _GEN_3257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3259 = 8'h8b == r_count_15_io_out ? io_r_139_b : _GEN_3258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3260 = 8'h8c == r_count_15_io_out ? io_r_140_b : _GEN_3259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3261 = 8'h8d == r_count_15_io_out ? io_r_141_b : _GEN_3260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3262 = 8'h8e == r_count_15_io_out ? io_r_142_b : _GEN_3261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3263 = 8'h8f == r_count_15_io_out ? io_r_143_b : _GEN_3262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3264 = 8'h90 == r_count_15_io_out ? io_r_144_b : _GEN_3263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3265 = 8'h91 == r_count_15_io_out ? io_r_145_b : _GEN_3264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3266 = 8'h92 == r_count_15_io_out ? io_r_146_b : _GEN_3265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3267 = 8'h93 == r_count_15_io_out ? io_r_147_b : _GEN_3266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3268 = 8'h94 == r_count_15_io_out ? io_r_148_b : _GEN_3267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3269 = 8'h95 == r_count_15_io_out ? io_r_149_b : _GEN_3268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3270 = 8'h96 == r_count_15_io_out ? io_r_150_b : _GEN_3269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3271 = 8'h97 == r_count_15_io_out ? io_r_151_b : _GEN_3270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3272 = 8'h98 == r_count_15_io_out ? io_r_152_b : _GEN_3271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3273 = 8'h99 == r_count_15_io_out ? io_r_153_b : _GEN_3272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3274 = 8'h9a == r_count_15_io_out ? io_r_154_b : _GEN_3273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3275 = 8'h9b == r_count_15_io_out ? io_r_155_b : _GEN_3274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3276 = 8'h9c == r_count_15_io_out ? io_r_156_b : _GEN_3275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3277 = 8'h9d == r_count_15_io_out ? io_r_157_b : _GEN_3276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3278 = 8'h9e == r_count_15_io_out ? io_r_158_b : _GEN_3277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3279 = 8'h9f == r_count_15_io_out ? io_r_159_b : _GEN_3278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3280 = 8'ha0 == r_count_15_io_out ? io_r_160_b : _GEN_3279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3281 = 8'ha1 == r_count_15_io_out ? io_r_161_b : _GEN_3280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3282 = 8'ha2 == r_count_15_io_out ? io_r_162_b : _GEN_3281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3283 = 8'ha3 == r_count_15_io_out ? io_r_163_b : _GEN_3282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3284 = 8'ha4 == r_count_15_io_out ? io_r_164_b : _GEN_3283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3285 = 8'ha5 == r_count_15_io_out ? io_r_165_b : _GEN_3284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3286 = 8'ha6 == r_count_15_io_out ? io_r_166_b : _GEN_3285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3287 = 8'ha7 == r_count_15_io_out ? io_r_167_b : _GEN_3286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3288 = 8'ha8 == r_count_15_io_out ? io_r_168_b : _GEN_3287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3289 = 8'ha9 == r_count_15_io_out ? io_r_169_b : _GEN_3288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3290 = 8'haa == r_count_15_io_out ? io_r_170_b : _GEN_3289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3291 = 8'hab == r_count_15_io_out ? io_r_171_b : _GEN_3290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3292 = 8'hac == r_count_15_io_out ? io_r_172_b : _GEN_3291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3293 = 8'had == r_count_15_io_out ? io_r_173_b : _GEN_3292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3294 = 8'hae == r_count_15_io_out ? io_r_174_b : _GEN_3293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3295 = 8'haf == r_count_15_io_out ? io_r_175_b : _GEN_3294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3296 = 8'hb0 == r_count_15_io_out ? io_r_176_b : _GEN_3295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3297 = 8'hb1 == r_count_15_io_out ? io_r_177_b : _GEN_3296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3298 = 8'hb2 == r_count_15_io_out ? io_r_178_b : _GEN_3297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3299 = 8'hb3 == r_count_15_io_out ? io_r_179_b : _GEN_3298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3300 = 8'hb4 == r_count_15_io_out ? io_r_180_b : _GEN_3299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3301 = 8'hb5 == r_count_15_io_out ? io_r_181_b : _GEN_3300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3302 = 8'hb6 == r_count_15_io_out ? io_r_182_b : _GEN_3301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3303 = 8'hb7 == r_count_15_io_out ? io_r_183_b : _GEN_3302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3304 = 8'hb8 == r_count_15_io_out ? io_r_184_b : _GEN_3303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3305 = 8'hb9 == r_count_15_io_out ? io_r_185_b : _GEN_3304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3306 = 8'hba == r_count_15_io_out ? io_r_186_b : _GEN_3305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3307 = 8'hbb == r_count_15_io_out ? io_r_187_b : _GEN_3306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3308 = 8'hbc == r_count_15_io_out ? io_r_188_b : _GEN_3307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3309 = 8'hbd == r_count_15_io_out ? io_r_189_b : _GEN_3308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3310 = 8'hbe == r_count_15_io_out ? io_r_190_b : _GEN_3309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3311 = 8'hbf == r_count_15_io_out ? io_r_191_b : _GEN_3310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3312 = 8'hc0 == r_count_15_io_out ? io_r_192_b : _GEN_3311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3313 = 8'hc1 == r_count_15_io_out ? io_r_193_b : _GEN_3312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3314 = 8'hc2 == r_count_15_io_out ? io_r_194_b : _GEN_3313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3315 = 8'hc3 == r_count_15_io_out ? io_r_195_b : _GEN_3314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3316 = 8'hc4 == r_count_15_io_out ? io_r_196_b : _GEN_3315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3317 = 8'hc5 == r_count_15_io_out ? io_r_197_b : _GEN_3316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3318 = 8'hc6 == r_count_15_io_out ? io_r_198_b : _GEN_3317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3321 = 8'h1 == r_count_16_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3322 = 8'h2 == r_count_16_io_out ? io_r_2_b : _GEN_3321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3323 = 8'h3 == r_count_16_io_out ? io_r_3_b : _GEN_3322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3324 = 8'h4 == r_count_16_io_out ? io_r_4_b : _GEN_3323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3325 = 8'h5 == r_count_16_io_out ? io_r_5_b : _GEN_3324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3326 = 8'h6 == r_count_16_io_out ? io_r_6_b : _GEN_3325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3327 = 8'h7 == r_count_16_io_out ? io_r_7_b : _GEN_3326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3328 = 8'h8 == r_count_16_io_out ? io_r_8_b : _GEN_3327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3329 = 8'h9 == r_count_16_io_out ? io_r_9_b : _GEN_3328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3330 = 8'ha == r_count_16_io_out ? io_r_10_b : _GEN_3329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3331 = 8'hb == r_count_16_io_out ? io_r_11_b : _GEN_3330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3332 = 8'hc == r_count_16_io_out ? io_r_12_b : _GEN_3331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3333 = 8'hd == r_count_16_io_out ? io_r_13_b : _GEN_3332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3334 = 8'he == r_count_16_io_out ? io_r_14_b : _GEN_3333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3335 = 8'hf == r_count_16_io_out ? io_r_15_b : _GEN_3334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3336 = 8'h10 == r_count_16_io_out ? io_r_16_b : _GEN_3335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3337 = 8'h11 == r_count_16_io_out ? io_r_17_b : _GEN_3336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3338 = 8'h12 == r_count_16_io_out ? io_r_18_b : _GEN_3337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3339 = 8'h13 == r_count_16_io_out ? io_r_19_b : _GEN_3338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3340 = 8'h14 == r_count_16_io_out ? io_r_20_b : _GEN_3339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3341 = 8'h15 == r_count_16_io_out ? io_r_21_b : _GEN_3340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3342 = 8'h16 == r_count_16_io_out ? io_r_22_b : _GEN_3341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3343 = 8'h17 == r_count_16_io_out ? io_r_23_b : _GEN_3342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3344 = 8'h18 == r_count_16_io_out ? io_r_24_b : _GEN_3343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3345 = 8'h19 == r_count_16_io_out ? io_r_25_b : _GEN_3344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3346 = 8'h1a == r_count_16_io_out ? io_r_26_b : _GEN_3345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3347 = 8'h1b == r_count_16_io_out ? io_r_27_b : _GEN_3346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3348 = 8'h1c == r_count_16_io_out ? io_r_28_b : _GEN_3347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3349 = 8'h1d == r_count_16_io_out ? io_r_29_b : _GEN_3348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3350 = 8'h1e == r_count_16_io_out ? io_r_30_b : _GEN_3349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3351 = 8'h1f == r_count_16_io_out ? io_r_31_b : _GEN_3350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3352 = 8'h20 == r_count_16_io_out ? io_r_32_b : _GEN_3351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3353 = 8'h21 == r_count_16_io_out ? io_r_33_b : _GEN_3352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3354 = 8'h22 == r_count_16_io_out ? io_r_34_b : _GEN_3353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3355 = 8'h23 == r_count_16_io_out ? io_r_35_b : _GEN_3354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3356 = 8'h24 == r_count_16_io_out ? io_r_36_b : _GEN_3355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3357 = 8'h25 == r_count_16_io_out ? io_r_37_b : _GEN_3356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3358 = 8'h26 == r_count_16_io_out ? io_r_38_b : _GEN_3357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3359 = 8'h27 == r_count_16_io_out ? io_r_39_b : _GEN_3358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3360 = 8'h28 == r_count_16_io_out ? io_r_40_b : _GEN_3359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3361 = 8'h29 == r_count_16_io_out ? io_r_41_b : _GEN_3360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3362 = 8'h2a == r_count_16_io_out ? io_r_42_b : _GEN_3361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3363 = 8'h2b == r_count_16_io_out ? io_r_43_b : _GEN_3362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3364 = 8'h2c == r_count_16_io_out ? io_r_44_b : _GEN_3363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3365 = 8'h2d == r_count_16_io_out ? io_r_45_b : _GEN_3364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3366 = 8'h2e == r_count_16_io_out ? io_r_46_b : _GEN_3365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3367 = 8'h2f == r_count_16_io_out ? io_r_47_b : _GEN_3366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3368 = 8'h30 == r_count_16_io_out ? io_r_48_b : _GEN_3367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3369 = 8'h31 == r_count_16_io_out ? io_r_49_b : _GEN_3368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3370 = 8'h32 == r_count_16_io_out ? io_r_50_b : _GEN_3369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3371 = 8'h33 == r_count_16_io_out ? io_r_51_b : _GEN_3370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3372 = 8'h34 == r_count_16_io_out ? io_r_52_b : _GEN_3371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3373 = 8'h35 == r_count_16_io_out ? io_r_53_b : _GEN_3372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3374 = 8'h36 == r_count_16_io_out ? io_r_54_b : _GEN_3373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3375 = 8'h37 == r_count_16_io_out ? io_r_55_b : _GEN_3374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3376 = 8'h38 == r_count_16_io_out ? io_r_56_b : _GEN_3375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3377 = 8'h39 == r_count_16_io_out ? io_r_57_b : _GEN_3376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3378 = 8'h3a == r_count_16_io_out ? io_r_58_b : _GEN_3377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3379 = 8'h3b == r_count_16_io_out ? io_r_59_b : _GEN_3378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3380 = 8'h3c == r_count_16_io_out ? io_r_60_b : _GEN_3379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3381 = 8'h3d == r_count_16_io_out ? io_r_61_b : _GEN_3380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3382 = 8'h3e == r_count_16_io_out ? io_r_62_b : _GEN_3381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3383 = 8'h3f == r_count_16_io_out ? io_r_63_b : _GEN_3382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3384 = 8'h40 == r_count_16_io_out ? io_r_64_b : _GEN_3383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3385 = 8'h41 == r_count_16_io_out ? io_r_65_b : _GEN_3384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3386 = 8'h42 == r_count_16_io_out ? io_r_66_b : _GEN_3385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3387 = 8'h43 == r_count_16_io_out ? io_r_67_b : _GEN_3386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3388 = 8'h44 == r_count_16_io_out ? io_r_68_b : _GEN_3387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3389 = 8'h45 == r_count_16_io_out ? io_r_69_b : _GEN_3388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3390 = 8'h46 == r_count_16_io_out ? io_r_70_b : _GEN_3389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3391 = 8'h47 == r_count_16_io_out ? io_r_71_b : _GEN_3390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3392 = 8'h48 == r_count_16_io_out ? io_r_72_b : _GEN_3391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3393 = 8'h49 == r_count_16_io_out ? io_r_73_b : _GEN_3392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3394 = 8'h4a == r_count_16_io_out ? io_r_74_b : _GEN_3393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3395 = 8'h4b == r_count_16_io_out ? io_r_75_b : _GEN_3394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3396 = 8'h4c == r_count_16_io_out ? io_r_76_b : _GEN_3395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3397 = 8'h4d == r_count_16_io_out ? io_r_77_b : _GEN_3396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3398 = 8'h4e == r_count_16_io_out ? io_r_78_b : _GEN_3397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3399 = 8'h4f == r_count_16_io_out ? io_r_79_b : _GEN_3398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3400 = 8'h50 == r_count_16_io_out ? io_r_80_b : _GEN_3399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3401 = 8'h51 == r_count_16_io_out ? io_r_81_b : _GEN_3400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3402 = 8'h52 == r_count_16_io_out ? io_r_82_b : _GEN_3401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3403 = 8'h53 == r_count_16_io_out ? io_r_83_b : _GEN_3402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3404 = 8'h54 == r_count_16_io_out ? io_r_84_b : _GEN_3403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3405 = 8'h55 == r_count_16_io_out ? io_r_85_b : _GEN_3404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3406 = 8'h56 == r_count_16_io_out ? io_r_86_b : _GEN_3405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3407 = 8'h57 == r_count_16_io_out ? io_r_87_b : _GEN_3406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3408 = 8'h58 == r_count_16_io_out ? io_r_88_b : _GEN_3407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3409 = 8'h59 == r_count_16_io_out ? io_r_89_b : _GEN_3408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3410 = 8'h5a == r_count_16_io_out ? io_r_90_b : _GEN_3409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3411 = 8'h5b == r_count_16_io_out ? io_r_91_b : _GEN_3410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3412 = 8'h5c == r_count_16_io_out ? io_r_92_b : _GEN_3411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3413 = 8'h5d == r_count_16_io_out ? io_r_93_b : _GEN_3412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3414 = 8'h5e == r_count_16_io_out ? io_r_94_b : _GEN_3413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3415 = 8'h5f == r_count_16_io_out ? io_r_95_b : _GEN_3414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3416 = 8'h60 == r_count_16_io_out ? io_r_96_b : _GEN_3415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3417 = 8'h61 == r_count_16_io_out ? io_r_97_b : _GEN_3416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3418 = 8'h62 == r_count_16_io_out ? io_r_98_b : _GEN_3417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3419 = 8'h63 == r_count_16_io_out ? io_r_99_b : _GEN_3418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3420 = 8'h64 == r_count_16_io_out ? io_r_100_b : _GEN_3419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3421 = 8'h65 == r_count_16_io_out ? io_r_101_b : _GEN_3420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3422 = 8'h66 == r_count_16_io_out ? io_r_102_b : _GEN_3421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3423 = 8'h67 == r_count_16_io_out ? io_r_103_b : _GEN_3422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3424 = 8'h68 == r_count_16_io_out ? io_r_104_b : _GEN_3423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3425 = 8'h69 == r_count_16_io_out ? io_r_105_b : _GEN_3424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3426 = 8'h6a == r_count_16_io_out ? io_r_106_b : _GEN_3425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3427 = 8'h6b == r_count_16_io_out ? io_r_107_b : _GEN_3426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3428 = 8'h6c == r_count_16_io_out ? io_r_108_b : _GEN_3427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3429 = 8'h6d == r_count_16_io_out ? io_r_109_b : _GEN_3428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3430 = 8'h6e == r_count_16_io_out ? io_r_110_b : _GEN_3429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3431 = 8'h6f == r_count_16_io_out ? io_r_111_b : _GEN_3430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3432 = 8'h70 == r_count_16_io_out ? io_r_112_b : _GEN_3431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3433 = 8'h71 == r_count_16_io_out ? io_r_113_b : _GEN_3432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3434 = 8'h72 == r_count_16_io_out ? io_r_114_b : _GEN_3433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3435 = 8'h73 == r_count_16_io_out ? io_r_115_b : _GEN_3434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3436 = 8'h74 == r_count_16_io_out ? io_r_116_b : _GEN_3435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3437 = 8'h75 == r_count_16_io_out ? io_r_117_b : _GEN_3436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3438 = 8'h76 == r_count_16_io_out ? io_r_118_b : _GEN_3437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3439 = 8'h77 == r_count_16_io_out ? io_r_119_b : _GEN_3438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3440 = 8'h78 == r_count_16_io_out ? io_r_120_b : _GEN_3439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3441 = 8'h79 == r_count_16_io_out ? io_r_121_b : _GEN_3440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3442 = 8'h7a == r_count_16_io_out ? io_r_122_b : _GEN_3441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3443 = 8'h7b == r_count_16_io_out ? io_r_123_b : _GEN_3442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3444 = 8'h7c == r_count_16_io_out ? io_r_124_b : _GEN_3443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3445 = 8'h7d == r_count_16_io_out ? io_r_125_b : _GEN_3444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3446 = 8'h7e == r_count_16_io_out ? io_r_126_b : _GEN_3445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3447 = 8'h7f == r_count_16_io_out ? io_r_127_b : _GEN_3446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3448 = 8'h80 == r_count_16_io_out ? io_r_128_b : _GEN_3447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3449 = 8'h81 == r_count_16_io_out ? io_r_129_b : _GEN_3448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3450 = 8'h82 == r_count_16_io_out ? io_r_130_b : _GEN_3449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3451 = 8'h83 == r_count_16_io_out ? io_r_131_b : _GEN_3450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3452 = 8'h84 == r_count_16_io_out ? io_r_132_b : _GEN_3451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3453 = 8'h85 == r_count_16_io_out ? io_r_133_b : _GEN_3452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3454 = 8'h86 == r_count_16_io_out ? io_r_134_b : _GEN_3453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3455 = 8'h87 == r_count_16_io_out ? io_r_135_b : _GEN_3454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3456 = 8'h88 == r_count_16_io_out ? io_r_136_b : _GEN_3455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3457 = 8'h89 == r_count_16_io_out ? io_r_137_b : _GEN_3456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3458 = 8'h8a == r_count_16_io_out ? io_r_138_b : _GEN_3457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3459 = 8'h8b == r_count_16_io_out ? io_r_139_b : _GEN_3458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3460 = 8'h8c == r_count_16_io_out ? io_r_140_b : _GEN_3459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3461 = 8'h8d == r_count_16_io_out ? io_r_141_b : _GEN_3460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3462 = 8'h8e == r_count_16_io_out ? io_r_142_b : _GEN_3461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3463 = 8'h8f == r_count_16_io_out ? io_r_143_b : _GEN_3462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3464 = 8'h90 == r_count_16_io_out ? io_r_144_b : _GEN_3463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3465 = 8'h91 == r_count_16_io_out ? io_r_145_b : _GEN_3464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3466 = 8'h92 == r_count_16_io_out ? io_r_146_b : _GEN_3465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3467 = 8'h93 == r_count_16_io_out ? io_r_147_b : _GEN_3466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3468 = 8'h94 == r_count_16_io_out ? io_r_148_b : _GEN_3467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3469 = 8'h95 == r_count_16_io_out ? io_r_149_b : _GEN_3468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3470 = 8'h96 == r_count_16_io_out ? io_r_150_b : _GEN_3469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3471 = 8'h97 == r_count_16_io_out ? io_r_151_b : _GEN_3470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3472 = 8'h98 == r_count_16_io_out ? io_r_152_b : _GEN_3471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3473 = 8'h99 == r_count_16_io_out ? io_r_153_b : _GEN_3472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3474 = 8'h9a == r_count_16_io_out ? io_r_154_b : _GEN_3473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3475 = 8'h9b == r_count_16_io_out ? io_r_155_b : _GEN_3474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3476 = 8'h9c == r_count_16_io_out ? io_r_156_b : _GEN_3475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3477 = 8'h9d == r_count_16_io_out ? io_r_157_b : _GEN_3476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3478 = 8'h9e == r_count_16_io_out ? io_r_158_b : _GEN_3477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3479 = 8'h9f == r_count_16_io_out ? io_r_159_b : _GEN_3478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3480 = 8'ha0 == r_count_16_io_out ? io_r_160_b : _GEN_3479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3481 = 8'ha1 == r_count_16_io_out ? io_r_161_b : _GEN_3480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3482 = 8'ha2 == r_count_16_io_out ? io_r_162_b : _GEN_3481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3483 = 8'ha3 == r_count_16_io_out ? io_r_163_b : _GEN_3482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3484 = 8'ha4 == r_count_16_io_out ? io_r_164_b : _GEN_3483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3485 = 8'ha5 == r_count_16_io_out ? io_r_165_b : _GEN_3484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3486 = 8'ha6 == r_count_16_io_out ? io_r_166_b : _GEN_3485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3487 = 8'ha7 == r_count_16_io_out ? io_r_167_b : _GEN_3486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3488 = 8'ha8 == r_count_16_io_out ? io_r_168_b : _GEN_3487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3489 = 8'ha9 == r_count_16_io_out ? io_r_169_b : _GEN_3488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3490 = 8'haa == r_count_16_io_out ? io_r_170_b : _GEN_3489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3491 = 8'hab == r_count_16_io_out ? io_r_171_b : _GEN_3490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3492 = 8'hac == r_count_16_io_out ? io_r_172_b : _GEN_3491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3493 = 8'had == r_count_16_io_out ? io_r_173_b : _GEN_3492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3494 = 8'hae == r_count_16_io_out ? io_r_174_b : _GEN_3493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3495 = 8'haf == r_count_16_io_out ? io_r_175_b : _GEN_3494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3496 = 8'hb0 == r_count_16_io_out ? io_r_176_b : _GEN_3495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3497 = 8'hb1 == r_count_16_io_out ? io_r_177_b : _GEN_3496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3498 = 8'hb2 == r_count_16_io_out ? io_r_178_b : _GEN_3497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3499 = 8'hb3 == r_count_16_io_out ? io_r_179_b : _GEN_3498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3500 = 8'hb4 == r_count_16_io_out ? io_r_180_b : _GEN_3499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3501 = 8'hb5 == r_count_16_io_out ? io_r_181_b : _GEN_3500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3502 = 8'hb6 == r_count_16_io_out ? io_r_182_b : _GEN_3501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3503 = 8'hb7 == r_count_16_io_out ? io_r_183_b : _GEN_3502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3504 = 8'hb8 == r_count_16_io_out ? io_r_184_b : _GEN_3503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3505 = 8'hb9 == r_count_16_io_out ? io_r_185_b : _GEN_3504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3506 = 8'hba == r_count_16_io_out ? io_r_186_b : _GEN_3505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3507 = 8'hbb == r_count_16_io_out ? io_r_187_b : _GEN_3506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3508 = 8'hbc == r_count_16_io_out ? io_r_188_b : _GEN_3507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3509 = 8'hbd == r_count_16_io_out ? io_r_189_b : _GEN_3508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3510 = 8'hbe == r_count_16_io_out ? io_r_190_b : _GEN_3509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3511 = 8'hbf == r_count_16_io_out ? io_r_191_b : _GEN_3510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3512 = 8'hc0 == r_count_16_io_out ? io_r_192_b : _GEN_3511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3513 = 8'hc1 == r_count_16_io_out ? io_r_193_b : _GEN_3512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3514 = 8'hc2 == r_count_16_io_out ? io_r_194_b : _GEN_3513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3515 = 8'hc3 == r_count_16_io_out ? io_r_195_b : _GEN_3514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3516 = 8'hc4 == r_count_16_io_out ? io_r_196_b : _GEN_3515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3517 = 8'hc5 == r_count_16_io_out ? io_r_197_b : _GEN_3516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3518 = 8'hc6 == r_count_16_io_out ? io_r_198_b : _GEN_3517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3521 = 8'h1 == r_count_17_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3522 = 8'h2 == r_count_17_io_out ? io_r_2_b : _GEN_3521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3523 = 8'h3 == r_count_17_io_out ? io_r_3_b : _GEN_3522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3524 = 8'h4 == r_count_17_io_out ? io_r_4_b : _GEN_3523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3525 = 8'h5 == r_count_17_io_out ? io_r_5_b : _GEN_3524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3526 = 8'h6 == r_count_17_io_out ? io_r_6_b : _GEN_3525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3527 = 8'h7 == r_count_17_io_out ? io_r_7_b : _GEN_3526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3528 = 8'h8 == r_count_17_io_out ? io_r_8_b : _GEN_3527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3529 = 8'h9 == r_count_17_io_out ? io_r_9_b : _GEN_3528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3530 = 8'ha == r_count_17_io_out ? io_r_10_b : _GEN_3529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3531 = 8'hb == r_count_17_io_out ? io_r_11_b : _GEN_3530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3532 = 8'hc == r_count_17_io_out ? io_r_12_b : _GEN_3531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3533 = 8'hd == r_count_17_io_out ? io_r_13_b : _GEN_3532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3534 = 8'he == r_count_17_io_out ? io_r_14_b : _GEN_3533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3535 = 8'hf == r_count_17_io_out ? io_r_15_b : _GEN_3534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3536 = 8'h10 == r_count_17_io_out ? io_r_16_b : _GEN_3535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3537 = 8'h11 == r_count_17_io_out ? io_r_17_b : _GEN_3536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3538 = 8'h12 == r_count_17_io_out ? io_r_18_b : _GEN_3537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3539 = 8'h13 == r_count_17_io_out ? io_r_19_b : _GEN_3538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3540 = 8'h14 == r_count_17_io_out ? io_r_20_b : _GEN_3539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3541 = 8'h15 == r_count_17_io_out ? io_r_21_b : _GEN_3540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3542 = 8'h16 == r_count_17_io_out ? io_r_22_b : _GEN_3541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3543 = 8'h17 == r_count_17_io_out ? io_r_23_b : _GEN_3542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3544 = 8'h18 == r_count_17_io_out ? io_r_24_b : _GEN_3543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3545 = 8'h19 == r_count_17_io_out ? io_r_25_b : _GEN_3544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3546 = 8'h1a == r_count_17_io_out ? io_r_26_b : _GEN_3545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3547 = 8'h1b == r_count_17_io_out ? io_r_27_b : _GEN_3546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3548 = 8'h1c == r_count_17_io_out ? io_r_28_b : _GEN_3547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3549 = 8'h1d == r_count_17_io_out ? io_r_29_b : _GEN_3548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3550 = 8'h1e == r_count_17_io_out ? io_r_30_b : _GEN_3549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3551 = 8'h1f == r_count_17_io_out ? io_r_31_b : _GEN_3550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3552 = 8'h20 == r_count_17_io_out ? io_r_32_b : _GEN_3551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3553 = 8'h21 == r_count_17_io_out ? io_r_33_b : _GEN_3552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3554 = 8'h22 == r_count_17_io_out ? io_r_34_b : _GEN_3553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3555 = 8'h23 == r_count_17_io_out ? io_r_35_b : _GEN_3554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3556 = 8'h24 == r_count_17_io_out ? io_r_36_b : _GEN_3555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3557 = 8'h25 == r_count_17_io_out ? io_r_37_b : _GEN_3556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3558 = 8'h26 == r_count_17_io_out ? io_r_38_b : _GEN_3557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3559 = 8'h27 == r_count_17_io_out ? io_r_39_b : _GEN_3558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3560 = 8'h28 == r_count_17_io_out ? io_r_40_b : _GEN_3559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3561 = 8'h29 == r_count_17_io_out ? io_r_41_b : _GEN_3560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3562 = 8'h2a == r_count_17_io_out ? io_r_42_b : _GEN_3561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3563 = 8'h2b == r_count_17_io_out ? io_r_43_b : _GEN_3562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3564 = 8'h2c == r_count_17_io_out ? io_r_44_b : _GEN_3563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3565 = 8'h2d == r_count_17_io_out ? io_r_45_b : _GEN_3564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3566 = 8'h2e == r_count_17_io_out ? io_r_46_b : _GEN_3565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3567 = 8'h2f == r_count_17_io_out ? io_r_47_b : _GEN_3566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3568 = 8'h30 == r_count_17_io_out ? io_r_48_b : _GEN_3567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3569 = 8'h31 == r_count_17_io_out ? io_r_49_b : _GEN_3568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3570 = 8'h32 == r_count_17_io_out ? io_r_50_b : _GEN_3569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3571 = 8'h33 == r_count_17_io_out ? io_r_51_b : _GEN_3570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3572 = 8'h34 == r_count_17_io_out ? io_r_52_b : _GEN_3571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3573 = 8'h35 == r_count_17_io_out ? io_r_53_b : _GEN_3572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3574 = 8'h36 == r_count_17_io_out ? io_r_54_b : _GEN_3573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3575 = 8'h37 == r_count_17_io_out ? io_r_55_b : _GEN_3574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3576 = 8'h38 == r_count_17_io_out ? io_r_56_b : _GEN_3575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3577 = 8'h39 == r_count_17_io_out ? io_r_57_b : _GEN_3576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3578 = 8'h3a == r_count_17_io_out ? io_r_58_b : _GEN_3577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3579 = 8'h3b == r_count_17_io_out ? io_r_59_b : _GEN_3578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3580 = 8'h3c == r_count_17_io_out ? io_r_60_b : _GEN_3579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3581 = 8'h3d == r_count_17_io_out ? io_r_61_b : _GEN_3580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3582 = 8'h3e == r_count_17_io_out ? io_r_62_b : _GEN_3581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3583 = 8'h3f == r_count_17_io_out ? io_r_63_b : _GEN_3582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3584 = 8'h40 == r_count_17_io_out ? io_r_64_b : _GEN_3583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3585 = 8'h41 == r_count_17_io_out ? io_r_65_b : _GEN_3584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3586 = 8'h42 == r_count_17_io_out ? io_r_66_b : _GEN_3585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3587 = 8'h43 == r_count_17_io_out ? io_r_67_b : _GEN_3586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3588 = 8'h44 == r_count_17_io_out ? io_r_68_b : _GEN_3587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3589 = 8'h45 == r_count_17_io_out ? io_r_69_b : _GEN_3588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3590 = 8'h46 == r_count_17_io_out ? io_r_70_b : _GEN_3589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3591 = 8'h47 == r_count_17_io_out ? io_r_71_b : _GEN_3590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3592 = 8'h48 == r_count_17_io_out ? io_r_72_b : _GEN_3591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3593 = 8'h49 == r_count_17_io_out ? io_r_73_b : _GEN_3592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3594 = 8'h4a == r_count_17_io_out ? io_r_74_b : _GEN_3593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3595 = 8'h4b == r_count_17_io_out ? io_r_75_b : _GEN_3594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3596 = 8'h4c == r_count_17_io_out ? io_r_76_b : _GEN_3595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3597 = 8'h4d == r_count_17_io_out ? io_r_77_b : _GEN_3596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3598 = 8'h4e == r_count_17_io_out ? io_r_78_b : _GEN_3597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3599 = 8'h4f == r_count_17_io_out ? io_r_79_b : _GEN_3598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3600 = 8'h50 == r_count_17_io_out ? io_r_80_b : _GEN_3599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3601 = 8'h51 == r_count_17_io_out ? io_r_81_b : _GEN_3600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3602 = 8'h52 == r_count_17_io_out ? io_r_82_b : _GEN_3601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3603 = 8'h53 == r_count_17_io_out ? io_r_83_b : _GEN_3602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3604 = 8'h54 == r_count_17_io_out ? io_r_84_b : _GEN_3603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3605 = 8'h55 == r_count_17_io_out ? io_r_85_b : _GEN_3604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3606 = 8'h56 == r_count_17_io_out ? io_r_86_b : _GEN_3605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3607 = 8'h57 == r_count_17_io_out ? io_r_87_b : _GEN_3606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3608 = 8'h58 == r_count_17_io_out ? io_r_88_b : _GEN_3607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3609 = 8'h59 == r_count_17_io_out ? io_r_89_b : _GEN_3608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3610 = 8'h5a == r_count_17_io_out ? io_r_90_b : _GEN_3609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3611 = 8'h5b == r_count_17_io_out ? io_r_91_b : _GEN_3610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3612 = 8'h5c == r_count_17_io_out ? io_r_92_b : _GEN_3611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3613 = 8'h5d == r_count_17_io_out ? io_r_93_b : _GEN_3612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3614 = 8'h5e == r_count_17_io_out ? io_r_94_b : _GEN_3613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3615 = 8'h5f == r_count_17_io_out ? io_r_95_b : _GEN_3614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3616 = 8'h60 == r_count_17_io_out ? io_r_96_b : _GEN_3615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3617 = 8'h61 == r_count_17_io_out ? io_r_97_b : _GEN_3616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3618 = 8'h62 == r_count_17_io_out ? io_r_98_b : _GEN_3617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3619 = 8'h63 == r_count_17_io_out ? io_r_99_b : _GEN_3618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3620 = 8'h64 == r_count_17_io_out ? io_r_100_b : _GEN_3619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3621 = 8'h65 == r_count_17_io_out ? io_r_101_b : _GEN_3620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3622 = 8'h66 == r_count_17_io_out ? io_r_102_b : _GEN_3621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3623 = 8'h67 == r_count_17_io_out ? io_r_103_b : _GEN_3622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3624 = 8'h68 == r_count_17_io_out ? io_r_104_b : _GEN_3623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3625 = 8'h69 == r_count_17_io_out ? io_r_105_b : _GEN_3624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3626 = 8'h6a == r_count_17_io_out ? io_r_106_b : _GEN_3625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3627 = 8'h6b == r_count_17_io_out ? io_r_107_b : _GEN_3626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3628 = 8'h6c == r_count_17_io_out ? io_r_108_b : _GEN_3627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3629 = 8'h6d == r_count_17_io_out ? io_r_109_b : _GEN_3628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3630 = 8'h6e == r_count_17_io_out ? io_r_110_b : _GEN_3629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3631 = 8'h6f == r_count_17_io_out ? io_r_111_b : _GEN_3630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3632 = 8'h70 == r_count_17_io_out ? io_r_112_b : _GEN_3631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3633 = 8'h71 == r_count_17_io_out ? io_r_113_b : _GEN_3632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3634 = 8'h72 == r_count_17_io_out ? io_r_114_b : _GEN_3633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3635 = 8'h73 == r_count_17_io_out ? io_r_115_b : _GEN_3634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3636 = 8'h74 == r_count_17_io_out ? io_r_116_b : _GEN_3635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3637 = 8'h75 == r_count_17_io_out ? io_r_117_b : _GEN_3636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3638 = 8'h76 == r_count_17_io_out ? io_r_118_b : _GEN_3637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3639 = 8'h77 == r_count_17_io_out ? io_r_119_b : _GEN_3638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3640 = 8'h78 == r_count_17_io_out ? io_r_120_b : _GEN_3639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3641 = 8'h79 == r_count_17_io_out ? io_r_121_b : _GEN_3640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3642 = 8'h7a == r_count_17_io_out ? io_r_122_b : _GEN_3641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3643 = 8'h7b == r_count_17_io_out ? io_r_123_b : _GEN_3642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3644 = 8'h7c == r_count_17_io_out ? io_r_124_b : _GEN_3643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3645 = 8'h7d == r_count_17_io_out ? io_r_125_b : _GEN_3644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3646 = 8'h7e == r_count_17_io_out ? io_r_126_b : _GEN_3645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3647 = 8'h7f == r_count_17_io_out ? io_r_127_b : _GEN_3646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3648 = 8'h80 == r_count_17_io_out ? io_r_128_b : _GEN_3647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3649 = 8'h81 == r_count_17_io_out ? io_r_129_b : _GEN_3648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3650 = 8'h82 == r_count_17_io_out ? io_r_130_b : _GEN_3649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3651 = 8'h83 == r_count_17_io_out ? io_r_131_b : _GEN_3650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3652 = 8'h84 == r_count_17_io_out ? io_r_132_b : _GEN_3651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3653 = 8'h85 == r_count_17_io_out ? io_r_133_b : _GEN_3652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3654 = 8'h86 == r_count_17_io_out ? io_r_134_b : _GEN_3653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3655 = 8'h87 == r_count_17_io_out ? io_r_135_b : _GEN_3654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3656 = 8'h88 == r_count_17_io_out ? io_r_136_b : _GEN_3655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3657 = 8'h89 == r_count_17_io_out ? io_r_137_b : _GEN_3656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3658 = 8'h8a == r_count_17_io_out ? io_r_138_b : _GEN_3657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3659 = 8'h8b == r_count_17_io_out ? io_r_139_b : _GEN_3658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3660 = 8'h8c == r_count_17_io_out ? io_r_140_b : _GEN_3659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3661 = 8'h8d == r_count_17_io_out ? io_r_141_b : _GEN_3660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3662 = 8'h8e == r_count_17_io_out ? io_r_142_b : _GEN_3661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3663 = 8'h8f == r_count_17_io_out ? io_r_143_b : _GEN_3662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3664 = 8'h90 == r_count_17_io_out ? io_r_144_b : _GEN_3663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3665 = 8'h91 == r_count_17_io_out ? io_r_145_b : _GEN_3664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3666 = 8'h92 == r_count_17_io_out ? io_r_146_b : _GEN_3665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3667 = 8'h93 == r_count_17_io_out ? io_r_147_b : _GEN_3666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3668 = 8'h94 == r_count_17_io_out ? io_r_148_b : _GEN_3667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3669 = 8'h95 == r_count_17_io_out ? io_r_149_b : _GEN_3668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3670 = 8'h96 == r_count_17_io_out ? io_r_150_b : _GEN_3669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3671 = 8'h97 == r_count_17_io_out ? io_r_151_b : _GEN_3670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3672 = 8'h98 == r_count_17_io_out ? io_r_152_b : _GEN_3671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3673 = 8'h99 == r_count_17_io_out ? io_r_153_b : _GEN_3672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3674 = 8'h9a == r_count_17_io_out ? io_r_154_b : _GEN_3673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3675 = 8'h9b == r_count_17_io_out ? io_r_155_b : _GEN_3674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3676 = 8'h9c == r_count_17_io_out ? io_r_156_b : _GEN_3675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3677 = 8'h9d == r_count_17_io_out ? io_r_157_b : _GEN_3676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3678 = 8'h9e == r_count_17_io_out ? io_r_158_b : _GEN_3677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3679 = 8'h9f == r_count_17_io_out ? io_r_159_b : _GEN_3678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3680 = 8'ha0 == r_count_17_io_out ? io_r_160_b : _GEN_3679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3681 = 8'ha1 == r_count_17_io_out ? io_r_161_b : _GEN_3680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3682 = 8'ha2 == r_count_17_io_out ? io_r_162_b : _GEN_3681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3683 = 8'ha3 == r_count_17_io_out ? io_r_163_b : _GEN_3682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3684 = 8'ha4 == r_count_17_io_out ? io_r_164_b : _GEN_3683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3685 = 8'ha5 == r_count_17_io_out ? io_r_165_b : _GEN_3684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3686 = 8'ha6 == r_count_17_io_out ? io_r_166_b : _GEN_3685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3687 = 8'ha7 == r_count_17_io_out ? io_r_167_b : _GEN_3686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3688 = 8'ha8 == r_count_17_io_out ? io_r_168_b : _GEN_3687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3689 = 8'ha9 == r_count_17_io_out ? io_r_169_b : _GEN_3688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3690 = 8'haa == r_count_17_io_out ? io_r_170_b : _GEN_3689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3691 = 8'hab == r_count_17_io_out ? io_r_171_b : _GEN_3690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3692 = 8'hac == r_count_17_io_out ? io_r_172_b : _GEN_3691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3693 = 8'had == r_count_17_io_out ? io_r_173_b : _GEN_3692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3694 = 8'hae == r_count_17_io_out ? io_r_174_b : _GEN_3693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3695 = 8'haf == r_count_17_io_out ? io_r_175_b : _GEN_3694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3696 = 8'hb0 == r_count_17_io_out ? io_r_176_b : _GEN_3695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3697 = 8'hb1 == r_count_17_io_out ? io_r_177_b : _GEN_3696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3698 = 8'hb2 == r_count_17_io_out ? io_r_178_b : _GEN_3697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3699 = 8'hb3 == r_count_17_io_out ? io_r_179_b : _GEN_3698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3700 = 8'hb4 == r_count_17_io_out ? io_r_180_b : _GEN_3699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3701 = 8'hb5 == r_count_17_io_out ? io_r_181_b : _GEN_3700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3702 = 8'hb6 == r_count_17_io_out ? io_r_182_b : _GEN_3701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3703 = 8'hb7 == r_count_17_io_out ? io_r_183_b : _GEN_3702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3704 = 8'hb8 == r_count_17_io_out ? io_r_184_b : _GEN_3703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3705 = 8'hb9 == r_count_17_io_out ? io_r_185_b : _GEN_3704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3706 = 8'hba == r_count_17_io_out ? io_r_186_b : _GEN_3705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3707 = 8'hbb == r_count_17_io_out ? io_r_187_b : _GEN_3706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3708 = 8'hbc == r_count_17_io_out ? io_r_188_b : _GEN_3707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3709 = 8'hbd == r_count_17_io_out ? io_r_189_b : _GEN_3708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3710 = 8'hbe == r_count_17_io_out ? io_r_190_b : _GEN_3709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3711 = 8'hbf == r_count_17_io_out ? io_r_191_b : _GEN_3710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3712 = 8'hc0 == r_count_17_io_out ? io_r_192_b : _GEN_3711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3713 = 8'hc1 == r_count_17_io_out ? io_r_193_b : _GEN_3712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3714 = 8'hc2 == r_count_17_io_out ? io_r_194_b : _GEN_3713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3715 = 8'hc3 == r_count_17_io_out ? io_r_195_b : _GEN_3714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3716 = 8'hc4 == r_count_17_io_out ? io_r_196_b : _GEN_3715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3717 = 8'hc5 == r_count_17_io_out ? io_r_197_b : _GEN_3716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3718 = 8'hc6 == r_count_17_io_out ? io_r_198_b : _GEN_3717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3721 = 8'h1 == r_count_18_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3722 = 8'h2 == r_count_18_io_out ? io_r_2_b : _GEN_3721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3723 = 8'h3 == r_count_18_io_out ? io_r_3_b : _GEN_3722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3724 = 8'h4 == r_count_18_io_out ? io_r_4_b : _GEN_3723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3725 = 8'h5 == r_count_18_io_out ? io_r_5_b : _GEN_3724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3726 = 8'h6 == r_count_18_io_out ? io_r_6_b : _GEN_3725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3727 = 8'h7 == r_count_18_io_out ? io_r_7_b : _GEN_3726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3728 = 8'h8 == r_count_18_io_out ? io_r_8_b : _GEN_3727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3729 = 8'h9 == r_count_18_io_out ? io_r_9_b : _GEN_3728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3730 = 8'ha == r_count_18_io_out ? io_r_10_b : _GEN_3729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3731 = 8'hb == r_count_18_io_out ? io_r_11_b : _GEN_3730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3732 = 8'hc == r_count_18_io_out ? io_r_12_b : _GEN_3731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3733 = 8'hd == r_count_18_io_out ? io_r_13_b : _GEN_3732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3734 = 8'he == r_count_18_io_out ? io_r_14_b : _GEN_3733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3735 = 8'hf == r_count_18_io_out ? io_r_15_b : _GEN_3734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3736 = 8'h10 == r_count_18_io_out ? io_r_16_b : _GEN_3735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3737 = 8'h11 == r_count_18_io_out ? io_r_17_b : _GEN_3736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3738 = 8'h12 == r_count_18_io_out ? io_r_18_b : _GEN_3737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3739 = 8'h13 == r_count_18_io_out ? io_r_19_b : _GEN_3738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3740 = 8'h14 == r_count_18_io_out ? io_r_20_b : _GEN_3739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3741 = 8'h15 == r_count_18_io_out ? io_r_21_b : _GEN_3740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3742 = 8'h16 == r_count_18_io_out ? io_r_22_b : _GEN_3741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3743 = 8'h17 == r_count_18_io_out ? io_r_23_b : _GEN_3742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3744 = 8'h18 == r_count_18_io_out ? io_r_24_b : _GEN_3743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3745 = 8'h19 == r_count_18_io_out ? io_r_25_b : _GEN_3744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3746 = 8'h1a == r_count_18_io_out ? io_r_26_b : _GEN_3745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3747 = 8'h1b == r_count_18_io_out ? io_r_27_b : _GEN_3746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3748 = 8'h1c == r_count_18_io_out ? io_r_28_b : _GEN_3747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3749 = 8'h1d == r_count_18_io_out ? io_r_29_b : _GEN_3748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3750 = 8'h1e == r_count_18_io_out ? io_r_30_b : _GEN_3749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3751 = 8'h1f == r_count_18_io_out ? io_r_31_b : _GEN_3750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3752 = 8'h20 == r_count_18_io_out ? io_r_32_b : _GEN_3751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3753 = 8'h21 == r_count_18_io_out ? io_r_33_b : _GEN_3752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3754 = 8'h22 == r_count_18_io_out ? io_r_34_b : _GEN_3753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3755 = 8'h23 == r_count_18_io_out ? io_r_35_b : _GEN_3754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3756 = 8'h24 == r_count_18_io_out ? io_r_36_b : _GEN_3755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3757 = 8'h25 == r_count_18_io_out ? io_r_37_b : _GEN_3756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3758 = 8'h26 == r_count_18_io_out ? io_r_38_b : _GEN_3757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3759 = 8'h27 == r_count_18_io_out ? io_r_39_b : _GEN_3758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3760 = 8'h28 == r_count_18_io_out ? io_r_40_b : _GEN_3759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3761 = 8'h29 == r_count_18_io_out ? io_r_41_b : _GEN_3760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3762 = 8'h2a == r_count_18_io_out ? io_r_42_b : _GEN_3761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3763 = 8'h2b == r_count_18_io_out ? io_r_43_b : _GEN_3762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3764 = 8'h2c == r_count_18_io_out ? io_r_44_b : _GEN_3763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3765 = 8'h2d == r_count_18_io_out ? io_r_45_b : _GEN_3764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3766 = 8'h2e == r_count_18_io_out ? io_r_46_b : _GEN_3765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3767 = 8'h2f == r_count_18_io_out ? io_r_47_b : _GEN_3766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3768 = 8'h30 == r_count_18_io_out ? io_r_48_b : _GEN_3767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3769 = 8'h31 == r_count_18_io_out ? io_r_49_b : _GEN_3768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3770 = 8'h32 == r_count_18_io_out ? io_r_50_b : _GEN_3769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3771 = 8'h33 == r_count_18_io_out ? io_r_51_b : _GEN_3770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3772 = 8'h34 == r_count_18_io_out ? io_r_52_b : _GEN_3771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3773 = 8'h35 == r_count_18_io_out ? io_r_53_b : _GEN_3772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3774 = 8'h36 == r_count_18_io_out ? io_r_54_b : _GEN_3773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3775 = 8'h37 == r_count_18_io_out ? io_r_55_b : _GEN_3774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3776 = 8'h38 == r_count_18_io_out ? io_r_56_b : _GEN_3775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3777 = 8'h39 == r_count_18_io_out ? io_r_57_b : _GEN_3776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3778 = 8'h3a == r_count_18_io_out ? io_r_58_b : _GEN_3777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3779 = 8'h3b == r_count_18_io_out ? io_r_59_b : _GEN_3778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3780 = 8'h3c == r_count_18_io_out ? io_r_60_b : _GEN_3779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3781 = 8'h3d == r_count_18_io_out ? io_r_61_b : _GEN_3780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3782 = 8'h3e == r_count_18_io_out ? io_r_62_b : _GEN_3781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3783 = 8'h3f == r_count_18_io_out ? io_r_63_b : _GEN_3782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3784 = 8'h40 == r_count_18_io_out ? io_r_64_b : _GEN_3783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3785 = 8'h41 == r_count_18_io_out ? io_r_65_b : _GEN_3784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3786 = 8'h42 == r_count_18_io_out ? io_r_66_b : _GEN_3785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3787 = 8'h43 == r_count_18_io_out ? io_r_67_b : _GEN_3786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3788 = 8'h44 == r_count_18_io_out ? io_r_68_b : _GEN_3787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3789 = 8'h45 == r_count_18_io_out ? io_r_69_b : _GEN_3788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3790 = 8'h46 == r_count_18_io_out ? io_r_70_b : _GEN_3789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3791 = 8'h47 == r_count_18_io_out ? io_r_71_b : _GEN_3790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3792 = 8'h48 == r_count_18_io_out ? io_r_72_b : _GEN_3791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3793 = 8'h49 == r_count_18_io_out ? io_r_73_b : _GEN_3792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3794 = 8'h4a == r_count_18_io_out ? io_r_74_b : _GEN_3793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3795 = 8'h4b == r_count_18_io_out ? io_r_75_b : _GEN_3794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3796 = 8'h4c == r_count_18_io_out ? io_r_76_b : _GEN_3795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3797 = 8'h4d == r_count_18_io_out ? io_r_77_b : _GEN_3796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3798 = 8'h4e == r_count_18_io_out ? io_r_78_b : _GEN_3797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3799 = 8'h4f == r_count_18_io_out ? io_r_79_b : _GEN_3798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3800 = 8'h50 == r_count_18_io_out ? io_r_80_b : _GEN_3799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3801 = 8'h51 == r_count_18_io_out ? io_r_81_b : _GEN_3800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3802 = 8'h52 == r_count_18_io_out ? io_r_82_b : _GEN_3801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3803 = 8'h53 == r_count_18_io_out ? io_r_83_b : _GEN_3802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3804 = 8'h54 == r_count_18_io_out ? io_r_84_b : _GEN_3803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3805 = 8'h55 == r_count_18_io_out ? io_r_85_b : _GEN_3804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3806 = 8'h56 == r_count_18_io_out ? io_r_86_b : _GEN_3805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3807 = 8'h57 == r_count_18_io_out ? io_r_87_b : _GEN_3806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3808 = 8'h58 == r_count_18_io_out ? io_r_88_b : _GEN_3807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3809 = 8'h59 == r_count_18_io_out ? io_r_89_b : _GEN_3808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3810 = 8'h5a == r_count_18_io_out ? io_r_90_b : _GEN_3809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3811 = 8'h5b == r_count_18_io_out ? io_r_91_b : _GEN_3810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3812 = 8'h5c == r_count_18_io_out ? io_r_92_b : _GEN_3811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3813 = 8'h5d == r_count_18_io_out ? io_r_93_b : _GEN_3812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3814 = 8'h5e == r_count_18_io_out ? io_r_94_b : _GEN_3813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3815 = 8'h5f == r_count_18_io_out ? io_r_95_b : _GEN_3814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3816 = 8'h60 == r_count_18_io_out ? io_r_96_b : _GEN_3815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3817 = 8'h61 == r_count_18_io_out ? io_r_97_b : _GEN_3816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3818 = 8'h62 == r_count_18_io_out ? io_r_98_b : _GEN_3817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3819 = 8'h63 == r_count_18_io_out ? io_r_99_b : _GEN_3818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3820 = 8'h64 == r_count_18_io_out ? io_r_100_b : _GEN_3819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3821 = 8'h65 == r_count_18_io_out ? io_r_101_b : _GEN_3820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3822 = 8'h66 == r_count_18_io_out ? io_r_102_b : _GEN_3821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3823 = 8'h67 == r_count_18_io_out ? io_r_103_b : _GEN_3822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3824 = 8'h68 == r_count_18_io_out ? io_r_104_b : _GEN_3823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3825 = 8'h69 == r_count_18_io_out ? io_r_105_b : _GEN_3824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3826 = 8'h6a == r_count_18_io_out ? io_r_106_b : _GEN_3825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3827 = 8'h6b == r_count_18_io_out ? io_r_107_b : _GEN_3826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3828 = 8'h6c == r_count_18_io_out ? io_r_108_b : _GEN_3827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3829 = 8'h6d == r_count_18_io_out ? io_r_109_b : _GEN_3828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3830 = 8'h6e == r_count_18_io_out ? io_r_110_b : _GEN_3829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3831 = 8'h6f == r_count_18_io_out ? io_r_111_b : _GEN_3830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3832 = 8'h70 == r_count_18_io_out ? io_r_112_b : _GEN_3831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3833 = 8'h71 == r_count_18_io_out ? io_r_113_b : _GEN_3832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3834 = 8'h72 == r_count_18_io_out ? io_r_114_b : _GEN_3833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3835 = 8'h73 == r_count_18_io_out ? io_r_115_b : _GEN_3834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3836 = 8'h74 == r_count_18_io_out ? io_r_116_b : _GEN_3835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3837 = 8'h75 == r_count_18_io_out ? io_r_117_b : _GEN_3836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3838 = 8'h76 == r_count_18_io_out ? io_r_118_b : _GEN_3837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3839 = 8'h77 == r_count_18_io_out ? io_r_119_b : _GEN_3838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3840 = 8'h78 == r_count_18_io_out ? io_r_120_b : _GEN_3839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3841 = 8'h79 == r_count_18_io_out ? io_r_121_b : _GEN_3840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3842 = 8'h7a == r_count_18_io_out ? io_r_122_b : _GEN_3841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3843 = 8'h7b == r_count_18_io_out ? io_r_123_b : _GEN_3842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3844 = 8'h7c == r_count_18_io_out ? io_r_124_b : _GEN_3843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3845 = 8'h7d == r_count_18_io_out ? io_r_125_b : _GEN_3844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3846 = 8'h7e == r_count_18_io_out ? io_r_126_b : _GEN_3845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3847 = 8'h7f == r_count_18_io_out ? io_r_127_b : _GEN_3846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3848 = 8'h80 == r_count_18_io_out ? io_r_128_b : _GEN_3847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3849 = 8'h81 == r_count_18_io_out ? io_r_129_b : _GEN_3848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3850 = 8'h82 == r_count_18_io_out ? io_r_130_b : _GEN_3849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3851 = 8'h83 == r_count_18_io_out ? io_r_131_b : _GEN_3850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3852 = 8'h84 == r_count_18_io_out ? io_r_132_b : _GEN_3851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3853 = 8'h85 == r_count_18_io_out ? io_r_133_b : _GEN_3852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3854 = 8'h86 == r_count_18_io_out ? io_r_134_b : _GEN_3853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3855 = 8'h87 == r_count_18_io_out ? io_r_135_b : _GEN_3854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3856 = 8'h88 == r_count_18_io_out ? io_r_136_b : _GEN_3855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3857 = 8'h89 == r_count_18_io_out ? io_r_137_b : _GEN_3856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3858 = 8'h8a == r_count_18_io_out ? io_r_138_b : _GEN_3857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3859 = 8'h8b == r_count_18_io_out ? io_r_139_b : _GEN_3858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3860 = 8'h8c == r_count_18_io_out ? io_r_140_b : _GEN_3859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3861 = 8'h8d == r_count_18_io_out ? io_r_141_b : _GEN_3860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3862 = 8'h8e == r_count_18_io_out ? io_r_142_b : _GEN_3861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3863 = 8'h8f == r_count_18_io_out ? io_r_143_b : _GEN_3862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3864 = 8'h90 == r_count_18_io_out ? io_r_144_b : _GEN_3863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3865 = 8'h91 == r_count_18_io_out ? io_r_145_b : _GEN_3864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3866 = 8'h92 == r_count_18_io_out ? io_r_146_b : _GEN_3865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3867 = 8'h93 == r_count_18_io_out ? io_r_147_b : _GEN_3866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3868 = 8'h94 == r_count_18_io_out ? io_r_148_b : _GEN_3867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3869 = 8'h95 == r_count_18_io_out ? io_r_149_b : _GEN_3868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3870 = 8'h96 == r_count_18_io_out ? io_r_150_b : _GEN_3869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3871 = 8'h97 == r_count_18_io_out ? io_r_151_b : _GEN_3870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3872 = 8'h98 == r_count_18_io_out ? io_r_152_b : _GEN_3871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3873 = 8'h99 == r_count_18_io_out ? io_r_153_b : _GEN_3872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3874 = 8'h9a == r_count_18_io_out ? io_r_154_b : _GEN_3873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3875 = 8'h9b == r_count_18_io_out ? io_r_155_b : _GEN_3874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3876 = 8'h9c == r_count_18_io_out ? io_r_156_b : _GEN_3875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3877 = 8'h9d == r_count_18_io_out ? io_r_157_b : _GEN_3876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3878 = 8'h9e == r_count_18_io_out ? io_r_158_b : _GEN_3877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3879 = 8'h9f == r_count_18_io_out ? io_r_159_b : _GEN_3878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3880 = 8'ha0 == r_count_18_io_out ? io_r_160_b : _GEN_3879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3881 = 8'ha1 == r_count_18_io_out ? io_r_161_b : _GEN_3880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3882 = 8'ha2 == r_count_18_io_out ? io_r_162_b : _GEN_3881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3883 = 8'ha3 == r_count_18_io_out ? io_r_163_b : _GEN_3882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3884 = 8'ha4 == r_count_18_io_out ? io_r_164_b : _GEN_3883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3885 = 8'ha5 == r_count_18_io_out ? io_r_165_b : _GEN_3884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3886 = 8'ha6 == r_count_18_io_out ? io_r_166_b : _GEN_3885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3887 = 8'ha7 == r_count_18_io_out ? io_r_167_b : _GEN_3886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3888 = 8'ha8 == r_count_18_io_out ? io_r_168_b : _GEN_3887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3889 = 8'ha9 == r_count_18_io_out ? io_r_169_b : _GEN_3888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3890 = 8'haa == r_count_18_io_out ? io_r_170_b : _GEN_3889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3891 = 8'hab == r_count_18_io_out ? io_r_171_b : _GEN_3890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3892 = 8'hac == r_count_18_io_out ? io_r_172_b : _GEN_3891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3893 = 8'had == r_count_18_io_out ? io_r_173_b : _GEN_3892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3894 = 8'hae == r_count_18_io_out ? io_r_174_b : _GEN_3893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3895 = 8'haf == r_count_18_io_out ? io_r_175_b : _GEN_3894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3896 = 8'hb0 == r_count_18_io_out ? io_r_176_b : _GEN_3895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3897 = 8'hb1 == r_count_18_io_out ? io_r_177_b : _GEN_3896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3898 = 8'hb2 == r_count_18_io_out ? io_r_178_b : _GEN_3897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3899 = 8'hb3 == r_count_18_io_out ? io_r_179_b : _GEN_3898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3900 = 8'hb4 == r_count_18_io_out ? io_r_180_b : _GEN_3899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3901 = 8'hb5 == r_count_18_io_out ? io_r_181_b : _GEN_3900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3902 = 8'hb6 == r_count_18_io_out ? io_r_182_b : _GEN_3901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3903 = 8'hb7 == r_count_18_io_out ? io_r_183_b : _GEN_3902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3904 = 8'hb8 == r_count_18_io_out ? io_r_184_b : _GEN_3903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3905 = 8'hb9 == r_count_18_io_out ? io_r_185_b : _GEN_3904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3906 = 8'hba == r_count_18_io_out ? io_r_186_b : _GEN_3905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3907 = 8'hbb == r_count_18_io_out ? io_r_187_b : _GEN_3906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3908 = 8'hbc == r_count_18_io_out ? io_r_188_b : _GEN_3907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3909 = 8'hbd == r_count_18_io_out ? io_r_189_b : _GEN_3908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3910 = 8'hbe == r_count_18_io_out ? io_r_190_b : _GEN_3909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3911 = 8'hbf == r_count_18_io_out ? io_r_191_b : _GEN_3910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3912 = 8'hc0 == r_count_18_io_out ? io_r_192_b : _GEN_3911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3913 = 8'hc1 == r_count_18_io_out ? io_r_193_b : _GEN_3912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3914 = 8'hc2 == r_count_18_io_out ? io_r_194_b : _GEN_3913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3915 = 8'hc3 == r_count_18_io_out ? io_r_195_b : _GEN_3914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3916 = 8'hc4 == r_count_18_io_out ? io_r_196_b : _GEN_3915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3917 = 8'hc5 == r_count_18_io_out ? io_r_197_b : _GEN_3916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3918 = 8'hc6 == r_count_18_io_out ? io_r_198_b : _GEN_3917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3921 = 8'h1 == r_count_19_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3922 = 8'h2 == r_count_19_io_out ? io_r_2_b : _GEN_3921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3923 = 8'h3 == r_count_19_io_out ? io_r_3_b : _GEN_3922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3924 = 8'h4 == r_count_19_io_out ? io_r_4_b : _GEN_3923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3925 = 8'h5 == r_count_19_io_out ? io_r_5_b : _GEN_3924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3926 = 8'h6 == r_count_19_io_out ? io_r_6_b : _GEN_3925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3927 = 8'h7 == r_count_19_io_out ? io_r_7_b : _GEN_3926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3928 = 8'h8 == r_count_19_io_out ? io_r_8_b : _GEN_3927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3929 = 8'h9 == r_count_19_io_out ? io_r_9_b : _GEN_3928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3930 = 8'ha == r_count_19_io_out ? io_r_10_b : _GEN_3929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3931 = 8'hb == r_count_19_io_out ? io_r_11_b : _GEN_3930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3932 = 8'hc == r_count_19_io_out ? io_r_12_b : _GEN_3931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3933 = 8'hd == r_count_19_io_out ? io_r_13_b : _GEN_3932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3934 = 8'he == r_count_19_io_out ? io_r_14_b : _GEN_3933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3935 = 8'hf == r_count_19_io_out ? io_r_15_b : _GEN_3934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3936 = 8'h10 == r_count_19_io_out ? io_r_16_b : _GEN_3935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3937 = 8'h11 == r_count_19_io_out ? io_r_17_b : _GEN_3936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3938 = 8'h12 == r_count_19_io_out ? io_r_18_b : _GEN_3937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3939 = 8'h13 == r_count_19_io_out ? io_r_19_b : _GEN_3938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3940 = 8'h14 == r_count_19_io_out ? io_r_20_b : _GEN_3939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3941 = 8'h15 == r_count_19_io_out ? io_r_21_b : _GEN_3940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3942 = 8'h16 == r_count_19_io_out ? io_r_22_b : _GEN_3941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3943 = 8'h17 == r_count_19_io_out ? io_r_23_b : _GEN_3942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3944 = 8'h18 == r_count_19_io_out ? io_r_24_b : _GEN_3943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3945 = 8'h19 == r_count_19_io_out ? io_r_25_b : _GEN_3944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3946 = 8'h1a == r_count_19_io_out ? io_r_26_b : _GEN_3945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3947 = 8'h1b == r_count_19_io_out ? io_r_27_b : _GEN_3946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3948 = 8'h1c == r_count_19_io_out ? io_r_28_b : _GEN_3947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3949 = 8'h1d == r_count_19_io_out ? io_r_29_b : _GEN_3948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3950 = 8'h1e == r_count_19_io_out ? io_r_30_b : _GEN_3949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3951 = 8'h1f == r_count_19_io_out ? io_r_31_b : _GEN_3950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3952 = 8'h20 == r_count_19_io_out ? io_r_32_b : _GEN_3951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3953 = 8'h21 == r_count_19_io_out ? io_r_33_b : _GEN_3952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3954 = 8'h22 == r_count_19_io_out ? io_r_34_b : _GEN_3953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3955 = 8'h23 == r_count_19_io_out ? io_r_35_b : _GEN_3954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3956 = 8'h24 == r_count_19_io_out ? io_r_36_b : _GEN_3955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3957 = 8'h25 == r_count_19_io_out ? io_r_37_b : _GEN_3956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3958 = 8'h26 == r_count_19_io_out ? io_r_38_b : _GEN_3957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3959 = 8'h27 == r_count_19_io_out ? io_r_39_b : _GEN_3958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3960 = 8'h28 == r_count_19_io_out ? io_r_40_b : _GEN_3959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3961 = 8'h29 == r_count_19_io_out ? io_r_41_b : _GEN_3960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3962 = 8'h2a == r_count_19_io_out ? io_r_42_b : _GEN_3961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3963 = 8'h2b == r_count_19_io_out ? io_r_43_b : _GEN_3962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3964 = 8'h2c == r_count_19_io_out ? io_r_44_b : _GEN_3963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3965 = 8'h2d == r_count_19_io_out ? io_r_45_b : _GEN_3964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3966 = 8'h2e == r_count_19_io_out ? io_r_46_b : _GEN_3965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3967 = 8'h2f == r_count_19_io_out ? io_r_47_b : _GEN_3966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3968 = 8'h30 == r_count_19_io_out ? io_r_48_b : _GEN_3967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3969 = 8'h31 == r_count_19_io_out ? io_r_49_b : _GEN_3968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3970 = 8'h32 == r_count_19_io_out ? io_r_50_b : _GEN_3969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3971 = 8'h33 == r_count_19_io_out ? io_r_51_b : _GEN_3970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3972 = 8'h34 == r_count_19_io_out ? io_r_52_b : _GEN_3971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3973 = 8'h35 == r_count_19_io_out ? io_r_53_b : _GEN_3972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3974 = 8'h36 == r_count_19_io_out ? io_r_54_b : _GEN_3973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3975 = 8'h37 == r_count_19_io_out ? io_r_55_b : _GEN_3974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3976 = 8'h38 == r_count_19_io_out ? io_r_56_b : _GEN_3975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3977 = 8'h39 == r_count_19_io_out ? io_r_57_b : _GEN_3976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3978 = 8'h3a == r_count_19_io_out ? io_r_58_b : _GEN_3977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3979 = 8'h3b == r_count_19_io_out ? io_r_59_b : _GEN_3978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3980 = 8'h3c == r_count_19_io_out ? io_r_60_b : _GEN_3979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3981 = 8'h3d == r_count_19_io_out ? io_r_61_b : _GEN_3980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3982 = 8'h3e == r_count_19_io_out ? io_r_62_b : _GEN_3981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3983 = 8'h3f == r_count_19_io_out ? io_r_63_b : _GEN_3982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3984 = 8'h40 == r_count_19_io_out ? io_r_64_b : _GEN_3983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3985 = 8'h41 == r_count_19_io_out ? io_r_65_b : _GEN_3984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3986 = 8'h42 == r_count_19_io_out ? io_r_66_b : _GEN_3985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3987 = 8'h43 == r_count_19_io_out ? io_r_67_b : _GEN_3986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3988 = 8'h44 == r_count_19_io_out ? io_r_68_b : _GEN_3987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3989 = 8'h45 == r_count_19_io_out ? io_r_69_b : _GEN_3988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3990 = 8'h46 == r_count_19_io_out ? io_r_70_b : _GEN_3989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3991 = 8'h47 == r_count_19_io_out ? io_r_71_b : _GEN_3990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3992 = 8'h48 == r_count_19_io_out ? io_r_72_b : _GEN_3991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3993 = 8'h49 == r_count_19_io_out ? io_r_73_b : _GEN_3992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3994 = 8'h4a == r_count_19_io_out ? io_r_74_b : _GEN_3993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3995 = 8'h4b == r_count_19_io_out ? io_r_75_b : _GEN_3994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3996 = 8'h4c == r_count_19_io_out ? io_r_76_b : _GEN_3995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3997 = 8'h4d == r_count_19_io_out ? io_r_77_b : _GEN_3996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3998 = 8'h4e == r_count_19_io_out ? io_r_78_b : _GEN_3997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3999 = 8'h4f == r_count_19_io_out ? io_r_79_b : _GEN_3998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4000 = 8'h50 == r_count_19_io_out ? io_r_80_b : _GEN_3999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4001 = 8'h51 == r_count_19_io_out ? io_r_81_b : _GEN_4000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4002 = 8'h52 == r_count_19_io_out ? io_r_82_b : _GEN_4001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4003 = 8'h53 == r_count_19_io_out ? io_r_83_b : _GEN_4002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4004 = 8'h54 == r_count_19_io_out ? io_r_84_b : _GEN_4003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4005 = 8'h55 == r_count_19_io_out ? io_r_85_b : _GEN_4004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4006 = 8'h56 == r_count_19_io_out ? io_r_86_b : _GEN_4005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4007 = 8'h57 == r_count_19_io_out ? io_r_87_b : _GEN_4006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4008 = 8'h58 == r_count_19_io_out ? io_r_88_b : _GEN_4007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4009 = 8'h59 == r_count_19_io_out ? io_r_89_b : _GEN_4008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4010 = 8'h5a == r_count_19_io_out ? io_r_90_b : _GEN_4009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4011 = 8'h5b == r_count_19_io_out ? io_r_91_b : _GEN_4010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4012 = 8'h5c == r_count_19_io_out ? io_r_92_b : _GEN_4011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4013 = 8'h5d == r_count_19_io_out ? io_r_93_b : _GEN_4012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4014 = 8'h5e == r_count_19_io_out ? io_r_94_b : _GEN_4013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4015 = 8'h5f == r_count_19_io_out ? io_r_95_b : _GEN_4014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4016 = 8'h60 == r_count_19_io_out ? io_r_96_b : _GEN_4015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4017 = 8'h61 == r_count_19_io_out ? io_r_97_b : _GEN_4016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4018 = 8'h62 == r_count_19_io_out ? io_r_98_b : _GEN_4017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4019 = 8'h63 == r_count_19_io_out ? io_r_99_b : _GEN_4018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4020 = 8'h64 == r_count_19_io_out ? io_r_100_b : _GEN_4019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4021 = 8'h65 == r_count_19_io_out ? io_r_101_b : _GEN_4020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4022 = 8'h66 == r_count_19_io_out ? io_r_102_b : _GEN_4021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4023 = 8'h67 == r_count_19_io_out ? io_r_103_b : _GEN_4022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4024 = 8'h68 == r_count_19_io_out ? io_r_104_b : _GEN_4023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4025 = 8'h69 == r_count_19_io_out ? io_r_105_b : _GEN_4024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4026 = 8'h6a == r_count_19_io_out ? io_r_106_b : _GEN_4025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4027 = 8'h6b == r_count_19_io_out ? io_r_107_b : _GEN_4026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4028 = 8'h6c == r_count_19_io_out ? io_r_108_b : _GEN_4027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4029 = 8'h6d == r_count_19_io_out ? io_r_109_b : _GEN_4028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4030 = 8'h6e == r_count_19_io_out ? io_r_110_b : _GEN_4029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4031 = 8'h6f == r_count_19_io_out ? io_r_111_b : _GEN_4030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4032 = 8'h70 == r_count_19_io_out ? io_r_112_b : _GEN_4031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4033 = 8'h71 == r_count_19_io_out ? io_r_113_b : _GEN_4032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4034 = 8'h72 == r_count_19_io_out ? io_r_114_b : _GEN_4033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4035 = 8'h73 == r_count_19_io_out ? io_r_115_b : _GEN_4034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4036 = 8'h74 == r_count_19_io_out ? io_r_116_b : _GEN_4035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4037 = 8'h75 == r_count_19_io_out ? io_r_117_b : _GEN_4036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4038 = 8'h76 == r_count_19_io_out ? io_r_118_b : _GEN_4037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4039 = 8'h77 == r_count_19_io_out ? io_r_119_b : _GEN_4038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4040 = 8'h78 == r_count_19_io_out ? io_r_120_b : _GEN_4039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4041 = 8'h79 == r_count_19_io_out ? io_r_121_b : _GEN_4040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4042 = 8'h7a == r_count_19_io_out ? io_r_122_b : _GEN_4041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4043 = 8'h7b == r_count_19_io_out ? io_r_123_b : _GEN_4042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4044 = 8'h7c == r_count_19_io_out ? io_r_124_b : _GEN_4043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4045 = 8'h7d == r_count_19_io_out ? io_r_125_b : _GEN_4044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4046 = 8'h7e == r_count_19_io_out ? io_r_126_b : _GEN_4045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4047 = 8'h7f == r_count_19_io_out ? io_r_127_b : _GEN_4046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4048 = 8'h80 == r_count_19_io_out ? io_r_128_b : _GEN_4047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4049 = 8'h81 == r_count_19_io_out ? io_r_129_b : _GEN_4048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4050 = 8'h82 == r_count_19_io_out ? io_r_130_b : _GEN_4049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4051 = 8'h83 == r_count_19_io_out ? io_r_131_b : _GEN_4050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4052 = 8'h84 == r_count_19_io_out ? io_r_132_b : _GEN_4051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4053 = 8'h85 == r_count_19_io_out ? io_r_133_b : _GEN_4052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4054 = 8'h86 == r_count_19_io_out ? io_r_134_b : _GEN_4053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4055 = 8'h87 == r_count_19_io_out ? io_r_135_b : _GEN_4054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4056 = 8'h88 == r_count_19_io_out ? io_r_136_b : _GEN_4055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4057 = 8'h89 == r_count_19_io_out ? io_r_137_b : _GEN_4056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4058 = 8'h8a == r_count_19_io_out ? io_r_138_b : _GEN_4057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4059 = 8'h8b == r_count_19_io_out ? io_r_139_b : _GEN_4058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4060 = 8'h8c == r_count_19_io_out ? io_r_140_b : _GEN_4059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4061 = 8'h8d == r_count_19_io_out ? io_r_141_b : _GEN_4060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4062 = 8'h8e == r_count_19_io_out ? io_r_142_b : _GEN_4061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4063 = 8'h8f == r_count_19_io_out ? io_r_143_b : _GEN_4062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4064 = 8'h90 == r_count_19_io_out ? io_r_144_b : _GEN_4063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4065 = 8'h91 == r_count_19_io_out ? io_r_145_b : _GEN_4064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4066 = 8'h92 == r_count_19_io_out ? io_r_146_b : _GEN_4065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4067 = 8'h93 == r_count_19_io_out ? io_r_147_b : _GEN_4066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4068 = 8'h94 == r_count_19_io_out ? io_r_148_b : _GEN_4067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4069 = 8'h95 == r_count_19_io_out ? io_r_149_b : _GEN_4068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4070 = 8'h96 == r_count_19_io_out ? io_r_150_b : _GEN_4069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4071 = 8'h97 == r_count_19_io_out ? io_r_151_b : _GEN_4070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4072 = 8'h98 == r_count_19_io_out ? io_r_152_b : _GEN_4071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4073 = 8'h99 == r_count_19_io_out ? io_r_153_b : _GEN_4072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4074 = 8'h9a == r_count_19_io_out ? io_r_154_b : _GEN_4073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4075 = 8'h9b == r_count_19_io_out ? io_r_155_b : _GEN_4074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4076 = 8'h9c == r_count_19_io_out ? io_r_156_b : _GEN_4075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4077 = 8'h9d == r_count_19_io_out ? io_r_157_b : _GEN_4076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4078 = 8'h9e == r_count_19_io_out ? io_r_158_b : _GEN_4077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4079 = 8'h9f == r_count_19_io_out ? io_r_159_b : _GEN_4078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4080 = 8'ha0 == r_count_19_io_out ? io_r_160_b : _GEN_4079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4081 = 8'ha1 == r_count_19_io_out ? io_r_161_b : _GEN_4080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4082 = 8'ha2 == r_count_19_io_out ? io_r_162_b : _GEN_4081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4083 = 8'ha3 == r_count_19_io_out ? io_r_163_b : _GEN_4082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4084 = 8'ha4 == r_count_19_io_out ? io_r_164_b : _GEN_4083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4085 = 8'ha5 == r_count_19_io_out ? io_r_165_b : _GEN_4084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4086 = 8'ha6 == r_count_19_io_out ? io_r_166_b : _GEN_4085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4087 = 8'ha7 == r_count_19_io_out ? io_r_167_b : _GEN_4086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4088 = 8'ha8 == r_count_19_io_out ? io_r_168_b : _GEN_4087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4089 = 8'ha9 == r_count_19_io_out ? io_r_169_b : _GEN_4088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4090 = 8'haa == r_count_19_io_out ? io_r_170_b : _GEN_4089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4091 = 8'hab == r_count_19_io_out ? io_r_171_b : _GEN_4090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4092 = 8'hac == r_count_19_io_out ? io_r_172_b : _GEN_4091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4093 = 8'had == r_count_19_io_out ? io_r_173_b : _GEN_4092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4094 = 8'hae == r_count_19_io_out ? io_r_174_b : _GEN_4093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4095 = 8'haf == r_count_19_io_out ? io_r_175_b : _GEN_4094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4096 = 8'hb0 == r_count_19_io_out ? io_r_176_b : _GEN_4095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4097 = 8'hb1 == r_count_19_io_out ? io_r_177_b : _GEN_4096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4098 = 8'hb2 == r_count_19_io_out ? io_r_178_b : _GEN_4097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4099 = 8'hb3 == r_count_19_io_out ? io_r_179_b : _GEN_4098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4100 = 8'hb4 == r_count_19_io_out ? io_r_180_b : _GEN_4099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4101 = 8'hb5 == r_count_19_io_out ? io_r_181_b : _GEN_4100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4102 = 8'hb6 == r_count_19_io_out ? io_r_182_b : _GEN_4101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4103 = 8'hb7 == r_count_19_io_out ? io_r_183_b : _GEN_4102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4104 = 8'hb8 == r_count_19_io_out ? io_r_184_b : _GEN_4103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4105 = 8'hb9 == r_count_19_io_out ? io_r_185_b : _GEN_4104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4106 = 8'hba == r_count_19_io_out ? io_r_186_b : _GEN_4105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4107 = 8'hbb == r_count_19_io_out ? io_r_187_b : _GEN_4106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4108 = 8'hbc == r_count_19_io_out ? io_r_188_b : _GEN_4107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4109 = 8'hbd == r_count_19_io_out ? io_r_189_b : _GEN_4108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4110 = 8'hbe == r_count_19_io_out ? io_r_190_b : _GEN_4109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4111 = 8'hbf == r_count_19_io_out ? io_r_191_b : _GEN_4110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4112 = 8'hc0 == r_count_19_io_out ? io_r_192_b : _GEN_4111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4113 = 8'hc1 == r_count_19_io_out ? io_r_193_b : _GEN_4112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4114 = 8'hc2 == r_count_19_io_out ? io_r_194_b : _GEN_4113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4115 = 8'hc3 == r_count_19_io_out ? io_r_195_b : _GEN_4114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4116 = 8'hc4 == r_count_19_io_out ? io_r_196_b : _GEN_4115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4117 = 8'hc5 == r_count_19_io_out ? io_r_197_b : _GEN_4116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4118 = 8'hc6 == r_count_19_io_out ? io_r_198_b : _GEN_4117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4121 = 8'h1 == r_count_20_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4122 = 8'h2 == r_count_20_io_out ? io_r_2_b : _GEN_4121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4123 = 8'h3 == r_count_20_io_out ? io_r_3_b : _GEN_4122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4124 = 8'h4 == r_count_20_io_out ? io_r_4_b : _GEN_4123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4125 = 8'h5 == r_count_20_io_out ? io_r_5_b : _GEN_4124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4126 = 8'h6 == r_count_20_io_out ? io_r_6_b : _GEN_4125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4127 = 8'h7 == r_count_20_io_out ? io_r_7_b : _GEN_4126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4128 = 8'h8 == r_count_20_io_out ? io_r_8_b : _GEN_4127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4129 = 8'h9 == r_count_20_io_out ? io_r_9_b : _GEN_4128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4130 = 8'ha == r_count_20_io_out ? io_r_10_b : _GEN_4129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4131 = 8'hb == r_count_20_io_out ? io_r_11_b : _GEN_4130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4132 = 8'hc == r_count_20_io_out ? io_r_12_b : _GEN_4131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4133 = 8'hd == r_count_20_io_out ? io_r_13_b : _GEN_4132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4134 = 8'he == r_count_20_io_out ? io_r_14_b : _GEN_4133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4135 = 8'hf == r_count_20_io_out ? io_r_15_b : _GEN_4134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4136 = 8'h10 == r_count_20_io_out ? io_r_16_b : _GEN_4135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4137 = 8'h11 == r_count_20_io_out ? io_r_17_b : _GEN_4136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4138 = 8'h12 == r_count_20_io_out ? io_r_18_b : _GEN_4137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4139 = 8'h13 == r_count_20_io_out ? io_r_19_b : _GEN_4138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4140 = 8'h14 == r_count_20_io_out ? io_r_20_b : _GEN_4139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4141 = 8'h15 == r_count_20_io_out ? io_r_21_b : _GEN_4140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4142 = 8'h16 == r_count_20_io_out ? io_r_22_b : _GEN_4141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4143 = 8'h17 == r_count_20_io_out ? io_r_23_b : _GEN_4142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4144 = 8'h18 == r_count_20_io_out ? io_r_24_b : _GEN_4143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4145 = 8'h19 == r_count_20_io_out ? io_r_25_b : _GEN_4144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4146 = 8'h1a == r_count_20_io_out ? io_r_26_b : _GEN_4145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4147 = 8'h1b == r_count_20_io_out ? io_r_27_b : _GEN_4146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4148 = 8'h1c == r_count_20_io_out ? io_r_28_b : _GEN_4147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4149 = 8'h1d == r_count_20_io_out ? io_r_29_b : _GEN_4148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4150 = 8'h1e == r_count_20_io_out ? io_r_30_b : _GEN_4149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4151 = 8'h1f == r_count_20_io_out ? io_r_31_b : _GEN_4150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4152 = 8'h20 == r_count_20_io_out ? io_r_32_b : _GEN_4151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4153 = 8'h21 == r_count_20_io_out ? io_r_33_b : _GEN_4152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4154 = 8'h22 == r_count_20_io_out ? io_r_34_b : _GEN_4153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4155 = 8'h23 == r_count_20_io_out ? io_r_35_b : _GEN_4154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4156 = 8'h24 == r_count_20_io_out ? io_r_36_b : _GEN_4155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4157 = 8'h25 == r_count_20_io_out ? io_r_37_b : _GEN_4156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4158 = 8'h26 == r_count_20_io_out ? io_r_38_b : _GEN_4157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4159 = 8'h27 == r_count_20_io_out ? io_r_39_b : _GEN_4158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4160 = 8'h28 == r_count_20_io_out ? io_r_40_b : _GEN_4159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4161 = 8'h29 == r_count_20_io_out ? io_r_41_b : _GEN_4160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4162 = 8'h2a == r_count_20_io_out ? io_r_42_b : _GEN_4161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4163 = 8'h2b == r_count_20_io_out ? io_r_43_b : _GEN_4162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4164 = 8'h2c == r_count_20_io_out ? io_r_44_b : _GEN_4163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4165 = 8'h2d == r_count_20_io_out ? io_r_45_b : _GEN_4164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4166 = 8'h2e == r_count_20_io_out ? io_r_46_b : _GEN_4165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4167 = 8'h2f == r_count_20_io_out ? io_r_47_b : _GEN_4166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4168 = 8'h30 == r_count_20_io_out ? io_r_48_b : _GEN_4167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4169 = 8'h31 == r_count_20_io_out ? io_r_49_b : _GEN_4168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4170 = 8'h32 == r_count_20_io_out ? io_r_50_b : _GEN_4169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4171 = 8'h33 == r_count_20_io_out ? io_r_51_b : _GEN_4170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4172 = 8'h34 == r_count_20_io_out ? io_r_52_b : _GEN_4171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4173 = 8'h35 == r_count_20_io_out ? io_r_53_b : _GEN_4172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4174 = 8'h36 == r_count_20_io_out ? io_r_54_b : _GEN_4173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4175 = 8'h37 == r_count_20_io_out ? io_r_55_b : _GEN_4174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4176 = 8'h38 == r_count_20_io_out ? io_r_56_b : _GEN_4175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4177 = 8'h39 == r_count_20_io_out ? io_r_57_b : _GEN_4176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4178 = 8'h3a == r_count_20_io_out ? io_r_58_b : _GEN_4177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4179 = 8'h3b == r_count_20_io_out ? io_r_59_b : _GEN_4178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4180 = 8'h3c == r_count_20_io_out ? io_r_60_b : _GEN_4179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4181 = 8'h3d == r_count_20_io_out ? io_r_61_b : _GEN_4180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4182 = 8'h3e == r_count_20_io_out ? io_r_62_b : _GEN_4181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4183 = 8'h3f == r_count_20_io_out ? io_r_63_b : _GEN_4182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4184 = 8'h40 == r_count_20_io_out ? io_r_64_b : _GEN_4183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4185 = 8'h41 == r_count_20_io_out ? io_r_65_b : _GEN_4184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4186 = 8'h42 == r_count_20_io_out ? io_r_66_b : _GEN_4185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4187 = 8'h43 == r_count_20_io_out ? io_r_67_b : _GEN_4186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4188 = 8'h44 == r_count_20_io_out ? io_r_68_b : _GEN_4187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4189 = 8'h45 == r_count_20_io_out ? io_r_69_b : _GEN_4188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4190 = 8'h46 == r_count_20_io_out ? io_r_70_b : _GEN_4189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4191 = 8'h47 == r_count_20_io_out ? io_r_71_b : _GEN_4190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4192 = 8'h48 == r_count_20_io_out ? io_r_72_b : _GEN_4191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4193 = 8'h49 == r_count_20_io_out ? io_r_73_b : _GEN_4192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4194 = 8'h4a == r_count_20_io_out ? io_r_74_b : _GEN_4193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4195 = 8'h4b == r_count_20_io_out ? io_r_75_b : _GEN_4194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4196 = 8'h4c == r_count_20_io_out ? io_r_76_b : _GEN_4195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4197 = 8'h4d == r_count_20_io_out ? io_r_77_b : _GEN_4196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4198 = 8'h4e == r_count_20_io_out ? io_r_78_b : _GEN_4197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4199 = 8'h4f == r_count_20_io_out ? io_r_79_b : _GEN_4198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4200 = 8'h50 == r_count_20_io_out ? io_r_80_b : _GEN_4199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4201 = 8'h51 == r_count_20_io_out ? io_r_81_b : _GEN_4200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4202 = 8'h52 == r_count_20_io_out ? io_r_82_b : _GEN_4201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4203 = 8'h53 == r_count_20_io_out ? io_r_83_b : _GEN_4202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4204 = 8'h54 == r_count_20_io_out ? io_r_84_b : _GEN_4203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4205 = 8'h55 == r_count_20_io_out ? io_r_85_b : _GEN_4204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4206 = 8'h56 == r_count_20_io_out ? io_r_86_b : _GEN_4205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4207 = 8'h57 == r_count_20_io_out ? io_r_87_b : _GEN_4206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4208 = 8'h58 == r_count_20_io_out ? io_r_88_b : _GEN_4207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4209 = 8'h59 == r_count_20_io_out ? io_r_89_b : _GEN_4208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4210 = 8'h5a == r_count_20_io_out ? io_r_90_b : _GEN_4209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4211 = 8'h5b == r_count_20_io_out ? io_r_91_b : _GEN_4210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4212 = 8'h5c == r_count_20_io_out ? io_r_92_b : _GEN_4211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4213 = 8'h5d == r_count_20_io_out ? io_r_93_b : _GEN_4212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4214 = 8'h5e == r_count_20_io_out ? io_r_94_b : _GEN_4213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4215 = 8'h5f == r_count_20_io_out ? io_r_95_b : _GEN_4214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4216 = 8'h60 == r_count_20_io_out ? io_r_96_b : _GEN_4215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4217 = 8'h61 == r_count_20_io_out ? io_r_97_b : _GEN_4216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4218 = 8'h62 == r_count_20_io_out ? io_r_98_b : _GEN_4217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4219 = 8'h63 == r_count_20_io_out ? io_r_99_b : _GEN_4218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4220 = 8'h64 == r_count_20_io_out ? io_r_100_b : _GEN_4219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4221 = 8'h65 == r_count_20_io_out ? io_r_101_b : _GEN_4220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4222 = 8'h66 == r_count_20_io_out ? io_r_102_b : _GEN_4221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4223 = 8'h67 == r_count_20_io_out ? io_r_103_b : _GEN_4222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4224 = 8'h68 == r_count_20_io_out ? io_r_104_b : _GEN_4223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4225 = 8'h69 == r_count_20_io_out ? io_r_105_b : _GEN_4224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4226 = 8'h6a == r_count_20_io_out ? io_r_106_b : _GEN_4225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4227 = 8'h6b == r_count_20_io_out ? io_r_107_b : _GEN_4226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4228 = 8'h6c == r_count_20_io_out ? io_r_108_b : _GEN_4227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4229 = 8'h6d == r_count_20_io_out ? io_r_109_b : _GEN_4228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4230 = 8'h6e == r_count_20_io_out ? io_r_110_b : _GEN_4229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4231 = 8'h6f == r_count_20_io_out ? io_r_111_b : _GEN_4230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4232 = 8'h70 == r_count_20_io_out ? io_r_112_b : _GEN_4231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4233 = 8'h71 == r_count_20_io_out ? io_r_113_b : _GEN_4232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4234 = 8'h72 == r_count_20_io_out ? io_r_114_b : _GEN_4233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4235 = 8'h73 == r_count_20_io_out ? io_r_115_b : _GEN_4234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4236 = 8'h74 == r_count_20_io_out ? io_r_116_b : _GEN_4235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4237 = 8'h75 == r_count_20_io_out ? io_r_117_b : _GEN_4236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4238 = 8'h76 == r_count_20_io_out ? io_r_118_b : _GEN_4237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4239 = 8'h77 == r_count_20_io_out ? io_r_119_b : _GEN_4238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4240 = 8'h78 == r_count_20_io_out ? io_r_120_b : _GEN_4239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4241 = 8'h79 == r_count_20_io_out ? io_r_121_b : _GEN_4240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4242 = 8'h7a == r_count_20_io_out ? io_r_122_b : _GEN_4241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4243 = 8'h7b == r_count_20_io_out ? io_r_123_b : _GEN_4242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4244 = 8'h7c == r_count_20_io_out ? io_r_124_b : _GEN_4243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4245 = 8'h7d == r_count_20_io_out ? io_r_125_b : _GEN_4244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4246 = 8'h7e == r_count_20_io_out ? io_r_126_b : _GEN_4245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4247 = 8'h7f == r_count_20_io_out ? io_r_127_b : _GEN_4246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4248 = 8'h80 == r_count_20_io_out ? io_r_128_b : _GEN_4247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4249 = 8'h81 == r_count_20_io_out ? io_r_129_b : _GEN_4248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4250 = 8'h82 == r_count_20_io_out ? io_r_130_b : _GEN_4249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4251 = 8'h83 == r_count_20_io_out ? io_r_131_b : _GEN_4250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4252 = 8'h84 == r_count_20_io_out ? io_r_132_b : _GEN_4251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4253 = 8'h85 == r_count_20_io_out ? io_r_133_b : _GEN_4252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4254 = 8'h86 == r_count_20_io_out ? io_r_134_b : _GEN_4253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4255 = 8'h87 == r_count_20_io_out ? io_r_135_b : _GEN_4254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4256 = 8'h88 == r_count_20_io_out ? io_r_136_b : _GEN_4255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4257 = 8'h89 == r_count_20_io_out ? io_r_137_b : _GEN_4256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4258 = 8'h8a == r_count_20_io_out ? io_r_138_b : _GEN_4257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4259 = 8'h8b == r_count_20_io_out ? io_r_139_b : _GEN_4258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4260 = 8'h8c == r_count_20_io_out ? io_r_140_b : _GEN_4259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4261 = 8'h8d == r_count_20_io_out ? io_r_141_b : _GEN_4260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4262 = 8'h8e == r_count_20_io_out ? io_r_142_b : _GEN_4261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4263 = 8'h8f == r_count_20_io_out ? io_r_143_b : _GEN_4262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4264 = 8'h90 == r_count_20_io_out ? io_r_144_b : _GEN_4263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4265 = 8'h91 == r_count_20_io_out ? io_r_145_b : _GEN_4264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4266 = 8'h92 == r_count_20_io_out ? io_r_146_b : _GEN_4265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4267 = 8'h93 == r_count_20_io_out ? io_r_147_b : _GEN_4266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4268 = 8'h94 == r_count_20_io_out ? io_r_148_b : _GEN_4267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4269 = 8'h95 == r_count_20_io_out ? io_r_149_b : _GEN_4268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4270 = 8'h96 == r_count_20_io_out ? io_r_150_b : _GEN_4269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4271 = 8'h97 == r_count_20_io_out ? io_r_151_b : _GEN_4270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4272 = 8'h98 == r_count_20_io_out ? io_r_152_b : _GEN_4271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4273 = 8'h99 == r_count_20_io_out ? io_r_153_b : _GEN_4272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4274 = 8'h9a == r_count_20_io_out ? io_r_154_b : _GEN_4273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4275 = 8'h9b == r_count_20_io_out ? io_r_155_b : _GEN_4274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4276 = 8'h9c == r_count_20_io_out ? io_r_156_b : _GEN_4275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4277 = 8'h9d == r_count_20_io_out ? io_r_157_b : _GEN_4276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4278 = 8'h9e == r_count_20_io_out ? io_r_158_b : _GEN_4277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4279 = 8'h9f == r_count_20_io_out ? io_r_159_b : _GEN_4278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4280 = 8'ha0 == r_count_20_io_out ? io_r_160_b : _GEN_4279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4281 = 8'ha1 == r_count_20_io_out ? io_r_161_b : _GEN_4280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4282 = 8'ha2 == r_count_20_io_out ? io_r_162_b : _GEN_4281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4283 = 8'ha3 == r_count_20_io_out ? io_r_163_b : _GEN_4282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4284 = 8'ha4 == r_count_20_io_out ? io_r_164_b : _GEN_4283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4285 = 8'ha5 == r_count_20_io_out ? io_r_165_b : _GEN_4284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4286 = 8'ha6 == r_count_20_io_out ? io_r_166_b : _GEN_4285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4287 = 8'ha7 == r_count_20_io_out ? io_r_167_b : _GEN_4286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4288 = 8'ha8 == r_count_20_io_out ? io_r_168_b : _GEN_4287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4289 = 8'ha9 == r_count_20_io_out ? io_r_169_b : _GEN_4288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4290 = 8'haa == r_count_20_io_out ? io_r_170_b : _GEN_4289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4291 = 8'hab == r_count_20_io_out ? io_r_171_b : _GEN_4290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4292 = 8'hac == r_count_20_io_out ? io_r_172_b : _GEN_4291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4293 = 8'had == r_count_20_io_out ? io_r_173_b : _GEN_4292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4294 = 8'hae == r_count_20_io_out ? io_r_174_b : _GEN_4293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4295 = 8'haf == r_count_20_io_out ? io_r_175_b : _GEN_4294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4296 = 8'hb0 == r_count_20_io_out ? io_r_176_b : _GEN_4295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4297 = 8'hb1 == r_count_20_io_out ? io_r_177_b : _GEN_4296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4298 = 8'hb2 == r_count_20_io_out ? io_r_178_b : _GEN_4297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4299 = 8'hb3 == r_count_20_io_out ? io_r_179_b : _GEN_4298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4300 = 8'hb4 == r_count_20_io_out ? io_r_180_b : _GEN_4299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4301 = 8'hb5 == r_count_20_io_out ? io_r_181_b : _GEN_4300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4302 = 8'hb6 == r_count_20_io_out ? io_r_182_b : _GEN_4301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4303 = 8'hb7 == r_count_20_io_out ? io_r_183_b : _GEN_4302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4304 = 8'hb8 == r_count_20_io_out ? io_r_184_b : _GEN_4303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4305 = 8'hb9 == r_count_20_io_out ? io_r_185_b : _GEN_4304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4306 = 8'hba == r_count_20_io_out ? io_r_186_b : _GEN_4305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4307 = 8'hbb == r_count_20_io_out ? io_r_187_b : _GEN_4306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4308 = 8'hbc == r_count_20_io_out ? io_r_188_b : _GEN_4307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4309 = 8'hbd == r_count_20_io_out ? io_r_189_b : _GEN_4308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4310 = 8'hbe == r_count_20_io_out ? io_r_190_b : _GEN_4309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4311 = 8'hbf == r_count_20_io_out ? io_r_191_b : _GEN_4310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4312 = 8'hc0 == r_count_20_io_out ? io_r_192_b : _GEN_4311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4313 = 8'hc1 == r_count_20_io_out ? io_r_193_b : _GEN_4312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4314 = 8'hc2 == r_count_20_io_out ? io_r_194_b : _GEN_4313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4315 = 8'hc3 == r_count_20_io_out ? io_r_195_b : _GEN_4314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4316 = 8'hc4 == r_count_20_io_out ? io_r_196_b : _GEN_4315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4317 = 8'hc5 == r_count_20_io_out ? io_r_197_b : _GEN_4316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4318 = 8'hc6 == r_count_20_io_out ? io_r_198_b : _GEN_4317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4321 = 8'h1 == r_count_21_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4322 = 8'h2 == r_count_21_io_out ? io_r_2_b : _GEN_4321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4323 = 8'h3 == r_count_21_io_out ? io_r_3_b : _GEN_4322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4324 = 8'h4 == r_count_21_io_out ? io_r_4_b : _GEN_4323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4325 = 8'h5 == r_count_21_io_out ? io_r_5_b : _GEN_4324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4326 = 8'h6 == r_count_21_io_out ? io_r_6_b : _GEN_4325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4327 = 8'h7 == r_count_21_io_out ? io_r_7_b : _GEN_4326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4328 = 8'h8 == r_count_21_io_out ? io_r_8_b : _GEN_4327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4329 = 8'h9 == r_count_21_io_out ? io_r_9_b : _GEN_4328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4330 = 8'ha == r_count_21_io_out ? io_r_10_b : _GEN_4329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4331 = 8'hb == r_count_21_io_out ? io_r_11_b : _GEN_4330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4332 = 8'hc == r_count_21_io_out ? io_r_12_b : _GEN_4331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4333 = 8'hd == r_count_21_io_out ? io_r_13_b : _GEN_4332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4334 = 8'he == r_count_21_io_out ? io_r_14_b : _GEN_4333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4335 = 8'hf == r_count_21_io_out ? io_r_15_b : _GEN_4334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4336 = 8'h10 == r_count_21_io_out ? io_r_16_b : _GEN_4335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4337 = 8'h11 == r_count_21_io_out ? io_r_17_b : _GEN_4336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4338 = 8'h12 == r_count_21_io_out ? io_r_18_b : _GEN_4337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4339 = 8'h13 == r_count_21_io_out ? io_r_19_b : _GEN_4338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4340 = 8'h14 == r_count_21_io_out ? io_r_20_b : _GEN_4339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4341 = 8'h15 == r_count_21_io_out ? io_r_21_b : _GEN_4340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4342 = 8'h16 == r_count_21_io_out ? io_r_22_b : _GEN_4341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4343 = 8'h17 == r_count_21_io_out ? io_r_23_b : _GEN_4342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4344 = 8'h18 == r_count_21_io_out ? io_r_24_b : _GEN_4343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4345 = 8'h19 == r_count_21_io_out ? io_r_25_b : _GEN_4344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4346 = 8'h1a == r_count_21_io_out ? io_r_26_b : _GEN_4345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4347 = 8'h1b == r_count_21_io_out ? io_r_27_b : _GEN_4346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4348 = 8'h1c == r_count_21_io_out ? io_r_28_b : _GEN_4347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4349 = 8'h1d == r_count_21_io_out ? io_r_29_b : _GEN_4348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4350 = 8'h1e == r_count_21_io_out ? io_r_30_b : _GEN_4349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4351 = 8'h1f == r_count_21_io_out ? io_r_31_b : _GEN_4350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4352 = 8'h20 == r_count_21_io_out ? io_r_32_b : _GEN_4351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4353 = 8'h21 == r_count_21_io_out ? io_r_33_b : _GEN_4352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4354 = 8'h22 == r_count_21_io_out ? io_r_34_b : _GEN_4353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4355 = 8'h23 == r_count_21_io_out ? io_r_35_b : _GEN_4354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4356 = 8'h24 == r_count_21_io_out ? io_r_36_b : _GEN_4355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4357 = 8'h25 == r_count_21_io_out ? io_r_37_b : _GEN_4356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4358 = 8'h26 == r_count_21_io_out ? io_r_38_b : _GEN_4357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4359 = 8'h27 == r_count_21_io_out ? io_r_39_b : _GEN_4358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4360 = 8'h28 == r_count_21_io_out ? io_r_40_b : _GEN_4359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4361 = 8'h29 == r_count_21_io_out ? io_r_41_b : _GEN_4360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4362 = 8'h2a == r_count_21_io_out ? io_r_42_b : _GEN_4361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4363 = 8'h2b == r_count_21_io_out ? io_r_43_b : _GEN_4362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4364 = 8'h2c == r_count_21_io_out ? io_r_44_b : _GEN_4363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4365 = 8'h2d == r_count_21_io_out ? io_r_45_b : _GEN_4364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4366 = 8'h2e == r_count_21_io_out ? io_r_46_b : _GEN_4365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4367 = 8'h2f == r_count_21_io_out ? io_r_47_b : _GEN_4366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4368 = 8'h30 == r_count_21_io_out ? io_r_48_b : _GEN_4367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4369 = 8'h31 == r_count_21_io_out ? io_r_49_b : _GEN_4368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4370 = 8'h32 == r_count_21_io_out ? io_r_50_b : _GEN_4369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4371 = 8'h33 == r_count_21_io_out ? io_r_51_b : _GEN_4370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4372 = 8'h34 == r_count_21_io_out ? io_r_52_b : _GEN_4371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4373 = 8'h35 == r_count_21_io_out ? io_r_53_b : _GEN_4372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4374 = 8'h36 == r_count_21_io_out ? io_r_54_b : _GEN_4373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4375 = 8'h37 == r_count_21_io_out ? io_r_55_b : _GEN_4374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4376 = 8'h38 == r_count_21_io_out ? io_r_56_b : _GEN_4375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4377 = 8'h39 == r_count_21_io_out ? io_r_57_b : _GEN_4376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4378 = 8'h3a == r_count_21_io_out ? io_r_58_b : _GEN_4377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4379 = 8'h3b == r_count_21_io_out ? io_r_59_b : _GEN_4378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4380 = 8'h3c == r_count_21_io_out ? io_r_60_b : _GEN_4379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4381 = 8'h3d == r_count_21_io_out ? io_r_61_b : _GEN_4380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4382 = 8'h3e == r_count_21_io_out ? io_r_62_b : _GEN_4381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4383 = 8'h3f == r_count_21_io_out ? io_r_63_b : _GEN_4382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4384 = 8'h40 == r_count_21_io_out ? io_r_64_b : _GEN_4383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4385 = 8'h41 == r_count_21_io_out ? io_r_65_b : _GEN_4384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4386 = 8'h42 == r_count_21_io_out ? io_r_66_b : _GEN_4385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4387 = 8'h43 == r_count_21_io_out ? io_r_67_b : _GEN_4386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4388 = 8'h44 == r_count_21_io_out ? io_r_68_b : _GEN_4387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4389 = 8'h45 == r_count_21_io_out ? io_r_69_b : _GEN_4388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4390 = 8'h46 == r_count_21_io_out ? io_r_70_b : _GEN_4389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4391 = 8'h47 == r_count_21_io_out ? io_r_71_b : _GEN_4390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4392 = 8'h48 == r_count_21_io_out ? io_r_72_b : _GEN_4391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4393 = 8'h49 == r_count_21_io_out ? io_r_73_b : _GEN_4392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4394 = 8'h4a == r_count_21_io_out ? io_r_74_b : _GEN_4393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4395 = 8'h4b == r_count_21_io_out ? io_r_75_b : _GEN_4394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4396 = 8'h4c == r_count_21_io_out ? io_r_76_b : _GEN_4395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4397 = 8'h4d == r_count_21_io_out ? io_r_77_b : _GEN_4396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4398 = 8'h4e == r_count_21_io_out ? io_r_78_b : _GEN_4397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4399 = 8'h4f == r_count_21_io_out ? io_r_79_b : _GEN_4398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4400 = 8'h50 == r_count_21_io_out ? io_r_80_b : _GEN_4399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4401 = 8'h51 == r_count_21_io_out ? io_r_81_b : _GEN_4400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4402 = 8'h52 == r_count_21_io_out ? io_r_82_b : _GEN_4401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4403 = 8'h53 == r_count_21_io_out ? io_r_83_b : _GEN_4402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4404 = 8'h54 == r_count_21_io_out ? io_r_84_b : _GEN_4403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4405 = 8'h55 == r_count_21_io_out ? io_r_85_b : _GEN_4404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4406 = 8'h56 == r_count_21_io_out ? io_r_86_b : _GEN_4405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4407 = 8'h57 == r_count_21_io_out ? io_r_87_b : _GEN_4406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4408 = 8'h58 == r_count_21_io_out ? io_r_88_b : _GEN_4407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4409 = 8'h59 == r_count_21_io_out ? io_r_89_b : _GEN_4408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4410 = 8'h5a == r_count_21_io_out ? io_r_90_b : _GEN_4409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4411 = 8'h5b == r_count_21_io_out ? io_r_91_b : _GEN_4410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4412 = 8'h5c == r_count_21_io_out ? io_r_92_b : _GEN_4411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4413 = 8'h5d == r_count_21_io_out ? io_r_93_b : _GEN_4412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4414 = 8'h5e == r_count_21_io_out ? io_r_94_b : _GEN_4413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4415 = 8'h5f == r_count_21_io_out ? io_r_95_b : _GEN_4414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4416 = 8'h60 == r_count_21_io_out ? io_r_96_b : _GEN_4415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4417 = 8'h61 == r_count_21_io_out ? io_r_97_b : _GEN_4416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4418 = 8'h62 == r_count_21_io_out ? io_r_98_b : _GEN_4417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4419 = 8'h63 == r_count_21_io_out ? io_r_99_b : _GEN_4418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4420 = 8'h64 == r_count_21_io_out ? io_r_100_b : _GEN_4419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4421 = 8'h65 == r_count_21_io_out ? io_r_101_b : _GEN_4420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4422 = 8'h66 == r_count_21_io_out ? io_r_102_b : _GEN_4421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4423 = 8'h67 == r_count_21_io_out ? io_r_103_b : _GEN_4422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4424 = 8'h68 == r_count_21_io_out ? io_r_104_b : _GEN_4423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4425 = 8'h69 == r_count_21_io_out ? io_r_105_b : _GEN_4424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4426 = 8'h6a == r_count_21_io_out ? io_r_106_b : _GEN_4425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4427 = 8'h6b == r_count_21_io_out ? io_r_107_b : _GEN_4426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4428 = 8'h6c == r_count_21_io_out ? io_r_108_b : _GEN_4427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4429 = 8'h6d == r_count_21_io_out ? io_r_109_b : _GEN_4428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4430 = 8'h6e == r_count_21_io_out ? io_r_110_b : _GEN_4429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4431 = 8'h6f == r_count_21_io_out ? io_r_111_b : _GEN_4430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4432 = 8'h70 == r_count_21_io_out ? io_r_112_b : _GEN_4431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4433 = 8'h71 == r_count_21_io_out ? io_r_113_b : _GEN_4432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4434 = 8'h72 == r_count_21_io_out ? io_r_114_b : _GEN_4433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4435 = 8'h73 == r_count_21_io_out ? io_r_115_b : _GEN_4434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4436 = 8'h74 == r_count_21_io_out ? io_r_116_b : _GEN_4435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4437 = 8'h75 == r_count_21_io_out ? io_r_117_b : _GEN_4436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4438 = 8'h76 == r_count_21_io_out ? io_r_118_b : _GEN_4437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4439 = 8'h77 == r_count_21_io_out ? io_r_119_b : _GEN_4438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4440 = 8'h78 == r_count_21_io_out ? io_r_120_b : _GEN_4439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4441 = 8'h79 == r_count_21_io_out ? io_r_121_b : _GEN_4440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4442 = 8'h7a == r_count_21_io_out ? io_r_122_b : _GEN_4441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4443 = 8'h7b == r_count_21_io_out ? io_r_123_b : _GEN_4442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4444 = 8'h7c == r_count_21_io_out ? io_r_124_b : _GEN_4443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4445 = 8'h7d == r_count_21_io_out ? io_r_125_b : _GEN_4444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4446 = 8'h7e == r_count_21_io_out ? io_r_126_b : _GEN_4445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4447 = 8'h7f == r_count_21_io_out ? io_r_127_b : _GEN_4446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4448 = 8'h80 == r_count_21_io_out ? io_r_128_b : _GEN_4447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4449 = 8'h81 == r_count_21_io_out ? io_r_129_b : _GEN_4448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4450 = 8'h82 == r_count_21_io_out ? io_r_130_b : _GEN_4449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4451 = 8'h83 == r_count_21_io_out ? io_r_131_b : _GEN_4450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4452 = 8'h84 == r_count_21_io_out ? io_r_132_b : _GEN_4451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4453 = 8'h85 == r_count_21_io_out ? io_r_133_b : _GEN_4452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4454 = 8'h86 == r_count_21_io_out ? io_r_134_b : _GEN_4453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4455 = 8'h87 == r_count_21_io_out ? io_r_135_b : _GEN_4454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4456 = 8'h88 == r_count_21_io_out ? io_r_136_b : _GEN_4455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4457 = 8'h89 == r_count_21_io_out ? io_r_137_b : _GEN_4456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4458 = 8'h8a == r_count_21_io_out ? io_r_138_b : _GEN_4457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4459 = 8'h8b == r_count_21_io_out ? io_r_139_b : _GEN_4458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4460 = 8'h8c == r_count_21_io_out ? io_r_140_b : _GEN_4459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4461 = 8'h8d == r_count_21_io_out ? io_r_141_b : _GEN_4460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4462 = 8'h8e == r_count_21_io_out ? io_r_142_b : _GEN_4461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4463 = 8'h8f == r_count_21_io_out ? io_r_143_b : _GEN_4462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4464 = 8'h90 == r_count_21_io_out ? io_r_144_b : _GEN_4463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4465 = 8'h91 == r_count_21_io_out ? io_r_145_b : _GEN_4464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4466 = 8'h92 == r_count_21_io_out ? io_r_146_b : _GEN_4465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4467 = 8'h93 == r_count_21_io_out ? io_r_147_b : _GEN_4466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4468 = 8'h94 == r_count_21_io_out ? io_r_148_b : _GEN_4467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4469 = 8'h95 == r_count_21_io_out ? io_r_149_b : _GEN_4468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4470 = 8'h96 == r_count_21_io_out ? io_r_150_b : _GEN_4469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4471 = 8'h97 == r_count_21_io_out ? io_r_151_b : _GEN_4470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4472 = 8'h98 == r_count_21_io_out ? io_r_152_b : _GEN_4471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4473 = 8'h99 == r_count_21_io_out ? io_r_153_b : _GEN_4472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4474 = 8'h9a == r_count_21_io_out ? io_r_154_b : _GEN_4473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4475 = 8'h9b == r_count_21_io_out ? io_r_155_b : _GEN_4474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4476 = 8'h9c == r_count_21_io_out ? io_r_156_b : _GEN_4475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4477 = 8'h9d == r_count_21_io_out ? io_r_157_b : _GEN_4476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4478 = 8'h9e == r_count_21_io_out ? io_r_158_b : _GEN_4477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4479 = 8'h9f == r_count_21_io_out ? io_r_159_b : _GEN_4478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4480 = 8'ha0 == r_count_21_io_out ? io_r_160_b : _GEN_4479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4481 = 8'ha1 == r_count_21_io_out ? io_r_161_b : _GEN_4480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4482 = 8'ha2 == r_count_21_io_out ? io_r_162_b : _GEN_4481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4483 = 8'ha3 == r_count_21_io_out ? io_r_163_b : _GEN_4482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4484 = 8'ha4 == r_count_21_io_out ? io_r_164_b : _GEN_4483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4485 = 8'ha5 == r_count_21_io_out ? io_r_165_b : _GEN_4484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4486 = 8'ha6 == r_count_21_io_out ? io_r_166_b : _GEN_4485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4487 = 8'ha7 == r_count_21_io_out ? io_r_167_b : _GEN_4486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4488 = 8'ha8 == r_count_21_io_out ? io_r_168_b : _GEN_4487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4489 = 8'ha9 == r_count_21_io_out ? io_r_169_b : _GEN_4488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4490 = 8'haa == r_count_21_io_out ? io_r_170_b : _GEN_4489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4491 = 8'hab == r_count_21_io_out ? io_r_171_b : _GEN_4490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4492 = 8'hac == r_count_21_io_out ? io_r_172_b : _GEN_4491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4493 = 8'had == r_count_21_io_out ? io_r_173_b : _GEN_4492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4494 = 8'hae == r_count_21_io_out ? io_r_174_b : _GEN_4493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4495 = 8'haf == r_count_21_io_out ? io_r_175_b : _GEN_4494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4496 = 8'hb0 == r_count_21_io_out ? io_r_176_b : _GEN_4495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4497 = 8'hb1 == r_count_21_io_out ? io_r_177_b : _GEN_4496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4498 = 8'hb2 == r_count_21_io_out ? io_r_178_b : _GEN_4497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4499 = 8'hb3 == r_count_21_io_out ? io_r_179_b : _GEN_4498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4500 = 8'hb4 == r_count_21_io_out ? io_r_180_b : _GEN_4499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4501 = 8'hb5 == r_count_21_io_out ? io_r_181_b : _GEN_4500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4502 = 8'hb6 == r_count_21_io_out ? io_r_182_b : _GEN_4501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4503 = 8'hb7 == r_count_21_io_out ? io_r_183_b : _GEN_4502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4504 = 8'hb8 == r_count_21_io_out ? io_r_184_b : _GEN_4503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4505 = 8'hb9 == r_count_21_io_out ? io_r_185_b : _GEN_4504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4506 = 8'hba == r_count_21_io_out ? io_r_186_b : _GEN_4505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4507 = 8'hbb == r_count_21_io_out ? io_r_187_b : _GEN_4506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4508 = 8'hbc == r_count_21_io_out ? io_r_188_b : _GEN_4507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4509 = 8'hbd == r_count_21_io_out ? io_r_189_b : _GEN_4508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4510 = 8'hbe == r_count_21_io_out ? io_r_190_b : _GEN_4509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4511 = 8'hbf == r_count_21_io_out ? io_r_191_b : _GEN_4510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4512 = 8'hc0 == r_count_21_io_out ? io_r_192_b : _GEN_4511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4513 = 8'hc1 == r_count_21_io_out ? io_r_193_b : _GEN_4512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4514 = 8'hc2 == r_count_21_io_out ? io_r_194_b : _GEN_4513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4515 = 8'hc3 == r_count_21_io_out ? io_r_195_b : _GEN_4514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4516 = 8'hc4 == r_count_21_io_out ? io_r_196_b : _GEN_4515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4517 = 8'hc5 == r_count_21_io_out ? io_r_197_b : _GEN_4516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4518 = 8'hc6 == r_count_21_io_out ? io_r_198_b : _GEN_4517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4521 = 8'h1 == r_count_22_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4522 = 8'h2 == r_count_22_io_out ? io_r_2_b : _GEN_4521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4523 = 8'h3 == r_count_22_io_out ? io_r_3_b : _GEN_4522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4524 = 8'h4 == r_count_22_io_out ? io_r_4_b : _GEN_4523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4525 = 8'h5 == r_count_22_io_out ? io_r_5_b : _GEN_4524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4526 = 8'h6 == r_count_22_io_out ? io_r_6_b : _GEN_4525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4527 = 8'h7 == r_count_22_io_out ? io_r_7_b : _GEN_4526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4528 = 8'h8 == r_count_22_io_out ? io_r_8_b : _GEN_4527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4529 = 8'h9 == r_count_22_io_out ? io_r_9_b : _GEN_4528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4530 = 8'ha == r_count_22_io_out ? io_r_10_b : _GEN_4529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4531 = 8'hb == r_count_22_io_out ? io_r_11_b : _GEN_4530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4532 = 8'hc == r_count_22_io_out ? io_r_12_b : _GEN_4531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4533 = 8'hd == r_count_22_io_out ? io_r_13_b : _GEN_4532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4534 = 8'he == r_count_22_io_out ? io_r_14_b : _GEN_4533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4535 = 8'hf == r_count_22_io_out ? io_r_15_b : _GEN_4534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4536 = 8'h10 == r_count_22_io_out ? io_r_16_b : _GEN_4535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4537 = 8'h11 == r_count_22_io_out ? io_r_17_b : _GEN_4536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4538 = 8'h12 == r_count_22_io_out ? io_r_18_b : _GEN_4537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4539 = 8'h13 == r_count_22_io_out ? io_r_19_b : _GEN_4538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4540 = 8'h14 == r_count_22_io_out ? io_r_20_b : _GEN_4539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4541 = 8'h15 == r_count_22_io_out ? io_r_21_b : _GEN_4540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4542 = 8'h16 == r_count_22_io_out ? io_r_22_b : _GEN_4541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4543 = 8'h17 == r_count_22_io_out ? io_r_23_b : _GEN_4542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4544 = 8'h18 == r_count_22_io_out ? io_r_24_b : _GEN_4543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4545 = 8'h19 == r_count_22_io_out ? io_r_25_b : _GEN_4544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4546 = 8'h1a == r_count_22_io_out ? io_r_26_b : _GEN_4545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4547 = 8'h1b == r_count_22_io_out ? io_r_27_b : _GEN_4546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4548 = 8'h1c == r_count_22_io_out ? io_r_28_b : _GEN_4547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4549 = 8'h1d == r_count_22_io_out ? io_r_29_b : _GEN_4548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4550 = 8'h1e == r_count_22_io_out ? io_r_30_b : _GEN_4549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4551 = 8'h1f == r_count_22_io_out ? io_r_31_b : _GEN_4550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4552 = 8'h20 == r_count_22_io_out ? io_r_32_b : _GEN_4551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4553 = 8'h21 == r_count_22_io_out ? io_r_33_b : _GEN_4552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4554 = 8'h22 == r_count_22_io_out ? io_r_34_b : _GEN_4553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4555 = 8'h23 == r_count_22_io_out ? io_r_35_b : _GEN_4554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4556 = 8'h24 == r_count_22_io_out ? io_r_36_b : _GEN_4555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4557 = 8'h25 == r_count_22_io_out ? io_r_37_b : _GEN_4556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4558 = 8'h26 == r_count_22_io_out ? io_r_38_b : _GEN_4557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4559 = 8'h27 == r_count_22_io_out ? io_r_39_b : _GEN_4558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4560 = 8'h28 == r_count_22_io_out ? io_r_40_b : _GEN_4559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4561 = 8'h29 == r_count_22_io_out ? io_r_41_b : _GEN_4560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4562 = 8'h2a == r_count_22_io_out ? io_r_42_b : _GEN_4561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4563 = 8'h2b == r_count_22_io_out ? io_r_43_b : _GEN_4562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4564 = 8'h2c == r_count_22_io_out ? io_r_44_b : _GEN_4563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4565 = 8'h2d == r_count_22_io_out ? io_r_45_b : _GEN_4564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4566 = 8'h2e == r_count_22_io_out ? io_r_46_b : _GEN_4565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4567 = 8'h2f == r_count_22_io_out ? io_r_47_b : _GEN_4566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4568 = 8'h30 == r_count_22_io_out ? io_r_48_b : _GEN_4567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4569 = 8'h31 == r_count_22_io_out ? io_r_49_b : _GEN_4568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4570 = 8'h32 == r_count_22_io_out ? io_r_50_b : _GEN_4569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4571 = 8'h33 == r_count_22_io_out ? io_r_51_b : _GEN_4570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4572 = 8'h34 == r_count_22_io_out ? io_r_52_b : _GEN_4571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4573 = 8'h35 == r_count_22_io_out ? io_r_53_b : _GEN_4572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4574 = 8'h36 == r_count_22_io_out ? io_r_54_b : _GEN_4573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4575 = 8'h37 == r_count_22_io_out ? io_r_55_b : _GEN_4574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4576 = 8'h38 == r_count_22_io_out ? io_r_56_b : _GEN_4575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4577 = 8'h39 == r_count_22_io_out ? io_r_57_b : _GEN_4576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4578 = 8'h3a == r_count_22_io_out ? io_r_58_b : _GEN_4577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4579 = 8'h3b == r_count_22_io_out ? io_r_59_b : _GEN_4578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4580 = 8'h3c == r_count_22_io_out ? io_r_60_b : _GEN_4579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4581 = 8'h3d == r_count_22_io_out ? io_r_61_b : _GEN_4580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4582 = 8'h3e == r_count_22_io_out ? io_r_62_b : _GEN_4581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4583 = 8'h3f == r_count_22_io_out ? io_r_63_b : _GEN_4582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4584 = 8'h40 == r_count_22_io_out ? io_r_64_b : _GEN_4583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4585 = 8'h41 == r_count_22_io_out ? io_r_65_b : _GEN_4584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4586 = 8'h42 == r_count_22_io_out ? io_r_66_b : _GEN_4585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4587 = 8'h43 == r_count_22_io_out ? io_r_67_b : _GEN_4586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4588 = 8'h44 == r_count_22_io_out ? io_r_68_b : _GEN_4587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4589 = 8'h45 == r_count_22_io_out ? io_r_69_b : _GEN_4588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4590 = 8'h46 == r_count_22_io_out ? io_r_70_b : _GEN_4589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4591 = 8'h47 == r_count_22_io_out ? io_r_71_b : _GEN_4590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4592 = 8'h48 == r_count_22_io_out ? io_r_72_b : _GEN_4591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4593 = 8'h49 == r_count_22_io_out ? io_r_73_b : _GEN_4592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4594 = 8'h4a == r_count_22_io_out ? io_r_74_b : _GEN_4593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4595 = 8'h4b == r_count_22_io_out ? io_r_75_b : _GEN_4594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4596 = 8'h4c == r_count_22_io_out ? io_r_76_b : _GEN_4595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4597 = 8'h4d == r_count_22_io_out ? io_r_77_b : _GEN_4596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4598 = 8'h4e == r_count_22_io_out ? io_r_78_b : _GEN_4597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4599 = 8'h4f == r_count_22_io_out ? io_r_79_b : _GEN_4598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4600 = 8'h50 == r_count_22_io_out ? io_r_80_b : _GEN_4599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4601 = 8'h51 == r_count_22_io_out ? io_r_81_b : _GEN_4600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4602 = 8'h52 == r_count_22_io_out ? io_r_82_b : _GEN_4601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4603 = 8'h53 == r_count_22_io_out ? io_r_83_b : _GEN_4602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4604 = 8'h54 == r_count_22_io_out ? io_r_84_b : _GEN_4603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4605 = 8'h55 == r_count_22_io_out ? io_r_85_b : _GEN_4604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4606 = 8'h56 == r_count_22_io_out ? io_r_86_b : _GEN_4605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4607 = 8'h57 == r_count_22_io_out ? io_r_87_b : _GEN_4606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4608 = 8'h58 == r_count_22_io_out ? io_r_88_b : _GEN_4607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4609 = 8'h59 == r_count_22_io_out ? io_r_89_b : _GEN_4608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4610 = 8'h5a == r_count_22_io_out ? io_r_90_b : _GEN_4609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4611 = 8'h5b == r_count_22_io_out ? io_r_91_b : _GEN_4610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4612 = 8'h5c == r_count_22_io_out ? io_r_92_b : _GEN_4611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4613 = 8'h5d == r_count_22_io_out ? io_r_93_b : _GEN_4612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4614 = 8'h5e == r_count_22_io_out ? io_r_94_b : _GEN_4613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4615 = 8'h5f == r_count_22_io_out ? io_r_95_b : _GEN_4614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4616 = 8'h60 == r_count_22_io_out ? io_r_96_b : _GEN_4615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4617 = 8'h61 == r_count_22_io_out ? io_r_97_b : _GEN_4616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4618 = 8'h62 == r_count_22_io_out ? io_r_98_b : _GEN_4617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4619 = 8'h63 == r_count_22_io_out ? io_r_99_b : _GEN_4618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4620 = 8'h64 == r_count_22_io_out ? io_r_100_b : _GEN_4619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4621 = 8'h65 == r_count_22_io_out ? io_r_101_b : _GEN_4620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4622 = 8'h66 == r_count_22_io_out ? io_r_102_b : _GEN_4621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4623 = 8'h67 == r_count_22_io_out ? io_r_103_b : _GEN_4622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4624 = 8'h68 == r_count_22_io_out ? io_r_104_b : _GEN_4623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4625 = 8'h69 == r_count_22_io_out ? io_r_105_b : _GEN_4624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4626 = 8'h6a == r_count_22_io_out ? io_r_106_b : _GEN_4625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4627 = 8'h6b == r_count_22_io_out ? io_r_107_b : _GEN_4626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4628 = 8'h6c == r_count_22_io_out ? io_r_108_b : _GEN_4627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4629 = 8'h6d == r_count_22_io_out ? io_r_109_b : _GEN_4628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4630 = 8'h6e == r_count_22_io_out ? io_r_110_b : _GEN_4629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4631 = 8'h6f == r_count_22_io_out ? io_r_111_b : _GEN_4630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4632 = 8'h70 == r_count_22_io_out ? io_r_112_b : _GEN_4631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4633 = 8'h71 == r_count_22_io_out ? io_r_113_b : _GEN_4632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4634 = 8'h72 == r_count_22_io_out ? io_r_114_b : _GEN_4633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4635 = 8'h73 == r_count_22_io_out ? io_r_115_b : _GEN_4634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4636 = 8'h74 == r_count_22_io_out ? io_r_116_b : _GEN_4635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4637 = 8'h75 == r_count_22_io_out ? io_r_117_b : _GEN_4636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4638 = 8'h76 == r_count_22_io_out ? io_r_118_b : _GEN_4637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4639 = 8'h77 == r_count_22_io_out ? io_r_119_b : _GEN_4638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4640 = 8'h78 == r_count_22_io_out ? io_r_120_b : _GEN_4639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4641 = 8'h79 == r_count_22_io_out ? io_r_121_b : _GEN_4640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4642 = 8'h7a == r_count_22_io_out ? io_r_122_b : _GEN_4641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4643 = 8'h7b == r_count_22_io_out ? io_r_123_b : _GEN_4642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4644 = 8'h7c == r_count_22_io_out ? io_r_124_b : _GEN_4643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4645 = 8'h7d == r_count_22_io_out ? io_r_125_b : _GEN_4644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4646 = 8'h7e == r_count_22_io_out ? io_r_126_b : _GEN_4645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4647 = 8'h7f == r_count_22_io_out ? io_r_127_b : _GEN_4646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4648 = 8'h80 == r_count_22_io_out ? io_r_128_b : _GEN_4647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4649 = 8'h81 == r_count_22_io_out ? io_r_129_b : _GEN_4648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4650 = 8'h82 == r_count_22_io_out ? io_r_130_b : _GEN_4649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4651 = 8'h83 == r_count_22_io_out ? io_r_131_b : _GEN_4650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4652 = 8'h84 == r_count_22_io_out ? io_r_132_b : _GEN_4651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4653 = 8'h85 == r_count_22_io_out ? io_r_133_b : _GEN_4652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4654 = 8'h86 == r_count_22_io_out ? io_r_134_b : _GEN_4653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4655 = 8'h87 == r_count_22_io_out ? io_r_135_b : _GEN_4654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4656 = 8'h88 == r_count_22_io_out ? io_r_136_b : _GEN_4655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4657 = 8'h89 == r_count_22_io_out ? io_r_137_b : _GEN_4656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4658 = 8'h8a == r_count_22_io_out ? io_r_138_b : _GEN_4657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4659 = 8'h8b == r_count_22_io_out ? io_r_139_b : _GEN_4658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4660 = 8'h8c == r_count_22_io_out ? io_r_140_b : _GEN_4659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4661 = 8'h8d == r_count_22_io_out ? io_r_141_b : _GEN_4660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4662 = 8'h8e == r_count_22_io_out ? io_r_142_b : _GEN_4661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4663 = 8'h8f == r_count_22_io_out ? io_r_143_b : _GEN_4662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4664 = 8'h90 == r_count_22_io_out ? io_r_144_b : _GEN_4663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4665 = 8'h91 == r_count_22_io_out ? io_r_145_b : _GEN_4664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4666 = 8'h92 == r_count_22_io_out ? io_r_146_b : _GEN_4665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4667 = 8'h93 == r_count_22_io_out ? io_r_147_b : _GEN_4666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4668 = 8'h94 == r_count_22_io_out ? io_r_148_b : _GEN_4667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4669 = 8'h95 == r_count_22_io_out ? io_r_149_b : _GEN_4668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4670 = 8'h96 == r_count_22_io_out ? io_r_150_b : _GEN_4669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4671 = 8'h97 == r_count_22_io_out ? io_r_151_b : _GEN_4670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4672 = 8'h98 == r_count_22_io_out ? io_r_152_b : _GEN_4671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4673 = 8'h99 == r_count_22_io_out ? io_r_153_b : _GEN_4672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4674 = 8'h9a == r_count_22_io_out ? io_r_154_b : _GEN_4673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4675 = 8'h9b == r_count_22_io_out ? io_r_155_b : _GEN_4674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4676 = 8'h9c == r_count_22_io_out ? io_r_156_b : _GEN_4675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4677 = 8'h9d == r_count_22_io_out ? io_r_157_b : _GEN_4676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4678 = 8'h9e == r_count_22_io_out ? io_r_158_b : _GEN_4677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4679 = 8'h9f == r_count_22_io_out ? io_r_159_b : _GEN_4678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4680 = 8'ha0 == r_count_22_io_out ? io_r_160_b : _GEN_4679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4681 = 8'ha1 == r_count_22_io_out ? io_r_161_b : _GEN_4680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4682 = 8'ha2 == r_count_22_io_out ? io_r_162_b : _GEN_4681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4683 = 8'ha3 == r_count_22_io_out ? io_r_163_b : _GEN_4682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4684 = 8'ha4 == r_count_22_io_out ? io_r_164_b : _GEN_4683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4685 = 8'ha5 == r_count_22_io_out ? io_r_165_b : _GEN_4684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4686 = 8'ha6 == r_count_22_io_out ? io_r_166_b : _GEN_4685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4687 = 8'ha7 == r_count_22_io_out ? io_r_167_b : _GEN_4686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4688 = 8'ha8 == r_count_22_io_out ? io_r_168_b : _GEN_4687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4689 = 8'ha9 == r_count_22_io_out ? io_r_169_b : _GEN_4688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4690 = 8'haa == r_count_22_io_out ? io_r_170_b : _GEN_4689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4691 = 8'hab == r_count_22_io_out ? io_r_171_b : _GEN_4690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4692 = 8'hac == r_count_22_io_out ? io_r_172_b : _GEN_4691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4693 = 8'had == r_count_22_io_out ? io_r_173_b : _GEN_4692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4694 = 8'hae == r_count_22_io_out ? io_r_174_b : _GEN_4693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4695 = 8'haf == r_count_22_io_out ? io_r_175_b : _GEN_4694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4696 = 8'hb0 == r_count_22_io_out ? io_r_176_b : _GEN_4695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4697 = 8'hb1 == r_count_22_io_out ? io_r_177_b : _GEN_4696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4698 = 8'hb2 == r_count_22_io_out ? io_r_178_b : _GEN_4697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4699 = 8'hb3 == r_count_22_io_out ? io_r_179_b : _GEN_4698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4700 = 8'hb4 == r_count_22_io_out ? io_r_180_b : _GEN_4699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4701 = 8'hb5 == r_count_22_io_out ? io_r_181_b : _GEN_4700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4702 = 8'hb6 == r_count_22_io_out ? io_r_182_b : _GEN_4701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4703 = 8'hb7 == r_count_22_io_out ? io_r_183_b : _GEN_4702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4704 = 8'hb8 == r_count_22_io_out ? io_r_184_b : _GEN_4703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4705 = 8'hb9 == r_count_22_io_out ? io_r_185_b : _GEN_4704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4706 = 8'hba == r_count_22_io_out ? io_r_186_b : _GEN_4705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4707 = 8'hbb == r_count_22_io_out ? io_r_187_b : _GEN_4706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4708 = 8'hbc == r_count_22_io_out ? io_r_188_b : _GEN_4707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4709 = 8'hbd == r_count_22_io_out ? io_r_189_b : _GEN_4708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4710 = 8'hbe == r_count_22_io_out ? io_r_190_b : _GEN_4709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4711 = 8'hbf == r_count_22_io_out ? io_r_191_b : _GEN_4710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4712 = 8'hc0 == r_count_22_io_out ? io_r_192_b : _GEN_4711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4713 = 8'hc1 == r_count_22_io_out ? io_r_193_b : _GEN_4712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4714 = 8'hc2 == r_count_22_io_out ? io_r_194_b : _GEN_4713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4715 = 8'hc3 == r_count_22_io_out ? io_r_195_b : _GEN_4714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4716 = 8'hc4 == r_count_22_io_out ? io_r_196_b : _GEN_4715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4717 = 8'hc5 == r_count_22_io_out ? io_r_197_b : _GEN_4716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4718 = 8'hc6 == r_count_22_io_out ? io_r_198_b : _GEN_4717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4721 = 8'h1 == r_count_23_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4722 = 8'h2 == r_count_23_io_out ? io_r_2_b : _GEN_4721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4723 = 8'h3 == r_count_23_io_out ? io_r_3_b : _GEN_4722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4724 = 8'h4 == r_count_23_io_out ? io_r_4_b : _GEN_4723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4725 = 8'h5 == r_count_23_io_out ? io_r_5_b : _GEN_4724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4726 = 8'h6 == r_count_23_io_out ? io_r_6_b : _GEN_4725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4727 = 8'h7 == r_count_23_io_out ? io_r_7_b : _GEN_4726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4728 = 8'h8 == r_count_23_io_out ? io_r_8_b : _GEN_4727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4729 = 8'h9 == r_count_23_io_out ? io_r_9_b : _GEN_4728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4730 = 8'ha == r_count_23_io_out ? io_r_10_b : _GEN_4729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4731 = 8'hb == r_count_23_io_out ? io_r_11_b : _GEN_4730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4732 = 8'hc == r_count_23_io_out ? io_r_12_b : _GEN_4731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4733 = 8'hd == r_count_23_io_out ? io_r_13_b : _GEN_4732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4734 = 8'he == r_count_23_io_out ? io_r_14_b : _GEN_4733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4735 = 8'hf == r_count_23_io_out ? io_r_15_b : _GEN_4734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4736 = 8'h10 == r_count_23_io_out ? io_r_16_b : _GEN_4735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4737 = 8'h11 == r_count_23_io_out ? io_r_17_b : _GEN_4736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4738 = 8'h12 == r_count_23_io_out ? io_r_18_b : _GEN_4737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4739 = 8'h13 == r_count_23_io_out ? io_r_19_b : _GEN_4738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4740 = 8'h14 == r_count_23_io_out ? io_r_20_b : _GEN_4739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4741 = 8'h15 == r_count_23_io_out ? io_r_21_b : _GEN_4740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4742 = 8'h16 == r_count_23_io_out ? io_r_22_b : _GEN_4741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4743 = 8'h17 == r_count_23_io_out ? io_r_23_b : _GEN_4742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4744 = 8'h18 == r_count_23_io_out ? io_r_24_b : _GEN_4743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4745 = 8'h19 == r_count_23_io_out ? io_r_25_b : _GEN_4744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4746 = 8'h1a == r_count_23_io_out ? io_r_26_b : _GEN_4745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4747 = 8'h1b == r_count_23_io_out ? io_r_27_b : _GEN_4746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4748 = 8'h1c == r_count_23_io_out ? io_r_28_b : _GEN_4747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4749 = 8'h1d == r_count_23_io_out ? io_r_29_b : _GEN_4748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4750 = 8'h1e == r_count_23_io_out ? io_r_30_b : _GEN_4749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4751 = 8'h1f == r_count_23_io_out ? io_r_31_b : _GEN_4750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4752 = 8'h20 == r_count_23_io_out ? io_r_32_b : _GEN_4751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4753 = 8'h21 == r_count_23_io_out ? io_r_33_b : _GEN_4752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4754 = 8'h22 == r_count_23_io_out ? io_r_34_b : _GEN_4753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4755 = 8'h23 == r_count_23_io_out ? io_r_35_b : _GEN_4754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4756 = 8'h24 == r_count_23_io_out ? io_r_36_b : _GEN_4755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4757 = 8'h25 == r_count_23_io_out ? io_r_37_b : _GEN_4756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4758 = 8'h26 == r_count_23_io_out ? io_r_38_b : _GEN_4757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4759 = 8'h27 == r_count_23_io_out ? io_r_39_b : _GEN_4758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4760 = 8'h28 == r_count_23_io_out ? io_r_40_b : _GEN_4759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4761 = 8'h29 == r_count_23_io_out ? io_r_41_b : _GEN_4760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4762 = 8'h2a == r_count_23_io_out ? io_r_42_b : _GEN_4761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4763 = 8'h2b == r_count_23_io_out ? io_r_43_b : _GEN_4762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4764 = 8'h2c == r_count_23_io_out ? io_r_44_b : _GEN_4763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4765 = 8'h2d == r_count_23_io_out ? io_r_45_b : _GEN_4764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4766 = 8'h2e == r_count_23_io_out ? io_r_46_b : _GEN_4765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4767 = 8'h2f == r_count_23_io_out ? io_r_47_b : _GEN_4766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4768 = 8'h30 == r_count_23_io_out ? io_r_48_b : _GEN_4767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4769 = 8'h31 == r_count_23_io_out ? io_r_49_b : _GEN_4768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4770 = 8'h32 == r_count_23_io_out ? io_r_50_b : _GEN_4769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4771 = 8'h33 == r_count_23_io_out ? io_r_51_b : _GEN_4770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4772 = 8'h34 == r_count_23_io_out ? io_r_52_b : _GEN_4771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4773 = 8'h35 == r_count_23_io_out ? io_r_53_b : _GEN_4772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4774 = 8'h36 == r_count_23_io_out ? io_r_54_b : _GEN_4773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4775 = 8'h37 == r_count_23_io_out ? io_r_55_b : _GEN_4774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4776 = 8'h38 == r_count_23_io_out ? io_r_56_b : _GEN_4775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4777 = 8'h39 == r_count_23_io_out ? io_r_57_b : _GEN_4776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4778 = 8'h3a == r_count_23_io_out ? io_r_58_b : _GEN_4777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4779 = 8'h3b == r_count_23_io_out ? io_r_59_b : _GEN_4778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4780 = 8'h3c == r_count_23_io_out ? io_r_60_b : _GEN_4779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4781 = 8'h3d == r_count_23_io_out ? io_r_61_b : _GEN_4780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4782 = 8'h3e == r_count_23_io_out ? io_r_62_b : _GEN_4781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4783 = 8'h3f == r_count_23_io_out ? io_r_63_b : _GEN_4782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4784 = 8'h40 == r_count_23_io_out ? io_r_64_b : _GEN_4783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4785 = 8'h41 == r_count_23_io_out ? io_r_65_b : _GEN_4784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4786 = 8'h42 == r_count_23_io_out ? io_r_66_b : _GEN_4785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4787 = 8'h43 == r_count_23_io_out ? io_r_67_b : _GEN_4786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4788 = 8'h44 == r_count_23_io_out ? io_r_68_b : _GEN_4787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4789 = 8'h45 == r_count_23_io_out ? io_r_69_b : _GEN_4788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4790 = 8'h46 == r_count_23_io_out ? io_r_70_b : _GEN_4789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4791 = 8'h47 == r_count_23_io_out ? io_r_71_b : _GEN_4790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4792 = 8'h48 == r_count_23_io_out ? io_r_72_b : _GEN_4791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4793 = 8'h49 == r_count_23_io_out ? io_r_73_b : _GEN_4792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4794 = 8'h4a == r_count_23_io_out ? io_r_74_b : _GEN_4793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4795 = 8'h4b == r_count_23_io_out ? io_r_75_b : _GEN_4794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4796 = 8'h4c == r_count_23_io_out ? io_r_76_b : _GEN_4795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4797 = 8'h4d == r_count_23_io_out ? io_r_77_b : _GEN_4796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4798 = 8'h4e == r_count_23_io_out ? io_r_78_b : _GEN_4797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4799 = 8'h4f == r_count_23_io_out ? io_r_79_b : _GEN_4798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4800 = 8'h50 == r_count_23_io_out ? io_r_80_b : _GEN_4799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4801 = 8'h51 == r_count_23_io_out ? io_r_81_b : _GEN_4800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4802 = 8'h52 == r_count_23_io_out ? io_r_82_b : _GEN_4801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4803 = 8'h53 == r_count_23_io_out ? io_r_83_b : _GEN_4802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4804 = 8'h54 == r_count_23_io_out ? io_r_84_b : _GEN_4803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4805 = 8'h55 == r_count_23_io_out ? io_r_85_b : _GEN_4804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4806 = 8'h56 == r_count_23_io_out ? io_r_86_b : _GEN_4805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4807 = 8'h57 == r_count_23_io_out ? io_r_87_b : _GEN_4806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4808 = 8'h58 == r_count_23_io_out ? io_r_88_b : _GEN_4807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4809 = 8'h59 == r_count_23_io_out ? io_r_89_b : _GEN_4808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4810 = 8'h5a == r_count_23_io_out ? io_r_90_b : _GEN_4809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4811 = 8'h5b == r_count_23_io_out ? io_r_91_b : _GEN_4810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4812 = 8'h5c == r_count_23_io_out ? io_r_92_b : _GEN_4811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4813 = 8'h5d == r_count_23_io_out ? io_r_93_b : _GEN_4812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4814 = 8'h5e == r_count_23_io_out ? io_r_94_b : _GEN_4813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4815 = 8'h5f == r_count_23_io_out ? io_r_95_b : _GEN_4814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4816 = 8'h60 == r_count_23_io_out ? io_r_96_b : _GEN_4815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4817 = 8'h61 == r_count_23_io_out ? io_r_97_b : _GEN_4816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4818 = 8'h62 == r_count_23_io_out ? io_r_98_b : _GEN_4817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4819 = 8'h63 == r_count_23_io_out ? io_r_99_b : _GEN_4818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4820 = 8'h64 == r_count_23_io_out ? io_r_100_b : _GEN_4819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4821 = 8'h65 == r_count_23_io_out ? io_r_101_b : _GEN_4820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4822 = 8'h66 == r_count_23_io_out ? io_r_102_b : _GEN_4821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4823 = 8'h67 == r_count_23_io_out ? io_r_103_b : _GEN_4822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4824 = 8'h68 == r_count_23_io_out ? io_r_104_b : _GEN_4823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4825 = 8'h69 == r_count_23_io_out ? io_r_105_b : _GEN_4824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4826 = 8'h6a == r_count_23_io_out ? io_r_106_b : _GEN_4825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4827 = 8'h6b == r_count_23_io_out ? io_r_107_b : _GEN_4826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4828 = 8'h6c == r_count_23_io_out ? io_r_108_b : _GEN_4827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4829 = 8'h6d == r_count_23_io_out ? io_r_109_b : _GEN_4828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4830 = 8'h6e == r_count_23_io_out ? io_r_110_b : _GEN_4829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4831 = 8'h6f == r_count_23_io_out ? io_r_111_b : _GEN_4830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4832 = 8'h70 == r_count_23_io_out ? io_r_112_b : _GEN_4831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4833 = 8'h71 == r_count_23_io_out ? io_r_113_b : _GEN_4832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4834 = 8'h72 == r_count_23_io_out ? io_r_114_b : _GEN_4833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4835 = 8'h73 == r_count_23_io_out ? io_r_115_b : _GEN_4834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4836 = 8'h74 == r_count_23_io_out ? io_r_116_b : _GEN_4835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4837 = 8'h75 == r_count_23_io_out ? io_r_117_b : _GEN_4836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4838 = 8'h76 == r_count_23_io_out ? io_r_118_b : _GEN_4837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4839 = 8'h77 == r_count_23_io_out ? io_r_119_b : _GEN_4838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4840 = 8'h78 == r_count_23_io_out ? io_r_120_b : _GEN_4839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4841 = 8'h79 == r_count_23_io_out ? io_r_121_b : _GEN_4840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4842 = 8'h7a == r_count_23_io_out ? io_r_122_b : _GEN_4841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4843 = 8'h7b == r_count_23_io_out ? io_r_123_b : _GEN_4842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4844 = 8'h7c == r_count_23_io_out ? io_r_124_b : _GEN_4843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4845 = 8'h7d == r_count_23_io_out ? io_r_125_b : _GEN_4844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4846 = 8'h7e == r_count_23_io_out ? io_r_126_b : _GEN_4845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4847 = 8'h7f == r_count_23_io_out ? io_r_127_b : _GEN_4846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4848 = 8'h80 == r_count_23_io_out ? io_r_128_b : _GEN_4847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4849 = 8'h81 == r_count_23_io_out ? io_r_129_b : _GEN_4848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4850 = 8'h82 == r_count_23_io_out ? io_r_130_b : _GEN_4849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4851 = 8'h83 == r_count_23_io_out ? io_r_131_b : _GEN_4850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4852 = 8'h84 == r_count_23_io_out ? io_r_132_b : _GEN_4851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4853 = 8'h85 == r_count_23_io_out ? io_r_133_b : _GEN_4852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4854 = 8'h86 == r_count_23_io_out ? io_r_134_b : _GEN_4853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4855 = 8'h87 == r_count_23_io_out ? io_r_135_b : _GEN_4854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4856 = 8'h88 == r_count_23_io_out ? io_r_136_b : _GEN_4855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4857 = 8'h89 == r_count_23_io_out ? io_r_137_b : _GEN_4856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4858 = 8'h8a == r_count_23_io_out ? io_r_138_b : _GEN_4857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4859 = 8'h8b == r_count_23_io_out ? io_r_139_b : _GEN_4858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4860 = 8'h8c == r_count_23_io_out ? io_r_140_b : _GEN_4859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4861 = 8'h8d == r_count_23_io_out ? io_r_141_b : _GEN_4860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4862 = 8'h8e == r_count_23_io_out ? io_r_142_b : _GEN_4861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4863 = 8'h8f == r_count_23_io_out ? io_r_143_b : _GEN_4862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4864 = 8'h90 == r_count_23_io_out ? io_r_144_b : _GEN_4863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4865 = 8'h91 == r_count_23_io_out ? io_r_145_b : _GEN_4864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4866 = 8'h92 == r_count_23_io_out ? io_r_146_b : _GEN_4865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4867 = 8'h93 == r_count_23_io_out ? io_r_147_b : _GEN_4866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4868 = 8'h94 == r_count_23_io_out ? io_r_148_b : _GEN_4867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4869 = 8'h95 == r_count_23_io_out ? io_r_149_b : _GEN_4868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4870 = 8'h96 == r_count_23_io_out ? io_r_150_b : _GEN_4869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4871 = 8'h97 == r_count_23_io_out ? io_r_151_b : _GEN_4870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4872 = 8'h98 == r_count_23_io_out ? io_r_152_b : _GEN_4871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4873 = 8'h99 == r_count_23_io_out ? io_r_153_b : _GEN_4872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4874 = 8'h9a == r_count_23_io_out ? io_r_154_b : _GEN_4873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4875 = 8'h9b == r_count_23_io_out ? io_r_155_b : _GEN_4874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4876 = 8'h9c == r_count_23_io_out ? io_r_156_b : _GEN_4875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4877 = 8'h9d == r_count_23_io_out ? io_r_157_b : _GEN_4876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4878 = 8'h9e == r_count_23_io_out ? io_r_158_b : _GEN_4877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4879 = 8'h9f == r_count_23_io_out ? io_r_159_b : _GEN_4878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4880 = 8'ha0 == r_count_23_io_out ? io_r_160_b : _GEN_4879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4881 = 8'ha1 == r_count_23_io_out ? io_r_161_b : _GEN_4880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4882 = 8'ha2 == r_count_23_io_out ? io_r_162_b : _GEN_4881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4883 = 8'ha3 == r_count_23_io_out ? io_r_163_b : _GEN_4882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4884 = 8'ha4 == r_count_23_io_out ? io_r_164_b : _GEN_4883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4885 = 8'ha5 == r_count_23_io_out ? io_r_165_b : _GEN_4884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4886 = 8'ha6 == r_count_23_io_out ? io_r_166_b : _GEN_4885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4887 = 8'ha7 == r_count_23_io_out ? io_r_167_b : _GEN_4886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4888 = 8'ha8 == r_count_23_io_out ? io_r_168_b : _GEN_4887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4889 = 8'ha9 == r_count_23_io_out ? io_r_169_b : _GEN_4888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4890 = 8'haa == r_count_23_io_out ? io_r_170_b : _GEN_4889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4891 = 8'hab == r_count_23_io_out ? io_r_171_b : _GEN_4890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4892 = 8'hac == r_count_23_io_out ? io_r_172_b : _GEN_4891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4893 = 8'had == r_count_23_io_out ? io_r_173_b : _GEN_4892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4894 = 8'hae == r_count_23_io_out ? io_r_174_b : _GEN_4893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4895 = 8'haf == r_count_23_io_out ? io_r_175_b : _GEN_4894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4896 = 8'hb0 == r_count_23_io_out ? io_r_176_b : _GEN_4895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4897 = 8'hb1 == r_count_23_io_out ? io_r_177_b : _GEN_4896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4898 = 8'hb2 == r_count_23_io_out ? io_r_178_b : _GEN_4897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4899 = 8'hb3 == r_count_23_io_out ? io_r_179_b : _GEN_4898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4900 = 8'hb4 == r_count_23_io_out ? io_r_180_b : _GEN_4899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4901 = 8'hb5 == r_count_23_io_out ? io_r_181_b : _GEN_4900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4902 = 8'hb6 == r_count_23_io_out ? io_r_182_b : _GEN_4901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4903 = 8'hb7 == r_count_23_io_out ? io_r_183_b : _GEN_4902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4904 = 8'hb8 == r_count_23_io_out ? io_r_184_b : _GEN_4903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4905 = 8'hb9 == r_count_23_io_out ? io_r_185_b : _GEN_4904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4906 = 8'hba == r_count_23_io_out ? io_r_186_b : _GEN_4905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4907 = 8'hbb == r_count_23_io_out ? io_r_187_b : _GEN_4906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4908 = 8'hbc == r_count_23_io_out ? io_r_188_b : _GEN_4907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4909 = 8'hbd == r_count_23_io_out ? io_r_189_b : _GEN_4908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4910 = 8'hbe == r_count_23_io_out ? io_r_190_b : _GEN_4909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4911 = 8'hbf == r_count_23_io_out ? io_r_191_b : _GEN_4910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4912 = 8'hc0 == r_count_23_io_out ? io_r_192_b : _GEN_4911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4913 = 8'hc1 == r_count_23_io_out ? io_r_193_b : _GEN_4912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4914 = 8'hc2 == r_count_23_io_out ? io_r_194_b : _GEN_4913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4915 = 8'hc3 == r_count_23_io_out ? io_r_195_b : _GEN_4914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4916 = 8'hc4 == r_count_23_io_out ? io_r_196_b : _GEN_4915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4917 = 8'hc5 == r_count_23_io_out ? io_r_197_b : _GEN_4916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4918 = 8'hc6 == r_count_23_io_out ? io_r_198_b : _GEN_4917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4921 = 8'h1 == r_count_24_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4922 = 8'h2 == r_count_24_io_out ? io_r_2_b : _GEN_4921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4923 = 8'h3 == r_count_24_io_out ? io_r_3_b : _GEN_4922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4924 = 8'h4 == r_count_24_io_out ? io_r_4_b : _GEN_4923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4925 = 8'h5 == r_count_24_io_out ? io_r_5_b : _GEN_4924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4926 = 8'h6 == r_count_24_io_out ? io_r_6_b : _GEN_4925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4927 = 8'h7 == r_count_24_io_out ? io_r_7_b : _GEN_4926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4928 = 8'h8 == r_count_24_io_out ? io_r_8_b : _GEN_4927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4929 = 8'h9 == r_count_24_io_out ? io_r_9_b : _GEN_4928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4930 = 8'ha == r_count_24_io_out ? io_r_10_b : _GEN_4929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4931 = 8'hb == r_count_24_io_out ? io_r_11_b : _GEN_4930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4932 = 8'hc == r_count_24_io_out ? io_r_12_b : _GEN_4931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4933 = 8'hd == r_count_24_io_out ? io_r_13_b : _GEN_4932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4934 = 8'he == r_count_24_io_out ? io_r_14_b : _GEN_4933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4935 = 8'hf == r_count_24_io_out ? io_r_15_b : _GEN_4934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4936 = 8'h10 == r_count_24_io_out ? io_r_16_b : _GEN_4935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4937 = 8'h11 == r_count_24_io_out ? io_r_17_b : _GEN_4936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4938 = 8'h12 == r_count_24_io_out ? io_r_18_b : _GEN_4937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4939 = 8'h13 == r_count_24_io_out ? io_r_19_b : _GEN_4938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4940 = 8'h14 == r_count_24_io_out ? io_r_20_b : _GEN_4939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4941 = 8'h15 == r_count_24_io_out ? io_r_21_b : _GEN_4940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4942 = 8'h16 == r_count_24_io_out ? io_r_22_b : _GEN_4941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4943 = 8'h17 == r_count_24_io_out ? io_r_23_b : _GEN_4942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4944 = 8'h18 == r_count_24_io_out ? io_r_24_b : _GEN_4943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4945 = 8'h19 == r_count_24_io_out ? io_r_25_b : _GEN_4944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4946 = 8'h1a == r_count_24_io_out ? io_r_26_b : _GEN_4945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4947 = 8'h1b == r_count_24_io_out ? io_r_27_b : _GEN_4946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4948 = 8'h1c == r_count_24_io_out ? io_r_28_b : _GEN_4947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4949 = 8'h1d == r_count_24_io_out ? io_r_29_b : _GEN_4948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4950 = 8'h1e == r_count_24_io_out ? io_r_30_b : _GEN_4949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4951 = 8'h1f == r_count_24_io_out ? io_r_31_b : _GEN_4950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4952 = 8'h20 == r_count_24_io_out ? io_r_32_b : _GEN_4951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4953 = 8'h21 == r_count_24_io_out ? io_r_33_b : _GEN_4952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4954 = 8'h22 == r_count_24_io_out ? io_r_34_b : _GEN_4953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4955 = 8'h23 == r_count_24_io_out ? io_r_35_b : _GEN_4954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4956 = 8'h24 == r_count_24_io_out ? io_r_36_b : _GEN_4955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4957 = 8'h25 == r_count_24_io_out ? io_r_37_b : _GEN_4956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4958 = 8'h26 == r_count_24_io_out ? io_r_38_b : _GEN_4957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4959 = 8'h27 == r_count_24_io_out ? io_r_39_b : _GEN_4958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4960 = 8'h28 == r_count_24_io_out ? io_r_40_b : _GEN_4959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4961 = 8'h29 == r_count_24_io_out ? io_r_41_b : _GEN_4960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4962 = 8'h2a == r_count_24_io_out ? io_r_42_b : _GEN_4961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4963 = 8'h2b == r_count_24_io_out ? io_r_43_b : _GEN_4962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4964 = 8'h2c == r_count_24_io_out ? io_r_44_b : _GEN_4963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4965 = 8'h2d == r_count_24_io_out ? io_r_45_b : _GEN_4964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4966 = 8'h2e == r_count_24_io_out ? io_r_46_b : _GEN_4965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4967 = 8'h2f == r_count_24_io_out ? io_r_47_b : _GEN_4966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4968 = 8'h30 == r_count_24_io_out ? io_r_48_b : _GEN_4967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4969 = 8'h31 == r_count_24_io_out ? io_r_49_b : _GEN_4968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4970 = 8'h32 == r_count_24_io_out ? io_r_50_b : _GEN_4969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4971 = 8'h33 == r_count_24_io_out ? io_r_51_b : _GEN_4970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4972 = 8'h34 == r_count_24_io_out ? io_r_52_b : _GEN_4971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4973 = 8'h35 == r_count_24_io_out ? io_r_53_b : _GEN_4972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4974 = 8'h36 == r_count_24_io_out ? io_r_54_b : _GEN_4973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4975 = 8'h37 == r_count_24_io_out ? io_r_55_b : _GEN_4974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4976 = 8'h38 == r_count_24_io_out ? io_r_56_b : _GEN_4975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4977 = 8'h39 == r_count_24_io_out ? io_r_57_b : _GEN_4976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4978 = 8'h3a == r_count_24_io_out ? io_r_58_b : _GEN_4977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4979 = 8'h3b == r_count_24_io_out ? io_r_59_b : _GEN_4978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4980 = 8'h3c == r_count_24_io_out ? io_r_60_b : _GEN_4979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4981 = 8'h3d == r_count_24_io_out ? io_r_61_b : _GEN_4980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4982 = 8'h3e == r_count_24_io_out ? io_r_62_b : _GEN_4981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4983 = 8'h3f == r_count_24_io_out ? io_r_63_b : _GEN_4982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4984 = 8'h40 == r_count_24_io_out ? io_r_64_b : _GEN_4983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4985 = 8'h41 == r_count_24_io_out ? io_r_65_b : _GEN_4984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4986 = 8'h42 == r_count_24_io_out ? io_r_66_b : _GEN_4985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4987 = 8'h43 == r_count_24_io_out ? io_r_67_b : _GEN_4986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4988 = 8'h44 == r_count_24_io_out ? io_r_68_b : _GEN_4987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4989 = 8'h45 == r_count_24_io_out ? io_r_69_b : _GEN_4988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4990 = 8'h46 == r_count_24_io_out ? io_r_70_b : _GEN_4989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4991 = 8'h47 == r_count_24_io_out ? io_r_71_b : _GEN_4990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4992 = 8'h48 == r_count_24_io_out ? io_r_72_b : _GEN_4991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4993 = 8'h49 == r_count_24_io_out ? io_r_73_b : _GEN_4992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4994 = 8'h4a == r_count_24_io_out ? io_r_74_b : _GEN_4993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4995 = 8'h4b == r_count_24_io_out ? io_r_75_b : _GEN_4994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4996 = 8'h4c == r_count_24_io_out ? io_r_76_b : _GEN_4995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4997 = 8'h4d == r_count_24_io_out ? io_r_77_b : _GEN_4996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4998 = 8'h4e == r_count_24_io_out ? io_r_78_b : _GEN_4997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4999 = 8'h4f == r_count_24_io_out ? io_r_79_b : _GEN_4998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5000 = 8'h50 == r_count_24_io_out ? io_r_80_b : _GEN_4999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5001 = 8'h51 == r_count_24_io_out ? io_r_81_b : _GEN_5000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5002 = 8'h52 == r_count_24_io_out ? io_r_82_b : _GEN_5001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5003 = 8'h53 == r_count_24_io_out ? io_r_83_b : _GEN_5002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5004 = 8'h54 == r_count_24_io_out ? io_r_84_b : _GEN_5003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5005 = 8'h55 == r_count_24_io_out ? io_r_85_b : _GEN_5004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5006 = 8'h56 == r_count_24_io_out ? io_r_86_b : _GEN_5005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5007 = 8'h57 == r_count_24_io_out ? io_r_87_b : _GEN_5006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5008 = 8'h58 == r_count_24_io_out ? io_r_88_b : _GEN_5007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5009 = 8'h59 == r_count_24_io_out ? io_r_89_b : _GEN_5008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5010 = 8'h5a == r_count_24_io_out ? io_r_90_b : _GEN_5009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5011 = 8'h5b == r_count_24_io_out ? io_r_91_b : _GEN_5010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5012 = 8'h5c == r_count_24_io_out ? io_r_92_b : _GEN_5011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5013 = 8'h5d == r_count_24_io_out ? io_r_93_b : _GEN_5012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5014 = 8'h5e == r_count_24_io_out ? io_r_94_b : _GEN_5013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5015 = 8'h5f == r_count_24_io_out ? io_r_95_b : _GEN_5014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5016 = 8'h60 == r_count_24_io_out ? io_r_96_b : _GEN_5015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5017 = 8'h61 == r_count_24_io_out ? io_r_97_b : _GEN_5016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5018 = 8'h62 == r_count_24_io_out ? io_r_98_b : _GEN_5017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5019 = 8'h63 == r_count_24_io_out ? io_r_99_b : _GEN_5018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5020 = 8'h64 == r_count_24_io_out ? io_r_100_b : _GEN_5019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5021 = 8'h65 == r_count_24_io_out ? io_r_101_b : _GEN_5020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5022 = 8'h66 == r_count_24_io_out ? io_r_102_b : _GEN_5021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5023 = 8'h67 == r_count_24_io_out ? io_r_103_b : _GEN_5022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5024 = 8'h68 == r_count_24_io_out ? io_r_104_b : _GEN_5023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5025 = 8'h69 == r_count_24_io_out ? io_r_105_b : _GEN_5024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5026 = 8'h6a == r_count_24_io_out ? io_r_106_b : _GEN_5025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5027 = 8'h6b == r_count_24_io_out ? io_r_107_b : _GEN_5026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5028 = 8'h6c == r_count_24_io_out ? io_r_108_b : _GEN_5027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5029 = 8'h6d == r_count_24_io_out ? io_r_109_b : _GEN_5028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5030 = 8'h6e == r_count_24_io_out ? io_r_110_b : _GEN_5029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5031 = 8'h6f == r_count_24_io_out ? io_r_111_b : _GEN_5030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5032 = 8'h70 == r_count_24_io_out ? io_r_112_b : _GEN_5031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5033 = 8'h71 == r_count_24_io_out ? io_r_113_b : _GEN_5032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5034 = 8'h72 == r_count_24_io_out ? io_r_114_b : _GEN_5033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5035 = 8'h73 == r_count_24_io_out ? io_r_115_b : _GEN_5034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5036 = 8'h74 == r_count_24_io_out ? io_r_116_b : _GEN_5035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5037 = 8'h75 == r_count_24_io_out ? io_r_117_b : _GEN_5036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5038 = 8'h76 == r_count_24_io_out ? io_r_118_b : _GEN_5037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5039 = 8'h77 == r_count_24_io_out ? io_r_119_b : _GEN_5038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5040 = 8'h78 == r_count_24_io_out ? io_r_120_b : _GEN_5039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5041 = 8'h79 == r_count_24_io_out ? io_r_121_b : _GEN_5040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5042 = 8'h7a == r_count_24_io_out ? io_r_122_b : _GEN_5041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5043 = 8'h7b == r_count_24_io_out ? io_r_123_b : _GEN_5042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5044 = 8'h7c == r_count_24_io_out ? io_r_124_b : _GEN_5043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5045 = 8'h7d == r_count_24_io_out ? io_r_125_b : _GEN_5044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5046 = 8'h7e == r_count_24_io_out ? io_r_126_b : _GEN_5045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5047 = 8'h7f == r_count_24_io_out ? io_r_127_b : _GEN_5046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5048 = 8'h80 == r_count_24_io_out ? io_r_128_b : _GEN_5047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5049 = 8'h81 == r_count_24_io_out ? io_r_129_b : _GEN_5048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5050 = 8'h82 == r_count_24_io_out ? io_r_130_b : _GEN_5049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5051 = 8'h83 == r_count_24_io_out ? io_r_131_b : _GEN_5050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5052 = 8'h84 == r_count_24_io_out ? io_r_132_b : _GEN_5051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5053 = 8'h85 == r_count_24_io_out ? io_r_133_b : _GEN_5052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5054 = 8'h86 == r_count_24_io_out ? io_r_134_b : _GEN_5053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5055 = 8'h87 == r_count_24_io_out ? io_r_135_b : _GEN_5054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5056 = 8'h88 == r_count_24_io_out ? io_r_136_b : _GEN_5055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5057 = 8'h89 == r_count_24_io_out ? io_r_137_b : _GEN_5056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5058 = 8'h8a == r_count_24_io_out ? io_r_138_b : _GEN_5057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5059 = 8'h8b == r_count_24_io_out ? io_r_139_b : _GEN_5058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5060 = 8'h8c == r_count_24_io_out ? io_r_140_b : _GEN_5059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5061 = 8'h8d == r_count_24_io_out ? io_r_141_b : _GEN_5060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5062 = 8'h8e == r_count_24_io_out ? io_r_142_b : _GEN_5061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5063 = 8'h8f == r_count_24_io_out ? io_r_143_b : _GEN_5062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5064 = 8'h90 == r_count_24_io_out ? io_r_144_b : _GEN_5063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5065 = 8'h91 == r_count_24_io_out ? io_r_145_b : _GEN_5064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5066 = 8'h92 == r_count_24_io_out ? io_r_146_b : _GEN_5065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5067 = 8'h93 == r_count_24_io_out ? io_r_147_b : _GEN_5066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5068 = 8'h94 == r_count_24_io_out ? io_r_148_b : _GEN_5067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5069 = 8'h95 == r_count_24_io_out ? io_r_149_b : _GEN_5068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5070 = 8'h96 == r_count_24_io_out ? io_r_150_b : _GEN_5069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5071 = 8'h97 == r_count_24_io_out ? io_r_151_b : _GEN_5070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5072 = 8'h98 == r_count_24_io_out ? io_r_152_b : _GEN_5071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5073 = 8'h99 == r_count_24_io_out ? io_r_153_b : _GEN_5072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5074 = 8'h9a == r_count_24_io_out ? io_r_154_b : _GEN_5073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5075 = 8'h9b == r_count_24_io_out ? io_r_155_b : _GEN_5074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5076 = 8'h9c == r_count_24_io_out ? io_r_156_b : _GEN_5075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5077 = 8'h9d == r_count_24_io_out ? io_r_157_b : _GEN_5076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5078 = 8'h9e == r_count_24_io_out ? io_r_158_b : _GEN_5077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5079 = 8'h9f == r_count_24_io_out ? io_r_159_b : _GEN_5078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5080 = 8'ha0 == r_count_24_io_out ? io_r_160_b : _GEN_5079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5081 = 8'ha1 == r_count_24_io_out ? io_r_161_b : _GEN_5080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5082 = 8'ha2 == r_count_24_io_out ? io_r_162_b : _GEN_5081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5083 = 8'ha3 == r_count_24_io_out ? io_r_163_b : _GEN_5082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5084 = 8'ha4 == r_count_24_io_out ? io_r_164_b : _GEN_5083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5085 = 8'ha5 == r_count_24_io_out ? io_r_165_b : _GEN_5084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5086 = 8'ha6 == r_count_24_io_out ? io_r_166_b : _GEN_5085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5087 = 8'ha7 == r_count_24_io_out ? io_r_167_b : _GEN_5086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5088 = 8'ha8 == r_count_24_io_out ? io_r_168_b : _GEN_5087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5089 = 8'ha9 == r_count_24_io_out ? io_r_169_b : _GEN_5088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5090 = 8'haa == r_count_24_io_out ? io_r_170_b : _GEN_5089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5091 = 8'hab == r_count_24_io_out ? io_r_171_b : _GEN_5090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5092 = 8'hac == r_count_24_io_out ? io_r_172_b : _GEN_5091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5093 = 8'had == r_count_24_io_out ? io_r_173_b : _GEN_5092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5094 = 8'hae == r_count_24_io_out ? io_r_174_b : _GEN_5093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5095 = 8'haf == r_count_24_io_out ? io_r_175_b : _GEN_5094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5096 = 8'hb0 == r_count_24_io_out ? io_r_176_b : _GEN_5095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5097 = 8'hb1 == r_count_24_io_out ? io_r_177_b : _GEN_5096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5098 = 8'hb2 == r_count_24_io_out ? io_r_178_b : _GEN_5097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5099 = 8'hb3 == r_count_24_io_out ? io_r_179_b : _GEN_5098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5100 = 8'hb4 == r_count_24_io_out ? io_r_180_b : _GEN_5099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5101 = 8'hb5 == r_count_24_io_out ? io_r_181_b : _GEN_5100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5102 = 8'hb6 == r_count_24_io_out ? io_r_182_b : _GEN_5101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5103 = 8'hb7 == r_count_24_io_out ? io_r_183_b : _GEN_5102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5104 = 8'hb8 == r_count_24_io_out ? io_r_184_b : _GEN_5103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5105 = 8'hb9 == r_count_24_io_out ? io_r_185_b : _GEN_5104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5106 = 8'hba == r_count_24_io_out ? io_r_186_b : _GEN_5105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5107 = 8'hbb == r_count_24_io_out ? io_r_187_b : _GEN_5106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5108 = 8'hbc == r_count_24_io_out ? io_r_188_b : _GEN_5107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5109 = 8'hbd == r_count_24_io_out ? io_r_189_b : _GEN_5108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5110 = 8'hbe == r_count_24_io_out ? io_r_190_b : _GEN_5109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5111 = 8'hbf == r_count_24_io_out ? io_r_191_b : _GEN_5110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5112 = 8'hc0 == r_count_24_io_out ? io_r_192_b : _GEN_5111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5113 = 8'hc1 == r_count_24_io_out ? io_r_193_b : _GEN_5112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5114 = 8'hc2 == r_count_24_io_out ? io_r_194_b : _GEN_5113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5115 = 8'hc3 == r_count_24_io_out ? io_r_195_b : _GEN_5114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5116 = 8'hc4 == r_count_24_io_out ? io_r_196_b : _GEN_5115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5117 = 8'hc5 == r_count_24_io_out ? io_r_197_b : _GEN_5116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5118 = 8'hc6 == r_count_24_io_out ? io_r_198_b : _GEN_5117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5121 = 8'h1 == r_count_25_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5122 = 8'h2 == r_count_25_io_out ? io_r_2_b : _GEN_5121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5123 = 8'h3 == r_count_25_io_out ? io_r_3_b : _GEN_5122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5124 = 8'h4 == r_count_25_io_out ? io_r_4_b : _GEN_5123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5125 = 8'h5 == r_count_25_io_out ? io_r_5_b : _GEN_5124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5126 = 8'h6 == r_count_25_io_out ? io_r_6_b : _GEN_5125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5127 = 8'h7 == r_count_25_io_out ? io_r_7_b : _GEN_5126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5128 = 8'h8 == r_count_25_io_out ? io_r_8_b : _GEN_5127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5129 = 8'h9 == r_count_25_io_out ? io_r_9_b : _GEN_5128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5130 = 8'ha == r_count_25_io_out ? io_r_10_b : _GEN_5129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5131 = 8'hb == r_count_25_io_out ? io_r_11_b : _GEN_5130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5132 = 8'hc == r_count_25_io_out ? io_r_12_b : _GEN_5131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5133 = 8'hd == r_count_25_io_out ? io_r_13_b : _GEN_5132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5134 = 8'he == r_count_25_io_out ? io_r_14_b : _GEN_5133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5135 = 8'hf == r_count_25_io_out ? io_r_15_b : _GEN_5134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5136 = 8'h10 == r_count_25_io_out ? io_r_16_b : _GEN_5135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5137 = 8'h11 == r_count_25_io_out ? io_r_17_b : _GEN_5136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5138 = 8'h12 == r_count_25_io_out ? io_r_18_b : _GEN_5137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5139 = 8'h13 == r_count_25_io_out ? io_r_19_b : _GEN_5138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5140 = 8'h14 == r_count_25_io_out ? io_r_20_b : _GEN_5139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5141 = 8'h15 == r_count_25_io_out ? io_r_21_b : _GEN_5140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5142 = 8'h16 == r_count_25_io_out ? io_r_22_b : _GEN_5141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5143 = 8'h17 == r_count_25_io_out ? io_r_23_b : _GEN_5142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5144 = 8'h18 == r_count_25_io_out ? io_r_24_b : _GEN_5143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5145 = 8'h19 == r_count_25_io_out ? io_r_25_b : _GEN_5144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5146 = 8'h1a == r_count_25_io_out ? io_r_26_b : _GEN_5145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5147 = 8'h1b == r_count_25_io_out ? io_r_27_b : _GEN_5146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5148 = 8'h1c == r_count_25_io_out ? io_r_28_b : _GEN_5147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5149 = 8'h1d == r_count_25_io_out ? io_r_29_b : _GEN_5148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5150 = 8'h1e == r_count_25_io_out ? io_r_30_b : _GEN_5149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5151 = 8'h1f == r_count_25_io_out ? io_r_31_b : _GEN_5150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5152 = 8'h20 == r_count_25_io_out ? io_r_32_b : _GEN_5151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5153 = 8'h21 == r_count_25_io_out ? io_r_33_b : _GEN_5152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5154 = 8'h22 == r_count_25_io_out ? io_r_34_b : _GEN_5153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5155 = 8'h23 == r_count_25_io_out ? io_r_35_b : _GEN_5154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5156 = 8'h24 == r_count_25_io_out ? io_r_36_b : _GEN_5155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5157 = 8'h25 == r_count_25_io_out ? io_r_37_b : _GEN_5156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5158 = 8'h26 == r_count_25_io_out ? io_r_38_b : _GEN_5157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5159 = 8'h27 == r_count_25_io_out ? io_r_39_b : _GEN_5158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5160 = 8'h28 == r_count_25_io_out ? io_r_40_b : _GEN_5159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5161 = 8'h29 == r_count_25_io_out ? io_r_41_b : _GEN_5160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5162 = 8'h2a == r_count_25_io_out ? io_r_42_b : _GEN_5161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5163 = 8'h2b == r_count_25_io_out ? io_r_43_b : _GEN_5162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5164 = 8'h2c == r_count_25_io_out ? io_r_44_b : _GEN_5163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5165 = 8'h2d == r_count_25_io_out ? io_r_45_b : _GEN_5164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5166 = 8'h2e == r_count_25_io_out ? io_r_46_b : _GEN_5165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5167 = 8'h2f == r_count_25_io_out ? io_r_47_b : _GEN_5166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5168 = 8'h30 == r_count_25_io_out ? io_r_48_b : _GEN_5167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5169 = 8'h31 == r_count_25_io_out ? io_r_49_b : _GEN_5168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5170 = 8'h32 == r_count_25_io_out ? io_r_50_b : _GEN_5169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5171 = 8'h33 == r_count_25_io_out ? io_r_51_b : _GEN_5170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5172 = 8'h34 == r_count_25_io_out ? io_r_52_b : _GEN_5171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5173 = 8'h35 == r_count_25_io_out ? io_r_53_b : _GEN_5172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5174 = 8'h36 == r_count_25_io_out ? io_r_54_b : _GEN_5173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5175 = 8'h37 == r_count_25_io_out ? io_r_55_b : _GEN_5174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5176 = 8'h38 == r_count_25_io_out ? io_r_56_b : _GEN_5175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5177 = 8'h39 == r_count_25_io_out ? io_r_57_b : _GEN_5176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5178 = 8'h3a == r_count_25_io_out ? io_r_58_b : _GEN_5177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5179 = 8'h3b == r_count_25_io_out ? io_r_59_b : _GEN_5178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5180 = 8'h3c == r_count_25_io_out ? io_r_60_b : _GEN_5179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5181 = 8'h3d == r_count_25_io_out ? io_r_61_b : _GEN_5180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5182 = 8'h3e == r_count_25_io_out ? io_r_62_b : _GEN_5181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5183 = 8'h3f == r_count_25_io_out ? io_r_63_b : _GEN_5182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5184 = 8'h40 == r_count_25_io_out ? io_r_64_b : _GEN_5183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5185 = 8'h41 == r_count_25_io_out ? io_r_65_b : _GEN_5184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5186 = 8'h42 == r_count_25_io_out ? io_r_66_b : _GEN_5185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5187 = 8'h43 == r_count_25_io_out ? io_r_67_b : _GEN_5186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5188 = 8'h44 == r_count_25_io_out ? io_r_68_b : _GEN_5187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5189 = 8'h45 == r_count_25_io_out ? io_r_69_b : _GEN_5188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5190 = 8'h46 == r_count_25_io_out ? io_r_70_b : _GEN_5189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5191 = 8'h47 == r_count_25_io_out ? io_r_71_b : _GEN_5190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5192 = 8'h48 == r_count_25_io_out ? io_r_72_b : _GEN_5191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5193 = 8'h49 == r_count_25_io_out ? io_r_73_b : _GEN_5192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5194 = 8'h4a == r_count_25_io_out ? io_r_74_b : _GEN_5193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5195 = 8'h4b == r_count_25_io_out ? io_r_75_b : _GEN_5194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5196 = 8'h4c == r_count_25_io_out ? io_r_76_b : _GEN_5195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5197 = 8'h4d == r_count_25_io_out ? io_r_77_b : _GEN_5196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5198 = 8'h4e == r_count_25_io_out ? io_r_78_b : _GEN_5197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5199 = 8'h4f == r_count_25_io_out ? io_r_79_b : _GEN_5198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5200 = 8'h50 == r_count_25_io_out ? io_r_80_b : _GEN_5199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5201 = 8'h51 == r_count_25_io_out ? io_r_81_b : _GEN_5200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5202 = 8'h52 == r_count_25_io_out ? io_r_82_b : _GEN_5201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5203 = 8'h53 == r_count_25_io_out ? io_r_83_b : _GEN_5202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5204 = 8'h54 == r_count_25_io_out ? io_r_84_b : _GEN_5203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5205 = 8'h55 == r_count_25_io_out ? io_r_85_b : _GEN_5204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5206 = 8'h56 == r_count_25_io_out ? io_r_86_b : _GEN_5205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5207 = 8'h57 == r_count_25_io_out ? io_r_87_b : _GEN_5206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5208 = 8'h58 == r_count_25_io_out ? io_r_88_b : _GEN_5207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5209 = 8'h59 == r_count_25_io_out ? io_r_89_b : _GEN_5208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5210 = 8'h5a == r_count_25_io_out ? io_r_90_b : _GEN_5209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5211 = 8'h5b == r_count_25_io_out ? io_r_91_b : _GEN_5210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5212 = 8'h5c == r_count_25_io_out ? io_r_92_b : _GEN_5211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5213 = 8'h5d == r_count_25_io_out ? io_r_93_b : _GEN_5212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5214 = 8'h5e == r_count_25_io_out ? io_r_94_b : _GEN_5213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5215 = 8'h5f == r_count_25_io_out ? io_r_95_b : _GEN_5214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5216 = 8'h60 == r_count_25_io_out ? io_r_96_b : _GEN_5215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5217 = 8'h61 == r_count_25_io_out ? io_r_97_b : _GEN_5216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5218 = 8'h62 == r_count_25_io_out ? io_r_98_b : _GEN_5217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5219 = 8'h63 == r_count_25_io_out ? io_r_99_b : _GEN_5218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5220 = 8'h64 == r_count_25_io_out ? io_r_100_b : _GEN_5219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5221 = 8'h65 == r_count_25_io_out ? io_r_101_b : _GEN_5220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5222 = 8'h66 == r_count_25_io_out ? io_r_102_b : _GEN_5221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5223 = 8'h67 == r_count_25_io_out ? io_r_103_b : _GEN_5222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5224 = 8'h68 == r_count_25_io_out ? io_r_104_b : _GEN_5223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5225 = 8'h69 == r_count_25_io_out ? io_r_105_b : _GEN_5224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5226 = 8'h6a == r_count_25_io_out ? io_r_106_b : _GEN_5225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5227 = 8'h6b == r_count_25_io_out ? io_r_107_b : _GEN_5226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5228 = 8'h6c == r_count_25_io_out ? io_r_108_b : _GEN_5227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5229 = 8'h6d == r_count_25_io_out ? io_r_109_b : _GEN_5228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5230 = 8'h6e == r_count_25_io_out ? io_r_110_b : _GEN_5229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5231 = 8'h6f == r_count_25_io_out ? io_r_111_b : _GEN_5230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5232 = 8'h70 == r_count_25_io_out ? io_r_112_b : _GEN_5231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5233 = 8'h71 == r_count_25_io_out ? io_r_113_b : _GEN_5232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5234 = 8'h72 == r_count_25_io_out ? io_r_114_b : _GEN_5233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5235 = 8'h73 == r_count_25_io_out ? io_r_115_b : _GEN_5234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5236 = 8'h74 == r_count_25_io_out ? io_r_116_b : _GEN_5235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5237 = 8'h75 == r_count_25_io_out ? io_r_117_b : _GEN_5236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5238 = 8'h76 == r_count_25_io_out ? io_r_118_b : _GEN_5237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5239 = 8'h77 == r_count_25_io_out ? io_r_119_b : _GEN_5238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5240 = 8'h78 == r_count_25_io_out ? io_r_120_b : _GEN_5239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5241 = 8'h79 == r_count_25_io_out ? io_r_121_b : _GEN_5240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5242 = 8'h7a == r_count_25_io_out ? io_r_122_b : _GEN_5241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5243 = 8'h7b == r_count_25_io_out ? io_r_123_b : _GEN_5242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5244 = 8'h7c == r_count_25_io_out ? io_r_124_b : _GEN_5243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5245 = 8'h7d == r_count_25_io_out ? io_r_125_b : _GEN_5244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5246 = 8'h7e == r_count_25_io_out ? io_r_126_b : _GEN_5245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5247 = 8'h7f == r_count_25_io_out ? io_r_127_b : _GEN_5246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5248 = 8'h80 == r_count_25_io_out ? io_r_128_b : _GEN_5247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5249 = 8'h81 == r_count_25_io_out ? io_r_129_b : _GEN_5248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5250 = 8'h82 == r_count_25_io_out ? io_r_130_b : _GEN_5249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5251 = 8'h83 == r_count_25_io_out ? io_r_131_b : _GEN_5250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5252 = 8'h84 == r_count_25_io_out ? io_r_132_b : _GEN_5251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5253 = 8'h85 == r_count_25_io_out ? io_r_133_b : _GEN_5252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5254 = 8'h86 == r_count_25_io_out ? io_r_134_b : _GEN_5253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5255 = 8'h87 == r_count_25_io_out ? io_r_135_b : _GEN_5254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5256 = 8'h88 == r_count_25_io_out ? io_r_136_b : _GEN_5255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5257 = 8'h89 == r_count_25_io_out ? io_r_137_b : _GEN_5256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5258 = 8'h8a == r_count_25_io_out ? io_r_138_b : _GEN_5257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5259 = 8'h8b == r_count_25_io_out ? io_r_139_b : _GEN_5258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5260 = 8'h8c == r_count_25_io_out ? io_r_140_b : _GEN_5259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5261 = 8'h8d == r_count_25_io_out ? io_r_141_b : _GEN_5260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5262 = 8'h8e == r_count_25_io_out ? io_r_142_b : _GEN_5261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5263 = 8'h8f == r_count_25_io_out ? io_r_143_b : _GEN_5262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5264 = 8'h90 == r_count_25_io_out ? io_r_144_b : _GEN_5263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5265 = 8'h91 == r_count_25_io_out ? io_r_145_b : _GEN_5264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5266 = 8'h92 == r_count_25_io_out ? io_r_146_b : _GEN_5265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5267 = 8'h93 == r_count_25_io_out ? io_r_147_b : _GEN_5266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5268 = 8'h94 == r_count_25_io_out ? io_r_148_b : _GEN_5267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5269 = 8'h95 == r_count_25_io_out ? io_r_149_b : _GEN_5268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5270 = 8'h96 == r_count_25_io_out ? io_r_150_b : _GEN_5269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5271 = 8'h97 == r_count_25_io_out ? io_r_151_b : _GEN_5270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5272 = 8'h98 == r_count_25_io_out ? io_r_152_b : _GEN_5271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5273 = 8'h99 == r_count_25_io_out ? io_r_153_b : _GEN_5272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5274 = 8'h9a == r_count_25_io_out ? io_r_154_b : _GEN_5273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5275 = 8'h9b == r_count_25_io_out ? io_r_155_b : _GEN_5274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5276 = 8'h9c == r_count_25_io_out ? io_r_156_b : _GEN_5275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5277 = 8'h9d == r_count_25_io_out ? io_r_157_b : _GEN_5276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5278 = 8'h9e == r_count_25_io_out ? io_r_158_b : _GEN_5277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5279 = 8'h9f == r_count_25_io_out ? io_r_159_b : _GEN_5278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5280 = 8'ha0 == r_count_25_io_out ? io_r_160_b : _GEN_5279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5281 = 8'ha1 == r_count_25_io_out ? io_r_161_b : _GEN_5280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5282 = 8'ha2 == r_count_25_io_out ? io_r_162_b : _GEN_5281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5283 = 8'ha3 == r_count_25_io_out ? io_r_163_b : _GEN_5282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5284 = 8'ha4 == r_count_25_io_out ? io_r_164_b : _GEN_5283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5285 = 8'ha5 == r_count_25_io_out ? io_r_165_b : _GEN_5284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5286 = 8'ha6 == r_count_25_io_out ? io_r_166_b : _GEN_5285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5287 = 8'ha7 == r_count_25_io_out ? io_r_167_b : _GEN_5286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5288 = 8'ha8 == r_count_25_io_out ? io_r_168_b : _GEN_5287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5289 = 8'ha9 == r_count_25_io_out ? io_r_169_b : _GEN_5288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5290 = 8'haa == r_count_25_io_out ? io_r_170_b : _GEN_5289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5291 = 8'hab == r_count_25_io_out ? io_r_171_b : _GEN_5290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5292 = 8'hac == r_count_25_io_out ? io_r_172_b : _GEN_5291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5293 = 8'had == r_count_25_io_out ? io_r_173_b : _GEN_5292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5294 = 8'hae == r_count_25_io_out ? io_r_174_b : _GEN_5293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5295 = 8'haf == r_count_25_io_out ? io_r_175_b : _GEN_5294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5296 = 8'hb0 == r_count_25_io_out ? io_r_176_b : _GEN_5295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5297 = 8'hb1 == r_count_25_io_out ? io_r_177_b : _GEN_5296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5298 = 8'hb2 == r_count_25_io_out ? io_r_178_b : _GEN_5297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5299 = 8'hb3 == r_count_25_io_out ? io_r_179_b : _GEN_5298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5300 = 8'hb4 == r_count_25_io_out ? io_r_180_b : _GEN_5299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5301 = 8'hb5 == r_count_25_io_out ? io_r_181_b : _GEN_5300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5302 = 8'hb6 == r_count_25_io_out ? io_r_182_b : _GEN_5301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5303 = 8'hb7 == r_count_25_io_out ? io_r_183_b : _GEN_5302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5304 = 8'hb8 == r_count_25_io_out ? io_r_184_b : _GEN_5303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5305 = 8'hb9 == r_count_25_io_out ? io_r_185_b : _GEN_5304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5306 = 8'hba == r_count_25_io_out ? io_r_186_b : _GEN_5305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5307 = 8'hbb == r_count_25_io_out ? io_r_187_b : _GEN_5306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5308 = 8'hbc == r_count_25_io_out ? io_r_188_b : _GEN_5307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5309 = 8'hbd == r_count_25_io_out ? io_r_189_b : _GEN_5308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5310 = 8'hbe == r_count_25_io_out ? io_r_190_b : _GEN_5309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5311 = 8'hbf == r_count_25_io_out ? io_r_191_b : _GEN_5310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5312 = 8'hc0 == r_count_25_io_out ? io_r_192_b : _GEN_5311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5313 = 8'hc1 == r_count_25_io_out ? io_r_193_b : _GEN_5312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5314 = 8'hc2 == r_count_25_io_out ? io_r_194_b : _GEN_5313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5315 = 8'hc3 == r_count_25_io_out ? io_r_195_b : _GEN_5314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5316 = 8'hc4 == r_count_25_io_out ? io_r_196_b : _GEN_5315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5317 = 8'hc5 == r_count_25_io_out ? io_r_197_b : _GEN_5316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5318 = 8'hc6 == r_count_25_io_out ? io_r_198_b : _GEN_5317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5321 = 8'h1 == r_count_26_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5322 = 8'h2 == r_count_26_io_out ? io_r_2_b : _GEN_5321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5323 = 8'h3 == r_count_26_io_out ? io_r_3_b : _GEN_5322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5324 = 8'h4 == r_count_26_io_out ? io_r_4_b : _GEN_5323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5325 = 8'h5 == r_count_26_io_out ? io_r_5_b : _GEN_5324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5326 = 8'h6 == r_count_26_io_out ? io_r_6_b : _GEN_5325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5327 = 8'h7 == r_count_26_io_out ? io_r_7_b : _GEN_5326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5328 = 8'h8 == r_count_26_io_out ? io_r_8_b : _GEN_5327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5329 = 8'h9 == r_count_26_io_out ? io_r_9_b : _GEN_5328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5330 = 8'ha == r_count_26_io_out ? io_r_10_b : _GEN_5329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5331 = 8'hb == r_count_26_io_out ? io_r_11_b : _GEN_5330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5332 = 8'hc == r_count_26_io_out ? io_r_12_b : _GEN_5331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5333 = 8'hd == r_count_26_io_out ? io_r_13_b : _GEN_5332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5334 = 8'he == r_count_26_io_out ? io_r_14_b : _GEN_5333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5335 = 8'hf == r_count_26_io_out ? io_r_15_b : _GEN_5334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5336 = 8'h10 == r_count_26_io_out ? io_r_16_b : _GEN_5335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5337 = 8'h11 == r_count_26_io_out ? io_r_17_b : _GEN_5336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5338 = 8'h12 == r_count_26_io_out ? io_r_18_b : _GEN_5337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5339 = 8'h13 == r_count_26_io_out ? io_r_19_b : _GEN_5338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5340 = 8'h14 == r_count_26_io_out ? io_r_20_b : _GEN_5339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5341 = 8'h15 == r_count_26_io_out ? io_r_21_b : _GEN_5340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5342 = 8'h16 == r_count_26_io_out ? io_r_22_b : _GEN_5341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5343 = 8'h17 == r_count_26_io_out ? io_r_23_b : _GEN_5342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5344 = 8'h18 == r_count_26_io_out ? io_r_24_b : _GEN_5343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5345 = 8'h19 == r_count_26_io_out ? io_r_25_b : _GEN_5344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5346 = 8'h1a == r_count_26_io_out ? io_r_26_b : _GEN_5345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5347 = 8'h1b == r_count_26_io_out ? io_r_27_b : _GEN_5346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5348 = 8'h1c == r_count_26_io_out ? io_r_28_b : _GEN_5347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5349 = 8'h1d == r_count_26_io_out ? io_r_29_b : _GEN_5348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5350 = 8'h1e == r_count_26_io_out ? io_r_30_b : _GEN_5349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5351 = 8'h1f == r_count_26_io_out ? io_r_31_b : _GEN_5350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5352 = 8'h20 == r_count_26_io_out ? io_r_32_b : _GEN_5351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5353 = 8'h21 == r_count_26_io_out ? io_r_33_b : _GEN_5352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5354 = 8'h22 == r_count_26_io_out ? io_r_34_b : _GEN_5353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5355 = 8'h23 == r_count_26_io_out ? io_r_35_b : _GEN_5354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5356 = 8'h24 == r_count_26_io_out ? io_r_36_b : _GEN_5355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5357 = 8'h25 == r_count_26_io_out ? io_r_37_b : _GEN_5356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5358 = 8'h26 == r_count_26_io_out ? io_r_38_b : _GEN_5357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5359 = 8'h27 == r_count_26_io_out ? io_r_39_b : _GEN_5358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5360 = 8'h28 == r_count_26_io_out ? io_r_40_b : _GEN_5359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5361 = 8'h29 == r_count_26_io_out ? io_r_41_b : _GEN_5360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5362 = 8'h2a == r_count_26_io_out ? io_r_42_b : _GEN_5361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5363 = 8'h2b == r_count_26_io_out ? io_r_43_b : _GEN_5362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5364 = 8'h2c == r_count_26_io_out ? io_r_44_b : _GEN_5363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5365 = 8'h2d == r_count_26_io_out ? io_r_45_b : _GEN_5364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5366 = 8'h2e == r_count_26_io_out ? io_r_46_b : _GEN_5365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5367 = 8'h2f == r_count_26_io_out ? io_r_47_b : _GEN_5366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5368 = 8'h30 == r_count_26_io_out ? io_r_48_b : _GEN_5367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5369 = 8'h31 == r_count_26_io_out ? io_r_49_b : _GEN_5368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5370 = 8'h32 == r_count_26_io_out ? io_r_50_b : _GEN_5369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5371 = 8'h33 == r_count_26_io_out ? io_r_51_b : _GEN_5370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5372 = 8'h34 == r_count_26_io_out ? io_r_52_b : _GEN_5371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5373 = 8'h35 == r_count_26_io_out ? io_r_53_b : _GEN_5372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5374 = 8'h36 == r_count_26_io_out ? io_r_54_b : _GEN_5373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5375 = 8'h37 == r_count_26_io_out ? io_r_55_b : _GEN_5374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5376 = 8'h38 == r_count_26_io_out ? io_r_56_b : _GEN_5375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5377 = 8'h39 == r_count_26_io_out ? io_r_57_b : _GEN_5376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5378 = 8'h3a == r_count_26_io_out ? io_r_58_b : _GEN_5377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5379 = 8'h3b == r_count_26_io_out ? io_r_59_b : _GEN_5378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5380 = 8'h3c == r_count_26_io_out ? io_r_60_b : _GEN_5379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5381 = 8'h3d == r_count_26_io_out ? io_r_61_b : _GEN_5380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5382 = 8'h3e == r_count_26_io_out ? io_r_62_b : _GEN_5381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5383 = 8'h3f == r_count_26_io_out ? io_r_63_b : _GEN_5382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5384 = 8'h40 == r_count_26_io_out ? io_r_64_b : _GEN_5383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5385 = 8'h41 == r_count_26_io_out ? io_r_65_b : _GEN_5384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5386 = 8'h42 == r_count_26_io_out ? io_r_66_b : _GEN_5385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5387 = 8'h43 == r_count_26_io_out ? io_r_67_b : _GEN_5386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5388 = 8'h44 == r_count_26_io_out ? io_r_68_b : _GEN_5387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5389 = 8'h45 == r_count_26_io_out ? io_r_69_b : _GEN_5388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5390 = 8'h46 == r_count_26_io_out ? io_r_70_b : _GEN_5389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5391 = 8'h47 == r_count_26_io_out ? io_r_71_b : _GEN_5390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5392 = 8'h48 == r_count_26_io_out ? io_r_72_b : _GEN_5391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5393 = 8'h49 == r_count_26_io_out ? io_r_73_b : _GEN_5392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5394 = 8'h4a == r_count_26_io_out ? io_r_74_b : _GEN_5393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5395 = 8'h4b == r_count_26_io_out ? io_r_75_b : _GEN_5394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5396 = 8'h4c == r_count_26_io_out ? io_r_76_b : _GEN_5395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5397 = 8'h4d == r_count_26_io_out ? io_r_77_b : _GEN_5396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5398 = 8'h4e == r_count_26_io_out ? io_r_78_b : _GEN_5397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5399 = 8'h4f == r_count_26_io_out ? io_r_79_b : _GEN_5398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5400 = 8'h50 == r_count_26_io_out ? io_r_80_b : _GEN_5399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5401 = 8'h51 == r_count_26_io_out ? io_r_81_b : _GEN_5400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5402 = 8'h52 == r_count_26_io_out ? io_r_82_b : _GEN_5401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5403 = 8'h53 == r_count_26_io_out ? io_r_83_b : _GEN_5402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5404 = 8'h54 == r_count_26_io_out ? io_r_84_b : _GEN_5403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5405 = 8'h55 == r_count_26_io_out ? io_r_85_b : _GEN_5404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5406 = 8'h56 == r_count_26_io_out ? io_r_86_b : _GEN_5405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5407 = 8'h57 == r_count_26_io_out ? io_r_87_b : _GEN_5406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5408 = 8'h58 == r_count_26_io_out ? io_r_88_b : _GEN_5407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5409 = 8'h59 == r_count_26_io_out ? io_r_89_b : _GEN_5408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5410 = 8'h5a == r_count_26_io_out ? io_r_90_b : _GEN_5409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5411 = 8'h5b == r_count_26_io_out ? io_r_91_b : _GEN_5410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5412 = 8'h5c == r_count_26_io_out ? io_r_92_b : _GEN_5411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5413 = 8'h5d == r_count_26_io_out ? io_r_93_b : _GEN_5412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5414 = 8'h5e == r_count_26_io_out ? io_r_94_b : _GEN_5413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5415 = 8'h5f == r_count_26_io_out ? io_r_95_b : _GEN_5414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5416 = 8'h60 == r_count_26_io_out ? io_r_96_b : _GEN_5415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5417 = 8'h61 == r_count_26_io_out ? io_r_97_b : _GEN_5416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5418 = 8'h62 == r_count_26_io_out ? io_r_98_b : _GEN_5417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5419 = 8'h63 == r_count_26_io_out ? io_r_99_b : _GEN_5418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5420 = 8'h64 == r_count_26_io_out ? io_r_100_b : _GEN_5419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5421 = 8'h65 == r_count_26_io_out ? io_r_101_b : _GEN_5420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5422 = 8'h66 == r_count_26_io_out ? io_r_102_b : _GEN_5421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5423 = 8'h67 == r_count_26_io_out ? io_r_103_b : _GEN_5422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5424 = 8'h68 == r_count_26_io_out ? io_r_104_b : _GEN_5423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5425 = 8'h69 == r_count_26_io_out ? io_r_105_b : _GEN_5424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5426 = 8'h6a == r_count_26_io_out ? io_r_106_b : _GEN_5425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5427 = 8'h6b == r_count_26_io_out ? io_r_107_b : _GEN_5426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5428 = 8'h6c == r_count_26_io_out ? io_r_108_b : _GEN_5427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5429 = 8'h6d == r_count_26_io_out ? io_r_109_b : _GEN_5428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5430 = 8'h6e == r_count_26_io_out ? io_r_110_b : _GEN_5429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5431 = 8'h6f == r_count_26_io_out ? io_r_111_b : _GEN_5430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5432 = 8'h70 == r_count_26_io_out ? io_r_112_b : _GEN_5431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5433 = 8'h71 == r_count_26_io_out ? io_r_113_b : _GEN_5432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5434 = 8'h72 == r_count_26_io_out ? io_r_114_b : _GEN_5433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5435 = 8'h73 == r_count_26_io_out ? io_r_115_b : _GEN_5434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5436 = 8'h74 == r_count_26_io_out ? io_r_116_b : _GEN_5435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5437 = 8'h75 == r_count_26_io_out ? io_r_117_b : _GEN_5436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5438 = 8'h76 == r_count_26_io_out ? io_r_118_b : _GEN_5437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5439 = 8'h77 == r_count_26_io_out ? io_r_119_b : _GEN_5438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5440 = 8'h78 == r_count_26_io_out ? io_r_120_b : _GEN_5439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5441 = 8'h79 == r_count_26_io_out ? io_r_121_b : _GEN_5440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5442 = 8'h7a == r_count_26_io_out ? io_r_122_b : _GEN_5441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5443 = 8'h7b == r_count_26_io_out ? io_r_123_b : _GEN_5442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5444 = 8'h7c == r_count_26_io_out ? io_r_124_b : _GEN_5443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5445 = 8'h7d == r_count_26_io_out ? io_r_125_b : _GEN_5444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5446 = 8'h7e == r_count_26_io_out ? io_r_126_b : _GEN_5445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5447 = 8'h7f == r_count_26_io_out ? io_r_127_b : _GEN_5446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5448 = 8'h80 == r_count_26_io_out ? io_r_128_b : _GEN_5447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5449 = 8'h81 == r_count_26_io_out ? io_r_129_b : _GEN_5448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5450 = 8'h82 == r_count_26_io_out ? io_r_130_b : _GEN_5449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5451 = 8'h83 == r_count_26_io_out ? io_r_131_b : _GEN_5450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5452 = 8'h84 == r_count_26_io_out ? io_r_132_b : _GEN_5451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5453 = 8'h85 == r_count_26_io_out ? io_r_133_b : _GEN_5452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5454 = 8'h86 == r_count_26_io_out ? io_r_134_b : _GEN_5453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5455 = 8'h87 == r_count_26_io_out ? io_r_135_b : _GEN_5454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5456 = 8'h88 == r_count_26_io_out ? io_r_136_b : _GEN_5455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5457 = 8'h89 == r_count_26_io_out ? io_r_137_b : _GEN_5456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5458 = 8'h8a == r_count_26_io_out ? io_r_138_b : _GEN_5457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5459 = 8'h8b == r_count_26_io_out ? io_r_139_b : _GEN_5458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5460 = 8'h8c == r_count_26_io_out ? io_r_140_b : _GEN_5459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5461 = 8'h8d == r_count_26_io_out ? io_r_141_b : _GEN_5460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5462 = 8'h8e == r_count_26_io_out ? io_r_142_b : _GEN_5461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5463 = 8'h8f == r_count_26_io_out ? io_r_143_b : _GEN_5462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5464 = 8'h90 == r_count_26_io_out ? io_r_144_b : _GEN_5463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5465 = 8'h91 == r_count_26_io_out ? io_r_145_b : _GEN_5464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5466 = 8'h92 == r_count_26_io_out ? io_r_146_b : _GEN_5465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5467 = 8'h93 == r_count_26_io_out ? io_r_147_b : _GEN_5466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5468 = 8'h94 == r_count_26_io_out ? io_r_148_b : _GEN_5467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5469 = 8'h95 == r_count_26_io_out ? io_r_149_b : _GEN_5468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5470 = 8'h96 == r_count_26_io_out ? io_r_150_b : _GEN_5469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5471 = 8'h97 == r_count_26_io_out ? io_r_151_b : _GEN_5470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5472 = 8'h98 == r_count_26_io_out ? io_r_152_b : _GEN_5471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5473 = 8'h99 == r_count_26_io_out ? io_r_153_b : _GEN_5472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5474 = 8'h9a == r_count_26_io_out ? io_r_154_b : _GEN_5473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5475 = 8'h9b == r_count_26_io_out ? io_r_155_b : _GEN_5474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5476 = 8'h9c == r_count_26_io_out ? io_r_156_b : _GEN_5475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5477 = 8'h9d == r_count_26_io_out ? io_r_157_b : _GEN_5476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5478 = 8'h9e == r_count_26_io_out ? io_r_158_b : _GEN_5477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5479 = 8'h9f == r_count_26_io_out ? io_r_159_b : _GEN_5478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5480 = 8'ha0 == r_count_26_io_out ? io_r_160_b : _GEN_5479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5481 = 8'ha1 == r_count_26_io_out ? io_r_161_b : _GEN_5480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5482 = 8'ha2 == r_count_26_io_out ? io_r_162_b : _GEN_5481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5483 = 8'ha3 == r_count_26_io_out ? io_r_163_b : _GEN_5482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5484 = 8'ha4 == r_count_26_io_out ? io_r_164_b : _GEN_5483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5485 = 8'ha5 == r_count_26_io_out ? io_r_165_b : _GEN_5484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5486 = 8'ha6 == r_count_26_io_out ? io_r_166_b : _GEN_5485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5487 = 8'ha7 == r_count_26_io_out ? io_r_167_b : _GEN_5486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5488 = 8'ha8 == r_count_26_io_out ? io_r_168_b : _GEN_5487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5489 = 8'ha9 == r_count_26_io_out ? io_r_169_b : _GEN_5488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5490 = 8'haa == r_count_26_io_out ? io_r_170_b : _GEN_5489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5491 = 8'hab == r_count_26_io_out ? io_r_171_b : _GEN_5490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5492 = 8'hac == r_count_26_io_out ? io_r_172_b : _GEN_5491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5493 = 8'had == r_count_26_io_out ? io_r_173_b : _GEN_5492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5494 = 8'hae == r_count_26_io_out ? io_r_174_b : _GEN_5493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5495 = 8'haf == r_count_26_io_out ? io_r_175_b : _GEN_5494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5496 = 8'hb0 == r_count_26_io_out ? io_r_176_b : _GEN_5495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5497 = 8'hb1 == r_count_26_io_out ? io_r_177_b : _GEN_5496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5498 = 8'hb2 == r_count_26_io_out ? io_r_178_b : _GEN_5497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5499 = 8'hb3 == r_count_26_io_out ? io_r_179_b : _GEN_5498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5500 = 8'hb4 == r_count_26_io_out ? io_r_180_b : _GEN_5499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5501 = 8'hb5 == r_count_26_io_out ? io_r_181_b : _GEN_5500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5502 = 8'hb6 == r_count_26_io_out ? io_r_182_b : _GEN_5501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5503 = 8'hb7 == r_count_26_io_out ? io_r_183_b : _GEN_5502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5504 = 8'hb8 == r_count_26_io_out ? io_r_184_b : _GEN_5503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5505 = 8'hb9 == r_count_26_io_out ? io_r_185_b : _GEN_5504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5506 = 8'hba == r_count_26_io_out ? io_r_186_b : _GEN_5505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5507 = 8'hbb == r_count_26_io_out ? io_r_187_b : _GEN_5506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5508 = 8'hbc == r_count_26_io_out ? io_r_188_b : _GEN_5507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5509 = 8'hbd == r_count_26_io_out ? io_r_189_b : _GEN_5508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5510 = 8'hbe == r_count_26_io_out ? io_r_190_b : _GEN_5509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5511 = 8'hbf == r_count_26_io_out ? io_r_191_b : _GEN_5510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5512 = 8'hc0 == r_count_26_io_out ? io_r_192_b : _GEN_5511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5513 = 8'hc1 == r_count_26_io_out ? io_r_193_b : _GEN_5512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5514 = 8'hc2 == r_count_26_io_out ? io_r_194_b : _GEN_5513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5515 = 8'hc3 == r_count_26_io_out ? io_r_195_b : _GEN_5514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5516 = 8'hc4 == r_count_26_io_out ? io_r_196_b : _GEN_5515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5517 = 8'hc5 == r_count_26_io_out ? io_r_197_b : _GEN_5516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5518 = 8'hc6 == r_count_26_io_out ? io_r_198_b : _GEN_5517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5521 = 8'h1 == r_count_27_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5522 = 8'h2 == r_count_27_io_out ? io_r_2_b : _GEN_5521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5523 = 8'h3 == r_count_27_io_out ? io_r_3_b : _GEN_5522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5524 = 8'h4 == r_count_27_io_out ? io_r_4_b : _GEN_5523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5525 = 8'h5 == r_count_27_io_out ? io_r_5_b : _GEN_5524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5526 = 8'h6 == r_count_27_io_out ? io_r_6_b : _GEN_5525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5527 = 8'h7 == r_count_27_io_out ? io_r_7_b : _GEN_5526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5528 = 8'h8 == r_count_27_io_out ? io_r_8_b : _GEN_5527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5529 = 8'h9 == r_count_27_io_out ? io_r_9_b : _GEN_5528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5530 = 8'ha == r_count_27_io_out ? io_r_10_b : _GEN_5529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5531 = 8'hb == r_count_27_io_out ? io_r_11_b : _GEN_5530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5532 = 8'hc == r_count_27_io_out ? io_r_12_b : _GEN_5531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5533 = 8'hd == r_count_27_io_out ? io_r_13_b : _GEN_5532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5534 = 8'he == r_count_27_io_out ? io_r_14_b : _GEN_5533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5535 = 8'hf == r_count_27_io_out ? io_r_15_b : _GEN_5534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5536 = 8'h10 == r_count_27_io_out ? io_r_16_b : _GEN_5535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5537 = 8'h11 == r_count_27_io_out ? io_r_17_b : _GEN_5536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5538 = 8'h12 == r_count_27_io_out ? io_r_18_b : _GEN_5537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5539 = 8'h13 == r_count_27_io_out ? io_r_19_b : _GEN_5538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5540 = 8'h14 == r_count_27_io_out ? io_r_20_b : _GEN_5539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5541 = 8'h15 == r_count_27_io_out ? io_r_21_b : _GEN_5540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5542 = 8'h16 == r_count_27_io_out ? io_r_22_b : _GEN_5541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5543 = 8'h17 == r_count_27_io_out ? io_r_23_b : _GEN_5542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5544 = 8'h18 == r_count_27_io_out ? io_r_24_b : _GEN_5543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5545 = 8'h19 == r_count_27_io_out ? io_r_25_b : _GEN_5544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5546 = 8'h1a == r_count_27_io_out ? io_r_26_b : _GEN_5545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5547 = 8'h1b == r_count_27_io_out ? io_r_27_b : _GEN_5546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5548 = 8'h1c == r_count_27_io_out ? io_r_28_b : _GEN_5547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5549 = 8'h1d == r_count_27_io_out ? io_r_29_b : _GEN_5548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5550 = 8'h1e == r_count_27_io_out ? io_r_30_b : _GEN_5549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5551 = 8'h1f == r_count_27_io_out ? io_r_31_b : _GEN_5550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5552 = 8'h20 == r_count_27_io_out ? io_r_32_b : _GEN_5551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5553 = 8'h21 == r_count_27_io_out ? io_r_33_b : _GEN_5552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5554 = 8'h22 == r_count_27_io_out ? io_r_34_b : _GEN_5553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5555 = 8'h23 == r_count_27_io_out ? io_r_35_b : _GEN_5554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5556 = 8'h24 == r_count_27_io_out ? io_r_36_b : _GEN_5555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5557 = 8'h25 == r_count_27_io_out ? io_r_37_b : _GEN_5556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5558 = 8'h26 == r_count_27_io_out ? io_r_38_b : _GEN_5557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5559 = 8'h27 == r_count_27_io_out ? io_r_39_b : _GEN_5558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5560 = 8'h28 == r_count_27_io_out ? io_r_40_b : _GEN_5559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5561 = 8'h29 == r_count_27_io_out ? io_r_41_b : _GEN_5560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5562 = 8'h2a == r_count_27_io_out ? io_r_42_b : _GEN_5561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5563 = 8'h2b == r_count_27_io_out ? io_r_43_b : _GEN_5562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5564 = 8'h2c == r_count_27_io_out ? io_r_44_b : _GEN_5563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5565 = 8'h2d == r_count_27_io_out ? io_r_45_b : _GEN_5564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5566 = 8'h2e == r_count_27_io_out ? io_r_46_b : _GEN_5565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5567 = 8'h2f == r_count_27_io_out ? io_r_47_b : _GEN_5566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5568 = 8'h30 == r_count_27_io_out ? io_r_48_b : _GEN_5567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5569 = 8'h31 == r_count_27_io_out ? io_r_49_b : _GEN_5568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5570 = 8'h32 == r_count_27_io_out ? io_r_50_b : _GEN_5569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5571 = 8'h33 == r_count_27_io_out ? io_r_51_b : _GEN_5570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5572 = 8'h34 == r_count_27_io_out ? io_r_52_b : _GEN_5571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5573 = 8'h35 == r_count_27_io_out ? io_r_53_b : _GEN_5572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5574 = 8'h36 == r_count_27_io_out ? io_r_54_b : _GEN_5573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5575 = 8'h37 == r_count_27_io_out ? io_r_55_b : _GEN_5574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5576 = 8'h38 == r_count_27_io_out ? io_r_56_b : _GEN_5575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5577 = 8'h39 == r_count_27_io_out ? io_r_57_b : _GEN_5576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5578 = 8'h3a == r_count_27_io_out ? io_r_58_b : _GEN_5577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5579 = 8'h3b == r_count_27_io_out ? io_r_59_b : _GEN_5578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5580 = 8'h3c == r_count_27_io_out ? io_r_60_b : _GEN_5579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5581 = 8'h3d == r_count_27_io_out ? io_r_61_b : _GEN_5580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5582 = 8'h3e == r_count_27_io_out ? io_r_62_b : _GEN_5581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5583 = 8'h3f == r_count_27_io_out ? io_r_63_b : _GEN_5582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5584 = 8'h40 == r_count_27_io_out ? io_r_64_b : _GEN_5583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5585 = 8'h41 == r_count_27_io_out ? io_r_65_b : _GEN_5584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5586 = 8'h42 == r_count_27_io_out ? io_r_66_b : _GEN_5585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5587 = 8'h43 == r_count_27_io_out ? io_r_67_b : _GEN_5586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5588 = 8'h44 == r_count_27_io_out ? io_r_68_b : _GEN_5587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5589 = 8'h45 == r_count_27_io_out ? io_r_69_b : _GEN_5588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5590 = 8'h46 == r_count_27_io_out ? io_r_70_b : _GEN_5589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5591 = 8'h47 == r_count_27_io_out ? io_r_71_b : _GEN_5590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5592 = 8'h48 == r_count_27_io_out ? io_r_72_b : _GEN_5591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5593 = 8'h49 == r_count_27_io_out ? io_r_73_b : _GEN_5592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5594 = 8'h4a == r_count_27_io_out ? io_r_74_b : _GEN_5593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5595 = 8'h4b == r_count_27_io_out ? io_r_75_b : _GEN_5594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5596 = 8'h4c == r_count_27_io_out ? io_r_76_b : _GEN_5595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5597 = 8'h4d == r_count_27_io_out ? io_r_77_b : _GEN_5596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5598 = 8'h4e == r_count_27_io_out ? io_r_78_b : _GEN_5597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5599 = 8'h4f == r_count_27_io_out ? io_r_79_b : _GEN_5598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5600 = 8'h50 == r_count_27_io_out ? io_r_80_b : _GEN_5599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5601 = 8'h51 == r_count_27_io_out ? io_r_81_b : _GEN_5600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5602 = 8'h52 == r_count_27_io_out ? io_r_82_b : _GEN_5601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5603 = 8'h53 == r_count_27_io_out ? io_r_83_b : _GEN_5602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5604 = 8'h54 == r_count_27_io_out ? io_r_84_b : _GEN_5603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5605 = 8'h55 == r_count_27_io_out ? io_r_85_b : _GEN_5604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5606 = 8'h56 == r_count_27_io_out ? io_r_86_b : _GEN_5605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5607 = 8'h57 == r_count_27_io_out ? io_r_87_b : _GEN_5606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5608 = 8'h58 == r_count_27_io_out ? io_r_88_b : _GEN_5607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5609 = 8'h59 == r_count_27_io_out ? io_r_89_b : _GEN_5608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5610 = 8'h5a == r_count_27_io_out ? io_r_90_b : _GEN_5609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5611 = 8'h5b == r_count_27_io_out ? io_r_91_b : _GEN_5610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5612 = 8'h5c == r_count_27_io_out ? io_r_92_b : _GEN_5611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5613 = 8'h5d == r_count_27_io_out ? io_r_93_b : _GEN_5612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5614 = 8'h5e == r_count_27_io_out ? io_r_94_b : _GEN_5613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5615 = 8'h5f == r_count_27_io_out ? io_r_95_b : _GEN_5614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5616 = 8'h60 == r_count_27_io_out ? io_r_96_b : _GEN_5615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5617 = 8'h61 == r_count_27_io_out ? io_r_97_b : _GEN_5616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5618 = 8'h62 == r_count_27_io_out ? io_r_98_b : _GEN_5617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5619 = 8'h63 == r_count_27_io_out ? io_r_99_b : _GEN_5618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5620 = 8'h64 == r_count_27_io_out ? io_r_100_b : _GEN_5619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5621 = 8'h65 == r_count_27_io_out ? io_r_101_b : _GEN_5620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5622 = 8'h66 == r_count_27_io_out ? io_r_102_b : _GEN_5621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5623 = 8'h67 == r_count_27_io_out ? io_r_103_b : _GEN_5622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5624 = 8'h68 == r_count_27_io_out ? io_r_104_b : _GEN_5623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5625 = 8'h69 == r_count_27_io_out ? io_r_105_b : _GEN_5624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5626 = 8'h6a == r_count_27_io_out ? io_r_106_b : _GEN_5625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5627 = 8'h6b == r_count_27_io_out ? io_r_107_b : _GEN_5626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5628 = 8'h6c == r_count_27_io_out ? io_r_108_b : _GEN_5627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5629 = 8'h6d == r_count_27_io_out ? io_r_109_b : _GEN_5628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5630 = 8'h6e == r_count_27_io_out ? io_r_110_b : _GEN_5629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5631 = 8'h6f == r_count_27_io_out ? io_r_111_b : _GEN_5630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5632 = 8'h70 == r_count_27_io_out ? io_r_112_b : _GEN_5631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5633 = 8'h71 == r_count_27_io_out ? io_r_113_b : _GEN_5632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5634 = 8'h72 == r_count_27_io_out ? io_r_114_b : _GEN_5633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5635 = 8'h73 == r_count_27_io_out ? io_r_115_b : _GEN_5634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5636 = 8'h74 == r_count_27_io_out ? io_r_116_b : _GEN_5635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5637 = 8'h75 == r_count_27_io_out ? io_r_117_b : _GEN_5636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5638 = 8'h76 == r_count_27_io_out ? io_r_118_b : _GEN_5637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5639 = 8'h77 == r_count_27_io_out ? io_r_119_b : _GEN_5638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5640 = 8'h78 == r_count_27_io_out ? io_r_120_b : _GEN_5639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5641 = 8'h79 == r_count_27_io_out ? io_r_121_b : _GEN_5640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5642 = 8'h7a == r_count_27_io_out ? io_r_122_b : _GEN_5641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5643 = 8'h7b == r_count_27_io_out ? io_r_123_b : _GEN_5642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5644 = 8'h7c == r_count_27_io_out ? io_r_124_b : _GEN_5643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5645 = 8'h7d == r_count_27_io_out ? io_r_125_b : _GEN_5644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5646 = 8'h7e == r_count_27_io_out ? io_r_126_b : _GEN_5645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5647 = 8'h7f == r_count_27_io_out ? io_r_127_b : _GEN_5646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5648 = 8'h80 == r_count_27_io_out ? io_r_128_b : _GEN_5647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5649 = 8'h81 == r_count_27_io_out ? io_r_129_b : _GEN_5648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5650 = 8'h82 == r_count_27_io_out ? io_r_130_b : _GEN_5649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5651 = 8'h83 == r_count_27_io_out ? io_r_131_b : _GEN_5650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5652 = 8'h84 == r_count_27_io_out ? io_r_132_b : _GEN_5651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5653 = 8'h85 == r_count_27_io_out ? io_r_133_b : _GEN_5652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5654 = 8'h86 == r_count_27_io_out ? io_r_134_b : _GEN_5653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5655 = 8'h87 == r_count_27_io_out ? io_r_135_b : _GEN_5654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5656 = 8'h88 == r_count_27_io_out ? io_r_136_b : _GEN_5655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5657 = 8'h89 == r_count_27_io_out ? io_r_137_b : _GEN_5656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5658 = 8'h8a == r_count_27_io_out ? io_r_138_b : _GEN_5657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5659 = 8'h8b == r_count_27_io_out ? io_r_139_b : _GEN_5658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5660 = 8'h8c == r_count_27_io_out ? io_r_140_b : _GEN_5659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5661 = 8'h8d == r_count_27_io_out ? io_r_141_b : _GEN_5660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5662 = 8'h8e == r_count_27_io_out ? io_r_142_b : _GEN_5661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5663 = 8'h8f == r_count_27_io_out ? io_r_143_b : _GEN_5662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5664 = 8'h90 == r_count_27_io_out ? io_r_144_b : _GEN_5663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5665 = 8'h91 == r_count_27_io_out ? io_r_145_b : _GEN_5664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5666 = 8'h92 == r_count_27_io_out ? io_r_146_b : _GEN_5665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5667 = 8'h93 == r_count_27_io_out ? io_r_147_b : _GEN_5666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5668 = 8'h94 == r_count_27_io_out ? io_r_148_b : _GEN_5667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5669 = 8'h95 == r_count_27_io_out ? io_r_149_b : _GEN_5668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5670 = 8'h96 == r_count_27_io_out ? io_r_150_b : _GEN_5669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5671 = 8'h97 == r_count_27_io_out ? io_r_151_b : _GEN_5670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5672 = 8'h98 == r_count_27_io_out ? io_r_152_b : _GEN_5671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5673 = 8'h99 == r_count_27_io_out ? io_r_153_b : _GEN_5672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5674 = 8'h9a == r_count_27_io_out ? io_r_154_b : _GEN_5673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5675 = 8'h9b == r_count_27_io_out ? io_r_155_b : _GEN_5674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5676 = 8'h9c == r_count_27_io_out ? io_r_156_b : _GEN_5675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5677 = 8'h9d == r_count_27_io_out ? io_r_157_b : _GEN_5676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5678 = 8'h9e == r_count_27_io_out ? io_r_158_b : _GEN_5677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5679 = 8'h9f == r_count_27_io_out ? io_r_159_b : _GEN_5678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5680 = 8'ha0 == r_count_27_io_out ? io_r_160_b : _GEN_5679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5681 = 8'ha1 == r_count_27_io_out ? io_r_161_b : _GEN_5680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5682 = 8'ha2 == r_count_27_io_out ? io_r_162_b : _GEN_5681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5683 = 8'ha3 == r_count_27_io_out ? io_r_163_b : _GEN_5682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5684 = 8'ha4 == r_count_27_io_out ? io_r_164_b : _GEN_5683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5685 = 8'ha5 == r_count_27_io_out ? io_r_165_b : _GEN_5684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5686 = 8'ha6 == r_count_27_io_out ? io_r_166_b : _GEN_5685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5687 = 8'ha7 == r_count_27_io_out ? io_r_167_b : _GEN_5686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5688 = 8'ha8 == r_count_27_io_out ? io_r_168_b : _GEN_5687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5689 = 8'ha9 == r_count_27_io_out ? io_r_169_b : _GEN_5688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5690 = 8'haa == r_count_27_io_out ? io_r_170_b : _GEN_5689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5691 = 8'hab == r_count_27_io_out ? io_r_171_b : _GEN_5690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5692 = 8'hac == r_count_27_io_out ? io_r_172_b : _GEN_5691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5693 = 8'had == r_count_27_io_out ? io_r_173_b : _GEN_5692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5694 = 8'hae == r_count_27_io_out ? io_r_174_b : _GEN_5693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5695 = 8'haf == r_count_27_io_out ? io_r_175_b : _GEN_5694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5696 = 8'hb0 == r_count_27_io_out ? io_r_176_b : _GEN_5695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5697 = 8'hb1 == r_count_27_io_out ? io_r_177_b : _GEN_5696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5698 = 8'hb2 == r_count_27_io_out ? io_r_178_b : _GEN_5697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5699 = 8'hb3 == r_count_27_io_out ? io_r_179_b : _GEN_5698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5700 = 8'hb4 == r_count_27_io_out ? io_r_180_b : _GEN_5699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5701 = 8'hb5 == r_count_27_io_out ? io_r_181_b : _GEN_5700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5702 = 8'hb6 == r_count_27_io_out ? io_r_182_b : _GEN_5701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5703 = 8'hb7 == r_count_27_io_out ? io_r_183_b : _GEN_5702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5704 = 8'hb8 == r_count_27_io_out ? io_r_184_b : _GEN_5703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5705 = 8'hb9 == r_count_27_io_out ? io_r_185_b : _GEN_5704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5706 = 8'hba == r_count_27_io_out ? io_r_186_b : _GEN_5705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5707 = 8'hbb == r_count_27_io_out ? io_r_187_b : _GEN_5706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5708 = 8'hbc == r_count_27_io_out ? io_r_188_b : _GEN_5707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5709 = 8'hbd == r_count_27_io_out ? io_r_189_b : _GEN_5708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5710 = 8'hbe == r_count_27_io_out ? io_r_190_b : _GEN_5709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5711 = 8'hbf == r_count_27_io_out ? io_r_191_b : _GEN_5710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5712 = 8'hc0 == r_count_27_io_out ? io_r_192_b : _GEN_5711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5713 = 8'hc1 == r_count_27_io_out ? io_r_193_b : _GEN_5712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5714 = 8'hc2 == r_count_27_io_out ? io_r_194_b : _GEN_5713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5715 = 8'hc3 == r_count_27_io_out ? io_r_195_b : _GEN_5714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5716 = 8'hc4 == r_count_27_io_out ? io_r_196_b : _GEN_5715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5717 = 8'hc5 == r_count_27_io_out ? io_r_197_b : _GEN_5716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5718 = 8'hc6 == r_count_27_io_out ? io_r_198_b : _GEN_5717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5721 = 8'h1 == r_count_28_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5722 = 8'h2 == r_count_28_io_out ? io_r_2_b : _GEN_5721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5723 = 8'h3 == r_count_28_io_out ? io_r_3_b : _GEN_5722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5724 = 8'h4 == r_count_28_io_out ? io_r_4_b : _GEN_5723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5725 = 8'h5 == r_count_28_io_out ? io_r_5_b : _GEN_5724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5726 = 8'h6 == r_count_28_io_out ? io_r_6_b : _GEN_5725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5727 = 8'h7 == r_count_28_io_out ? io_r_7_b : _GEN_5726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5728 = 8'h8 == r_count_28_io_out ? io_r_8_b : _GEN_5727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5729 = 8'h9 == r_count_28_io_out ? io_r_9_b : _GEN_5728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5730 = 8'ha == r_count_28_io_out ? io_r_10_b : _GEN_5729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5731 = 8'hb == r_count_28_io_out ? io_r_11_b : _GEN_5730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5732 = 8'hc == r_count_28_io_out ? io_r_12_b : _GEN_5731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5733 = 8'hd == r_count_28_io_out ? io_r_13_b : _GEN_5732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5734 = 8'he == r_count_28_io_out ? io_r_14_b : _GEN_5733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5735 = 8'hf == r_count_28_io_out ? io_r_15_b : _GEN_5734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5736 = 8'h10 == r_count_28_io_out ? io_r_16_b : _GEN_5735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5737 = 8'h11 == r_count_28_io_out ? io_r_17_b : _GEN_5736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5738 = 8'h12 == r_count_28_io_out ? io_r_18_b : _GEN_5737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5739 = 8'h13 == r_count_28_io_out ? io_r_19_b : _GEN_5738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5740 = 8'h14 == r_count_28_io_out ? io_r_20_b : _GEN_5739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5741 = 8'h15 == r_count_28_io_out ? io_r_21_b : _GEN_5740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5742 = 8'h16 == r_count_28_io_out ? io_r_22_b : _GEN_5741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5743 = 8'h17 == r_count_28_io_out ? io_r_23_b : _GEN_5742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5744 = 8'h18 == r_count_28_io_out ? io_r_24_b : _GEN_5743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5745 = 8'h19 == r_count_28_io_out ? io_r_25_b : _GEN_5744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5746 = 8'h1a == r_count_28_io_out ? io_r_26_b : _GEN_5745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5747 = 8'h1b == r_count_28_io_out ? io_r_27_b : _GEN_5746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5748 = 8'h1c == r_count_28_io_out ? io_r_28_b : _GEN_5747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5749 = 8'h1d == r_count_28_io_out ? io_r_29_b : _GEN_5748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5750 = 8'h1e == r_count_28_io_out ? io_r_30_b : _GEN_5749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5751 = 8'h1f == r_count_28_io_out ? io_r_31_b : _GEN_5750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5752 = 8'h20 == r_count_28_io_out ? io_r_32_b : _GEN_5751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5753 = 8'h21 == r_count_28_io_out ? io_r_33_b : _GEN_5752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5754 = 8'h22 == r_count_28_io_out ? io_r_34_b : _GEN_5753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5755 = 8'h23 == r_count_28_io_out ? io_r_35_b : _GEN_5754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5756 = 8'h24 == r_count_28_io_out ? io_r_36_b : _GEN_5755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5757 = 8'h25 == r_count_28_io_out ? io_r_37_b : _GEN_5756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5758 = 8'h26 == r_count_28_io_out ? io_r_38_b : _GEN_5757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5759 = 8'h27 == r_count_28_io_out ? io_r_39_b : _GEN_5758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5760 = 8'h28 == r_count_28_io_out ? io_r_40_b : _GEN_5759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5761 = 8'h29 == r_count_28_io_out ? io_r_41_b : _GEN_5760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5762 = 8'h2a == r_count_28_io_out ? io_r_42_b : _GEN_5761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5763 = 8'h2b == r_count_28_io_out ? io_r_43_b : _GEN_5762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5764 = 8'h2c == r_count_28_io_out ? io_r_44_b : _GEN_5763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5765 = 8'h2d == r_count_28_io_out ? io_r_45_b : _GEN_5764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5766 = 8'h2e == r_count_28_io_out ? io_r_46_b : _GEN_5765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5767 = 8'h2f == r_count_28_io_out ? io_r_47_b : _GEN_5766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5768 = 8'h30 == r_count_28_io_out ? io_r_48_b : _GEN_5767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5769 = 8'h31 == r_count_28_io_out ? io_r_49_b : _GEN_5768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5770 = 8'h32 == r_count_28_io_out ? io_r_50_b : _GEN_5769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5771 = 8'h33 == r_count_28_io_out ? io_r_51_b : _GEN_5770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5772 = 8'h34 == r_count_28_io_out ? io_r_52_b : _GEN_5771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5773 = 8'h35 == r_count_28_io_out ? io_r_53_b : _GEN_5772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5774 = 8'h36 == r_count_28_io_out ? io_r_54_b : _GEN_5773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5775 = 8'h37 == r_count_28_io_out ? io_r_55_b : _GEN_5774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5776 = 8'h38 == r_count_28_io_out ? io_r_56_b : _GEN_5775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5777 = 8'h39 == r_count_28_io_out ? io_r_57_b : _GEN_5776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5778 = 8'h3a == r_count_28_io_out ? io_r_58_b : _GEN_5777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5779 = 8'h3b == r_count_28_io_out ? io_r_59_b : _GEN_5778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5780 = 8'h3c == r_count_28_io_out ? io_r_60_b : _GEN_5779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5781 = 8'h3d == r_count_28_io_out ? io_r_61_b : _GEN_5780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5782 = 8'h3e == r_count_28_io_out ? io_r_62_b : _GEN_5781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5783 = 8'h3f == r_count_28_io_out ? io_r_63_b : _GEN_5782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5784 = 8'h40 == r_count_28_io_out ? io_r_64_b : _GEN_5783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5785 = 8'h41 == r_count_28_io_out ? io_r_65_b : _GEN_5784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5786 = 8'h42 == r_count_28_io_out ? io_r_66_b : _GEN_5785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5787 = 8'h43 == r_count_28_io_out ? io_r_67_b : _GEN_5786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5788 = 8'h44 == r_count_28_io_out ? io_r_68_b : _GEN_5787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5789 = 8'h45 == r_count_28_io_out ? io_r_69_b : _GEN_5788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5790 = 8'h46 == r_count_28_io_out ? io_r_70_b : _GEN_5789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5791 = 8'h47 == r_count_28_io_out ? io_r_71_b : _GEN_5790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5792 = 8'h48 == r_count_28_io_out ? io_r_72_b : _GEN_5791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5793 = 8'h49 == r_count_28_io_out ? io_r_73_b : _GEN_5792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5794 = 8'h4a == r_count_28_io_out ? io_r_74_b : _GEN_5793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5795 = 8'h4b == r_count_28_io_out ? io_r_75_b : _GEN_5794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5796 = 8'h4c == r_count_28_io_out ? io_r_76_b : _GEN_5795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5797 = 8'h4d == r_count_28_io_out ? io_r_77_b : _GEN_5796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5798 = 8'h4e == r_count_28_io_out ? io_r_78_b : _GEN_5797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5799 = 8'h4f == r_count_28_io_out ? io_r_79_b : _GEN_5798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5800 = 8'h50 == r_count_28_io_out ? io_r_80_b : _GEN_5799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5801 = 8'h51 == r_count_28_io_out ? io_r_81_b : _GEN_5800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5802 = 8'h52 == r_count_28_io_out ? io_r_82_b : _GEN_5801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5803 = 8'h53 == r_count_28_io_out ? io_r_83_b : _GEN_5802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5804 = 8'h54 == r_count_28_io_out ? io_r_84_b : _GEN_5803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5805 = 8'h55 == r_count_28_io_out ? io_r_85_b : _GEN_5804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5806 = 8'h56 == r_count_28_io_out ? io_r_86_b : _GEN_5805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5807 = 8'h57 == r_count_28_io_out ? io_r_87_b : _GEN_5806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5808 = 8'h58 == r_count_28_io_out ? io_r_88_b : _GEN_5807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5809 = 8'h59 == r_count_28_io_out ? io_r_89_b : _GEN_5808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5810 = 8'h5a == r_count_28_io_out ? io_r_90_b : _GEN_5809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5811 = 8'h5b == r_count_28_io_out ? io_r_91_b : _GEN_5810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5812 = 8'h5c == r_count_28_io_out ? io_r_92_b : _GEN_5811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5813 = 8'h5d == r_count_28_io_out ? io_r_93_b : _GEN_5812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5814 = 8'h5e == r_count_28_io_out ? io_r_94_b : _GEN_5813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5815 = 8'h5f == r_count_28_io_out ? io_r_95_b : _GEN_5814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5816 = 8'h60 == r_count_28_io_out ? io_r_96_b : _GEN_5815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5817 = 8'h61 == r_count_28_io_out ? io_r_97_b : _GEN_5816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5818 = 8'h62 == r_count_28_io_out ? io_r_98_b : _GEN_5817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5819 = 8'h63 == r_count_28_io_out ? io_r_99_b : _GEN_5818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5820 = 8'h64 == r_count_28_io_out ? io_r_100_b : _GEN_5819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5821 = 8'h65 == r_count_28_io_out ? io_r_101_b : _GEN_5820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5822 = 8'h66 == r_count_28_io_out ? io_r_102_b : _GEN_5821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5823 = 8'h67 == r_count_28_io_out ? io_r_103_b : _GEN_5822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5824 = 8'h68 == r_count_28_io_out ? io_r_104_b : _GEN_5823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5825 = 8'h69 == r_count_28_io_out ? io_r_105_b : _GEN_5824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5826 = 8'h6a == r_count_28_io_out ? io_r_106_b : _GEN_5825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5827 = 8'h6b == r_count_28_io_out ? io_r_107_b : _GEN_5826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5828 = 8'h6c == r_count_28_io_out ? io_r_108_b : _GEN_5827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5829 = 8'h6d == r_count_28_io_out ? io_r_109_b : _GEN_5828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5830 = 8'h6e == r_count_28_io_out ? io_r_110_b : _GEN_5829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5831 = 8'h6f == r_count_28_io_out ? io_r_111_b : _GEN_5830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5832 = 8'h70 == r_count_28_io_out ? io_r_112_b : _GEN_5831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5833 = 8'h71 == r_count_28_io_out ? io_r_113_b : _GEN_5832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5834 = 8'h72 == r_count_28_io_out ? io_r_114_b : _GEN_5833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5835 = 8'h73 == r_count_28_io_out ? io_r_115_b : _GEN_5834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5836 = 8'h74 == r_count_28_io_out ? io_r_116_b : _GEN_5835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5837 = 8'h75 == r_count_28_io_out ? io_r_117_b : _GEN_5836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5838 = 8'h76 == r_count_28_io_out ? io_r_118_b : _GEN_5837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5839 = 8'h77 == r_count_28_io_out ? io_r_119_b : _GEN_5838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5840 = 8'h78 == r_count_28_io_out ? io_r_120_b : _GEN_5839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5841 = 8'h79 == r_count_28_io_out ? io_r_121_b : _GEN_5840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5842 = 8'h7a == r_count_28_io_out ? io_r_122_b : _GEN_5841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5843 = 8'h7b == r_count_28_io_out ? io_r_123_b : _GEN_5842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5844 = 8'h7c == r_count_28_io_out ? io_r_124_b : _GEN_5843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5845 = 8'h7d == r_count_28_io_out ? io_r_125_b : _GEN_5844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5846 = 8'h7e == r_count_28_io_out ? io_r_126_b : _GEN_5845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5847 = 8'h7f == r_count_28_io_out ? io_r_127_b : _GEN_5846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5848 = 8'h80 == r_count_28_io_out ? io_r_128_b : _GEN_5847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5849 = 8'h81 == r_count_28_io_out ? io_r_129_b : _GEN_5848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5850 = 8'h82 == r_count_28_io_out ? io_r_130_b : _GEN_5849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5851 = 8'h83 == r_count_28_io_out ? io_r_131_b : _GEN_5850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5852 = 8'h84 == r_count_28_io_out ? io_r_132_b : _GEN_5851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5853 = 8'h85 == r_count_28_io_out ? io_r_133_b : _GEN_5852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5854 = 8'h86 == r_count_28_io_out ? io_r_134_b : _GEN_5853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5855 = 8'h87 == r_count_28_io_out ? io_r_135_b : _GEN_5854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5856 = 8'h88 == r_count_28_io_out ? io_r_136_b : _GEN_5855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5857 = 8'h89 == r_count_28_io_out ? io_r_137_b : _GEN_5856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5858 = 8'h8a == r_count_28_io_out ? io_r_138_b : _GEN_5857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5859 = 8'h8b == r_count_28_io_out ? io_r_139_b : _GEN_5858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5860 = 8'h8c == r_count_28_io_out ? io_r_140_b : _GEN_5859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5861 = 8'h8d == r_count_28_io_out ? io_r_141_b : _GEN_5860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5862 = 8'h8e == r_count_28_io_out ? io_r_142_b : _GEN_5861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5863 = 8'h8f == r_count_28_io_out ? io_r_143_b : _GEN_5862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5864 = 8'h90 == r_count_28_io_out ? io_r_144_b : _GEN_5863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5865 = 8'h91 == r_count_28_io_out ? io_r_145_b : _GEN_5864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5866 = 8'h92 == r_count_28_io_out ? io_r_146_b : _GEN_5865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5867 = 8'h93 == r_count_28_io_out ? io_r_147_b : _GEN_5866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5868 = 8'h94 == r_count_28_io_out ? io_r_148_b : _GEN_5867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5869 = 8'h95 == r_count_28_io_out ? io_r_149_b : _GEN_5868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5870 = 8'h96 == r_count_28_io_out ? io_r_150_b : _GEN_5869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5871 = 8'h97 == r_count_28_io_out ? io_r_151_b : _GEN_5870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5872 = 8'h98 == r_count_28_io_out ? io_r_152_b : _GEN_5871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5873 = 8'h99 == r_count_28_io_out ? io_r_153_b : _GEN_5872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5874 = 8'h9a == r_count_28_io_out ? io_r_154_b : _GEN_5873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5875 = 8'h9b == r_count_28_io_out ? io_r_155_b : _GEN_5874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5876 = 8'h9c == r_count_28_io_out ? io_r_156_b : _GEN_5875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5877 = 8'h9d == r_count_28_io_out ? io_r_157_b : _GEN_5876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5878 = 8'h9e == r_count_28_io_out ? io_r_158_b : _GEN_5877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5879 = 8'h9f == r_count_28_io_out ? io_r_159_b : _GEN_5878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5880 = 8'ha0 == r_count_28_io_out ? io_r_160_b : _GEN_5879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5881 = 8'ha1 == r_count_28_io_out ? io_r_161_b : _GEN_5880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5882 = 8'ha2 == r_count_28_io_out ? io_r_162_b : _GEN_5881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5883 = 8'ha3 == r_count_28_io_out ? io_r_163_b : _GEN_5882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5884 = 8'ha4 == r_count_28_io_out ? io_r_164_b : _GEN_5883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5885 = 8'ha5 == r_count_28_io_out ? io_r_165_b : _GEN_5884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5886 = 8'ha6 == r_count_28_io_out ? io_r_166_b : _GEN_5885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5887 = 8'ha7 == r_count_28_io_out ? io_r_167_b : _GEN_5886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5888 = 8'ha8 == r_count_28_io_out ? io_r_168_b : _GEN_5887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5889 = 8'ha9 == r_count_28_io_out ? io_r_169_b : _GEN_5888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5890 = 8'haa == r_count_28_io_out ? io_r_170_b : _GEN_5889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5891 = 8'hab == r_count_28_io_out ? io_r_171_b : _GEN_5890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5892 = 8'hac == r_count_28_io_out ? io_r_172_b : _GEN_5891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5893 = 8'had == r_count_28_io_out ? io_r_173_b : _GEN_5892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5894 = 8'hae == r_count_28_io_out ? io_r_174_b : _GEN_5893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5895 = 8'haf == r_count_28_io_out ? io_r_175_b : _GEN_5894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5896 = 8'hb0 == r_count_28_io_out ? io_r_176_b : _GEN_5895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5897 = 8'hb1 == r_count_28_io_out ? io_r_177_b : _GEN_5896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5898 = 8'hb2 == r_count_28_io_out ? io_r_178_b : _GEN_5897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5899 = 8'hb3 == r_count_28_io_out ? io_r_179_b : _GEN_5898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5900 = 8'hb4 == r_count_28_io_out ? io_r_180_b : _GEN_5899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5901 = 8'hb5 == r_count_28_io_out ? io_r_181_b : _GEN_5900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5902 = 8'hb6 == r_count_28_io_out ? io_r_182_b : _GEN_5901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5903 = 8'hb7 == r_count_28_io_out ? io_r_183_b : _GEN_5902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5904 = 8'hb8 == r_count_28_io_out ? io_r_184_b : _GEN_5903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5905 = 8'hb9 == r_count_28_io_out ? io_r_185_b : _GEN_5904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5906 = 8'hba == r_count_28_io_out ? io_r_186_b : _GEN_5905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5907 = 8'hbb == r_count_28_io_out ? io_r_187_b : _GEN_5906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5908 = 8'hbc == r_count_28_io_out ? io_r_188_b : _GEN_5907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5909 = 8'hbd == r_count_28_io_out ? io_r_189_b : _GEN_5908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5910 = 8'hbe == r_count_28_io_out ? io_r_190_b : _GEN_5909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5911 = 8'hbf == r_count_28_io_out ? io_r_191_b : _GEN_5910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5912 = 8'hc0 == r_count_28_io_out ? io_r_192_b : _GEN_5911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5913 = 8'hc1 == r_count_28_io_out ? io_r_193_b : _GEN_5912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5914 = 8'hc2 == r_count_28_io_out ? io_r_194_b : _GEN_5913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5915 = 8'hc3 == r_count_28_io_out ? io_r_195_b : _GEN_5914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5916 = 8'hc4 == r_count_28_io_out ? io_r_196_b : _GEN_5915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5917 = 8'hc5 == r_count_28_io_out ? io_r_197_b : _GEN_5916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5918 = 8'hc6 == r_count_28_io_out ? io_r_198_b : _GEN_5917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5921 = 8'h1 == r_count_29_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5922 = 8'h2 == r_count_29_io_out ? io_r_2_b : _GEN_5921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5923 = 8'h3 == r_count_29_io_out ? io_r_3_b : _GEN_5922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5924 = 8'h4 == r_count_29_io_out ? io_r_4_b : _GEN_5923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5925 = 8'h5 == r_count_29_io_out ? io_r_5_b : _GEN_5924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5926 = 8'h6 == r_count_29_io_out ? io_r_6_b : _GEN_5925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5927 = 8'h7 == r_count_29_io_out ? io_r_7_b : _GEN_5926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5928 = 8'h8 == r_count_29_io_out ? io_r_8_b : _GEN_5927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5929 = 8'h9 == r_count_29_io_out ? io_r_9_b : _GEN_5928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5930 = 8'ha == r_count_29_io_out ? io_r_10_b : _GEN_5929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5931 = 8'hb == r_count_29_io_out ? io_r_11_b : _GEN_5930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5932 = 8'hc == r_count_29_io_out ? io_r_12_b : _GEN_5931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5933 = 8'hd == r_count_29_io_out ? io_r_13_b : _GEN_5932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5934 = 8'he == r_count_29_io_out ? io_r_14_b : _GEN_5933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5935 = 8'hf == r_count_29_io_out ? io_r_15_b : _GEN_5934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5936 = 8'h10 == r_count_29_io_out ? io_r_16_b : _GEN_5935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5937 = 8'h11 == r_count_29_io_out ? io_r_17_b : _GEN_5936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5938 = 8'h12 == r_count_29_io_out ? io_r_18_b : _GEN_5937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5939 = 8'h13 == r_count_29_io_out ? io_r_19_b : _GEN_5938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5940 = 8'h14 == r_count_29_io_out ? io_r_20_b : _GEN_5939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5941 = 8'h15 == r_count_29_io_out ? io_r_21_b : _GEN_5940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5942 = 8'h16 == r_count_29_io_out ? io_r_22_b : _GEN_5941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5943 = 8'h17 == r_count_29_io_out ? io_r_23_b : _GEN_5942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5944 = 8'h18 == r_count_29_io_out ? io_r_24_b : _GEN_5943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5945 = 8'h19 == r_count_29_io_out ? io_r_25_b : _GEN_5944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5946 = 8'h1a == r_count_29_io_out ? io_r_26_b : _GEN_5945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5947 = 8'h1b == r_count_29_io_out ? io_r_27_b : _GEN_5946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5948 = 8'h1c == r_count_29_io_out ? io_r_28_b : _GEN_5947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5949 = 8'h1d == r_count_29_io_out ? io_r_29_b : _GEN_5948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5950 = 8'h1e == r_count_29_io_out ? io_r_30_b : _GEN_5949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5951 = 8'h1f == r_count_29_io_out ? io_r_31_b : _GEN_5950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5952 = 8'h20 == r_count_29_io_out ? io_r_32_b : _GEN_5951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5953 = 8'h21 == r_count_29_io_out ? io_r_33_b : _GEN_5952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5954 = 8'h22 == r_count_29_io_out ? io_r_34_b : _GEN_5953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5955 = 8'h23 == r_count_29_io_out ? io_r_35_b : _GEN_5954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5956 = 8'h24 == r_count_29_io_out ? io_r_36_b : _GEN_5955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5957 = 8'h25 == r_count_29_io_out ? io_r_37_b : _GEN_5956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5958 = 8'h26 == r_count_29_io_out ? io_r_38_b : _GEN_5957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5959 = 8'h27 == r_count_29_io_out ? io_r_39_b : _GEN_5958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5960 = 8'h28 == r_count_29_io_out ? io_r_40_b : _GEN_5959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5961 = 8'h29 == r_count_29_io_out ? io_r_41_b : _GEN_5960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5962 = 8'h2a == r_count_29_io_out ? io_r_42_b : _GEN_5961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5963 = 8'h2b == r_count_29_io_out ? io_r_43_b : _GEN_5962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5964 = 8'h2c == r_count_29_io_out ? io_r_44_b : _GEN_5963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5965 = 8'h2d == r_count_29_io_out ? io_r_45_b : _GEN_5964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5966 = 8'h2e == r_count_29_io_out ? io_r_46_b : _GEN_5965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5967 = 8'h2f == r_count_29_io_out ? io_r_47_b : _GEN_5966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5968 = 8'h30 == r_count_29_io_out ? io_r_48_b : _GEN_5967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5969 = 8'h31 == r_count_29_io_out ? io_r_49_b : _GEN_5968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5970 = 8'h32 == r_count_29_io_out ? io_r_50_b : _GEN_5969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5971 = 8'h33 == r_count_29_io_out ? io_r_51_b : _GEN_5970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5972 = 8'h34 == r_count_29_io_out ? io_r_52_b : _GEN_5971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5973 = 8'h35 == r_count_29_io_out ? io_r_53_b : _GEN_5972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5974 = 8'h36 == r_count_29_io_out ? io_r_54_b : _GEN_5973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5975 = 8'h37 == r_count_29_io_out ? io_r_55_b : _GEN_5974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5976 = 8'h38 == r_count_29_io_out ? io_r_56_b : _GEN_5975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5977 = 8'h39 == r_count_29_io_out ? io_r_57_b : _GEN_5976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5978 = 8'h3a == r_count_29_io_out ? io_r_58_b : _GEN_5977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5979 = 8'h3b == r_count_29_io_out ? io_r_59_b : _GEN_5978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5980 = 8'h3c == r_count_29_io_out ? io_r_60_b : _GEN_5979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5981 = 8'h3d == r_count_29_io_out ? io_r_61_b : _GEN_5980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5982 = 8'h3e == r_count_29_io_out ? io_r_62_b : _GEN_5981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5983 = 8'h3f == r_count_29_io_out ? io_r_63_b : _GEN_5982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5984 = 8'h40 == r_count_29_io_out ? io_r_64_b : _GEN_5983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5985 = 8'h41 == r_count_29_io_out ? io_r_65_b : _GEN_5984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5986 = 8'h42 == r_count_29_io_out ? io_r_66_b : _GEN_5985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5987 = 8'h43 == r_count_29_io_out ? io_r_67_b : _GEN_5986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5988 = 8'h44 == r_count_29_io_out ? io_r_68_b : _GEN_5987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5989 = 8'h45 == r_count_29_io_out ? io_r_69_b : _GEN_5988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5990 = 8'h46 == r_count_29_io_out ? io_r_70_b : _GEN_5989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5991 = 8'h47 == r_count_29_io_out ? io_r_71_b : _GEN_5990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5992 = 8'h48 == r_count_29_io_out ? io_r_72_b : _GEN_5991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5993 = 8'h49 == r_count_29_io_out ? io_r_73_b : _GEN_5992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5994 = 8'h4a == r_count_29_io_out ? io_r_74_b : _GEN_5993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5995 = 8'h4b == r_count_29_io_out ? io_r_75_b : _GEN_5994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5996 = 8'h4c == r_count_29_io_out ? io_r_76_b : _GEN_5995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5997 = 8'h4d == r_count_29_io_out ? io_r_77_b : _GEN_5996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5998 = 8'h4e == r_count_29_io_out ? io_r_78_b : _GEN_5997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5999 = 8'h4f == r_count_29_io_out ? io_r_79_b : _GEN_5998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6000 = 8'h50 == r_count_29_io_out ? io_r_80_b : _GEN_5999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6001 = 8'h51 == r_count_29_io_out ? io_r_81_b : _GEN_6000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6002 = 8'h52 == r_count_29_io_out ? io_r_82_b : _GEN_6001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6003 = 8'h53 == r_count_29_io_out ? io_r_83_b : _GEN_6002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6004 = 8'h54 == r_count_29_io_out ? io_r_84_b : _GEN_6003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6005 = 8'h55 == r_count_29_io_out ? io_r_85_b : _GEN_6004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6006 = 8'h56 == r_count_29_io_out ? io_r_86_b : _GEN_6005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6007 = 8'h57 == r_count_29_io_out ? io_r_87_b : _GEN_6006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6008 = 8'h58 == r_count_29_io_out ? io_r_88_b : _GEN_6007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6009 = 8'h59 == r_count_29_io_out ? io_r_89_b : _GEN_6008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6010 = 8'h5a == r_count_29_io_out ? io_r_90_b : _GEN_6009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6011 = 8'h5b == r_count_29_io_out ? io_r_91_b : _GEN_6010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6012 = 8'h5c == r_count_29_io_out ? io_r_92_b : _GEN_6011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6013 = 8'h5d == r_count_29_io_out ? io_r_93_b : _GEN_6012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6014 = 8'h5e == r_count_29_io_out ? io_r_94_b : _GEN_6013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6015 = 8'h5f == r_count_29_io_out ? io_r_95_b : _GEN_6014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6016 = 8'h60 == r_count_29_io_out ? io_r_96_b : _GEN_6015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6017 = 8'h61 == r_count_29_io_out ? io_r_97_b : _GEN_6016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6018 = 8'h62 == r_count_29_io_out ? io_r_98_b : _GEN_6017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6019 = 8'h63 == r_count_29_io_out ? io_r_99_b : _GEN_6018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6020 = 8'h64 == r_count_29_io_out ? io_r_100_b : _GEN_6019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6021 = 8'h65 == r_count_29_io_out ? io_r_101_b : _GEN_6020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6022 = 8'h66 == r_count_29_io_out ? io_r_102_b : _GEN_6021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6023 = 8'h67 == r_count_29_io_out ? io_r_103_b : _GEN_6022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6024 = 8'h68 == r_count_29_io_out ? io_r_104_b : _GEN_6023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6025 = 8'h69 == r_count_29_io_out ? io_r_105_b : _GEN_6024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6026 = 8'h6a == r_count_29_io_out ? io_r_106_b : _GEN_6025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6027 = 8'h6b == r_count_29_io_out ? io_r_107_b : _GEN_6026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6028 = 8'h6c == r_count_29_io_out ? io_r_108_b : _GEN_6027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6029 = 8'h6d == r_count_29_io_out ? io_r_109_b : _GEN_6028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6030 = 8'h6e == r_count_29_io_out ? io_r_110_b : _GEN_6029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6031 = 8'h6f == r_count_29_io_out ? io_r_111_b : _GEN_6030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6032 = 8'h70 == r_count_29_io_out ? io_r_112_b : _GEN_6031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6033 = 8'h71 == r_count_29_io_out ? io_r_113_b : _GEN_6032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6034 = 8'h72 == r_count_29_io_out ? io_r_114_b : _GEN_6033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6035 = 8'h73 == r_count_29_io_out ? io_r_115_b : _GEN_6034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6036 = 8'h74 == r_count_29_io_out ? io_r_116_b : _GEN_6035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6037 = 8'h75 == r_count_29_io_out ? io_r_117_b : _GEN_6036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6038 = 8'h76 == r_count_29_io_out ? io_r_118_b : _GEN_6037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6039 = 8'h77 == r_count_29_io_out ? io_r_119_b : _GEN_6038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6040 = 8'h78 == r_count_29_io_out ? io_r_120_b : _GEN_6039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6041 = 8'h79 == r_count_29_io_out ? io_r_121_b : _GEN_6040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6042 = 8'h7a == r_count_29_io_out ? io_r_122_b : _GEN_6041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6043 = 8'h7b == r_count_29_io_out ? io_r_123_b : _GEN_6042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6044 = 8'h7c == r_count_29_io_out ? io_r_124_b : _GEN_6043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6045 = 8'h7d == r_count_29_io_out ? io_r_125_b : _GEN_6044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6046 = 8'h7e == r_count_29_io_out ? io_r_126_b : _GEN_6045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6047 = 8'h7f == r_count_29_io_out ? io_r_127_b : _GEN_6046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6048 = 8'h80 == r_count_29_io_out ? io_r_128_b : _GEN_6047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6049 = 8'h81 == r_count_29_io_out ? io_r_129_b : _GEN_6048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6050 = 8'h82 == r_count_29_io_out ? io_r_130_b : _GEN_6049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6051 = 8'h83 == r_count_29_io_out ? io_r_131_b : _GEN_6050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6052 = 8'h84 == r_count_29_io_out ? io_r_132_b : _GEN_6051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6053 = 8'h85 == r_count_29_io_out ? io_r_133_b : _GEN_6052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6054 = 8'h86 == r_count_29_io_out ? io_r_134_b : _GEN_6053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6055 = 8'h87 == r_count_29_io_out ? io_r_135_b : _GEN_6054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6056 = 8'h88 == r_count_29_io_out ? io_r_136_b : _GEN_6055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6057 = 8'h89 == r_count_29_io_out ? io_r_137_b : _GEN_6056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6058 = 8'h8a == r_count_29_io_out ? io_r_138_b : _GEN_6057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6059 = 8'h8b == r_count_29_io_out ? io_r_139_b : _GEN_6058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6060 = 8'h8c == r_count_29_io_out ? io_r_140_b : _GEN_6059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6061 = 8'h8d == r_count_29_io_out ? io_r_141_b : _GEN_6060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6062 = 8'h8e == r_count_29_io_out ? io_r_142_b : _GEN_6061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6063 = 8'h8f == r_count_29_io_out ? io_r_143_b : _GEN_6062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6064 = 8'h90 == r_count_29_io_out ? io_r_144_b : _GEN_6063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6065 = 8'h91 == r_count_29_io_out ? io_r_145_b : _GEN_6064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6066 = 8'h92 == r_count_29_io_out ? io_r_146_b : _GEN_6065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6067 = 8'h93 == r_count_29_io_out ? io_r_147_b : _GEN_6066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6068 = 8'h94 == r_count_29_io_out ? io_r_148_b : _GEN_6067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6069 = 8'h95 == r_count_29_io_out ? io_r_149_b : _GEN_6068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6070 = 8'h96 == r_count_29_io_out ? io_r_150_b : _GEN_6069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6071 = 8'h97 == r_count_29_io_out ? io_r_151_b : _GEN_6070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6072 = 8'h98 == r_count_29_io_out ? io_r_152_b : _GEN_6071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6073 = 8'h99 == r_count_29_io_out ? io_r_153_b : _GEN_6072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6074 = 8'h9a == r_count_29_io_out ? io_r_154_b : _GEN_6073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6075 = 8'h9b == r_count_29_io_out ? io_r_155_b : _GEN_6074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6076 = 8'h9c == r_count_29_io_out ? io_r_156_b : _GEN_6075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6077 = 8'h9d == r_count_29_io_out ? io_r_157_b : _GEN_6076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6078 = 8'h9e == r_count_29_io_out ? io_r_158_b : _GEN_6077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6079 = 8'h9f == r_count_29_io_out ? io_r_159_b : _GEN_6078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6080 = 8'ha0 == r_count_29_io_out ? io_r_160_b : _GEN_6079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6081 = 8'ha1 == r_count_29_io_out ? io_r_161_b : _GEN_6080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6082 = 8'ha2 == r_count_29_io_out ? io_r_162_b : _GEN_6081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6083 = 8'ha3 == r_count_29_io_out ? io_r_163_b : _GEN_6082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6084 = 8'ha4 == r_count_29_io_out ? io_r_164_b : _GEN_6083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6085 = 8'ha5 == r_count_29_io_out ? io_r_165_b : _GEN_6084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6086 = 8'ha6 == r_count_29_io_out ? io_r_166_b : _GEN_6085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6087 = 8'ha7 == r_count_29_io_out ? io_r_167_b : _GEN_6086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6088 = 8'ha8 == r_count_29_io_out ? io_r_168_b : _GEN_6087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6089 = 8'ha9 == r_count_29_io_out ? io_r_169_b : _GEN_6088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6090 = 8'haa == r_count_29_io_out ? io_r_170_b : _GEN_6089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6091 = 8'hab == r_count_29_io_out ? io_r_171_b : _GEN_6090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6092 = 8'hac == r_count_29_io_out ? io_r_172_b : _GEN_6091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6093 = 8'had == r_count_29_io_out ? io_r_173_b : _GEN_6092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6094 = 8'hae == r_count_29_io_out ? io_r_174_b : _GEN_6093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6095 = 8'haf == r_count_29_io_out ? io_r_175_b : _GEN_6094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6096 = 8'hb0 == r_count_29_io_out ? io_r_176_b : _GEN_6095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6097 = 8'hb1 == r_count_29_io_out ? io_r_177_b : _GEN_6096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6098 = 8'hb2 == r_count_29_io_out ? io_r_178_b : _GEN_6097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6099 = 8'hb3 == r_count_29_io_out ? io_r_179_b : _GEN_6098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6100 = 8'hb4 == r_count_29_io_out ? io_r_180_b : _GEN_6099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6101 = 8'hb5 == r_count_29_io_out ? io_r_181_b : _GEN_6100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6102 = 8'hb6 == r_count_29_io_out ? io_r_182_b : _GEN_6101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6103 = 8'hb7 == r_count_29_io_out ? io_r_183_b : _GEN_6102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6104 = 8'hb8 == r_count_29_io_out ? io_r_184_b : _GEN_6103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6105 = 8'hb9 == r_count_29_io_out ? io_r_185_b : _GEN_6104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6106 = 8'hba == r_count_29_io_out ? io_r_186_b : _GEN_6105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6107 = 8'hbb == r_count_29_io_out ? io_r_187_b : _GEN_6106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6108 = 8'hbc == r_count_29_io_out ? io_r_188_b : _GEN_6107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6109 = 8'hbd == r_count_29_io_out ? io_r_189_b : _GEN_6108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6110 = 8'hbe == r_count_29_io_out ? io_r_190_b : _GEN_6109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6111 = 8'hbf == r_count_29_io_out ? io_r_191_b : _GEN_6110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6112 = 8'hc0 == r_count_29_io_out ? io_r_192_b : _GEN_6111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6113 = 8'hc1 == r_count_29_io_out ? io_r_193_b : _GEN_6112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6114 = 8'hc2 == r_count_29_io_out ? io_r_194_b : _GEN_6113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6115 = 8'hc3 == r_count_29_io_out ? io_r_195_b : _GEN_6114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6116 = 8'hc4 == r_count_29_io_out ? io_r_196_b : _GEN_6115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6117 = 8'hc5 == r_count_29_io_out ? io_r_197_b : _GEN_6116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6118 = 8'hc6 == r_count_29_io_out ? io_r_198_b : _GEN_6117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6121 = 8'h1 == r_count_30_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6122 = 8'h2 == r_count_30_io_out ? io_r_2_b : _GEN_6121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6123 = 8'h3 == r_count_30_io_out ? io_r_3_b : _GEN_6122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6124 = 8'h4 == r_count_30_io_out ? io_r_4_b : _GEN_6123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6125 = 8'h5 == r_count_30_io_out ? io_r_5_b : _GEN_6124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6126 = 8'h6 == r_count_30_io_out ? io_r_6_b : _GEN_6125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6127 = 8'h7 == r_count_30_io_out ? io_r_7_b : _GEN_6126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6128 = 8'h8 == r_count_30_io_out ? io_r_8_b : _GEN_6127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6129 = 8'h9 == r_count_30_io_out ? io_r_9_b : _GEN_6128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6130 = 8'ha == r_count_30_io_out ? io_r_10_b : _GEN_6129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6131 = 8'hb == r_count_30_io_out ? io_r_11_b : _GEN_6130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6132 = 8'hc == r_count_30_io_out ? io_r_12_b : _GEN_6131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6133 = 8'hd == r_count_30_io_out ? io_r_13_b : _GEN_6132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6134 = 8'he == r_count_30_io_out ? io_r_14_b : _GEN_6133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6135 = 8'hf == r_count_30_io_out ? io_r_15_b : _GEN_6134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6136 = 8'h10 == r_count_30_io_out ? io_r_16_b : _GEN_6135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6137 = 8'h11 == r_count_30_io_out ? io_r_17_b : _GEN_6136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6138 = 8'h12 == r_count_30_io_out ? io_r_18_b : _GEN_6137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6139 = 8'h13 == r_count_30_io_out ? io_r_19_b : _GEN_6138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6140 = 8'h14 == r_count_30_io_out ? io_r_20_b : _GEN_6139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6141 = 8'h15 == r_count_30_io_out ? io_r_21_b : _GEN_6140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6142 = 8'h16 == r_count_30_io_out ? io_r_22_b : _GEN_6141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6143 = 8'h17 == r_count_30_io_out ? io_r_23_b : _GEN_6142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6144 = 8'h18 == r_count_30_io_out ? io_r_24_b : _GEN_6143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6145 = 8'h19 == r_count_30_io_out ? io_r_25_b : _GEN_6144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6146 = 8'h1a == r_count_30_io_out ? io_r_26_b : _GEN_6145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6147 = 8'h1b == r_count_30_io_out ? io_r_27_b : _GEN_6146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6148 = 8'h1c == r_count_30_io_out ? io_r_28_b : _GEN_6147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6149 = 8'h1d == r_count_30_io_out ? io_r_29_b : _GEN_6148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6150 = 8'h1e == r_count_30_io_out ? io_r_30_b : _GEN_6149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6151 = 8'h1f == r_count_30_io_out ? io_r_31_b : _GEN_6150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6152 = 8'h20 == r_count_30_io_out ? io_r_32_b : _GEN_6151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6153 = 8'h21 == r_count_30_io_out ? io_r_33_b : _GEN_6152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6154 = 8'h22 == r_count_30_io_out ? io_r_34_b : _GEN_6153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6155 = 8'h23 == r_count_30_io_out ? io_r_35_b : _GEN_6154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6156 = 8'h24 == r_count_30_io_out ? io_r_36_b : _GEN_6155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6157 = 8'h25 == r_count_30_io_out ? io_r_37_b : _GEN_6156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6158 = 8'h26 == r_count_30_io_out ? io_r_38_b : _GEN_6157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6159 = 8'h27 == r_count_30_io_out ? io_r_39_b : _GEN_6158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6160 = 8'h28 == r_count_30_io_out ? io_r_40_b : _GEN_6159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6161 = 8'h29 == r_count_30_io_out ? io_r_41_b : _GEN_6160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6162 = 8'h2a == r_count_30_io_out ? io_r_42_b : _GEN_6161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6163 = 8'h2b == r_count_30_io_out ? io_r_43_b : _GEN_6162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6164 = 8'h2c == r_count_30_io_out ? io_r_44_b : _GEN_6163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6165 = 8'h2d == r_count_30_io_out ? io_r_45_b : _GEN_6164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6166 = 8'h2e == r_count_30_io_out ? io_r_46_b : _GEN_6165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6167 = 8'h2f == r_count_30_io_out ? io_r_47_b : _GEN_6166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6168 = 8'h30 == r_count_30_io_out ? io_r_48_b : _GEN_6167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6169 = 8'h31 == r_count_30_io_out ? io_r_49_b : _GEN_6168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6170 = 8'h32 == r_count_30_io_out ? io_r_50_b : _GEN_6169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6171 = 8'h33 == r_count_30_io_out ? io_r_51_b : _GEN_6170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6172 = 8'h34 == r_count_30_io_out ? io_r_52_b : _GEN_6171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6173 = 8'h35 == r_count_30_io_out ? io_r_53_b : _GEN_6172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6174 = 8'h36 == r_count_30_io_out ? io_r_54_b : _GEN_6173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6175 = 8'h37 == r_count_30_io_out ? io_r_55_b : _GEN_6174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6176 = 8'h38 == r_count_30_io_out ? io_r_56_b : _GEN_6175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6177 = 8'h39 == r_count_30_io_out ? io_r_57_b : _GEN_6176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6178 = 8'h3a == r_count_30_io_out ? io_r_58_b : _GEN_6177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6179 = 8'h3b == r_count_30_io_out ? io_r_59_b : _GEN_6178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6180 = 8'h3c == r_count_30_io_out ? io_r_60_b : _GEN_6179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6181 = 8'h3d == r_count_30_io_out ? io_r_61_b : _GEN_6180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6182 = 8'h3e == r_count_30_io_out ? io_r_62_b : _GEN_6181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6183 = 8'h3f == r_count_30_io_out ? io_r_63_b : _GEN_6182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6184 = 8'h40 == r_count_30_io_out ? io_r_64_b : _GEN_6183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6185 = 8'h41 == r_count_30_io_out ? io_r_65_b : _GEN_6184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6186 = 8'h42 == r_count_30_io_out ? io_r_66_b : _GEN_6185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6187 = 8'h43 == r_count_30_io_out ? io_r_67_b : _GEN_6186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6188 = 8'h44 == r_count_30_io_out ? io_r_68_b : _GEN_6187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6189 = 8'h45 == r_count_30_io_out ? io_r_69_b : _GEN_6188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6190 = 8'h46 == r_count_30_io_out ? io_r_70_b : _GEN_6189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6191 = 8'h47 == r_count_30_io_out ? io_r_71_b : _GEN_6190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6192 = 8'h48 == r_count_30_io_out ? io_r_72_b : _GEN_6191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6193 = 8'h49 == r_count_30_io_out ? io_r_73_b : _GEN_6192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6194 = 8'h4a == r_count_30_io_out ? io_r_74_b : _GEN_6193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6195 = 8'h4b == r_count_30_io_out ? io_r_75_b : _GEN_6194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6196 = 8'h4c == r_count_30_io_out ? io_r_76_b : _GEN_6195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6197 = 8'h4d == r_count_30_io_out ? io_r_77_b : _GEN_6196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6198 = 8'h4e == r_count_30_io_out ? io_r_78_b : _GEN_6197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6199 = 8'h4f == r_count_30_io_out ? io_r_79_b : _GEN_6198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6200 = 8'h50 == r_count_30_io_out ? io_r_80_b : _GEN_6199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6201 = 8'h51 == r_count_30_io_out ? io_r_81_b : _GEN_6200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6202 = 8'h52 == r_count_30_io_out ? io_r_82_b : _GEN_6201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6203 = 8'h53 == r_count_30_io_out ? io_r_83_b : _GEN_6202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6204 = 8'h54 == r_count_30_io_out ? io_r_84_b : _GEN_6203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6205 = 8'h55 == r_count_30_io_out ? io_r_85_b : _GEN_6204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6206 = 8'h56 == r_count_30_io_out ? io_r_86_b : _GEN_6205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6207 = 8'h57 == r_count_30_io_out ? io_r_87_b : _GEN_6206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6208 = 8'h58 == r_count_30_io_out ? io_r_88_b : _GEN_6207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6209 = 8'h59 == r_count_30_io_out ? io_r_89_b : _GEN_6208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6210 = 8'h5a == r_count_30_io_out ? io_r_90_b : _GEN_6209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6211 = 8'h5b == r_count_30_io_out ? io_r_91_b : _GEN_6210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6212 = 8'h5c == r_count_30_io_out ? io_r_92_b : _GEN_6211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6213 = 8'h5d == r_count_30_io_out ? io_r_93_b : _GEN_6212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6214 = 8'h5e == r_count_30_io_out ? io_r_94_b : _GEN_6213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6215 = 8'h5f == r_count_30_io_out ? io_r_95_b : _GEN_6214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6216 = 8'h60 == r_count_30_io_out ? io_r_96_b : _GEN_6215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6217 = 8'h61 == r_count_30_io_out ? io_r_97_b : _GEN_6216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6218 = 8'h62 == r_count_30_io_out ? io_r_98_b : _GEN_6217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6219 = 8'h63 == r_count_30_io_out ? io_r_99_b : _GEN_6218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6220 = 8'h64 == r_count_30_io_out ? io_r_100_b : _GEN_6219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6221 = 8'h65 == r_count_30_io_out ? io_r_101_b : _GEN_6220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6222 = 8'h66 == r_count_30_io_out ? io_r_102_b : _GEN_6221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6223 = 8'h67 == r_count_30_io_out ? io_r_103_b : _GEN_6222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6224 = 8'h68 == r_count_30_io_out ? io_r_104_b : _GEN_6223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6225 = 8'h69 == r_count_30_io_out ? io_r_105_b : _GEN_6224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6226 = 8'h6a == r_count_30_io_out ? io_r_106_b : _GEN_6225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6227 = 8'h6b == r_count_30_io_out ? io_r_107_b : _GEN_6226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6228 = 8'h6c == r_count_30_io_out ? io_r_108_b : _GEN_6227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6229 = 8'h6d == r_count_30_io_out ? io_r_109_b : _GEN_6228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6230 = 8'h6e == r_count_30_io_out ? io_r_110_b : _GEN_6229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6231 = 8'h6f == r_count_30_io_out ? io_r_111_b : _GEN_6230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6232 = 8'h70 == r_count_30_io_out ? io_r_112_b : _GEN_6231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6233 = 8'h71 == r_count_30_io_out ? io_r_113_b : _GEN_6232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6234 = 8'h72 == r_count_30_io_out ? io_r_114_b : _GEN_6233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6235 = 8'h73 == r_count_30_io_out ? io_r_115_b : _GEN_6234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6236 = 8'h74 == r_count_30_io_out ? io_r_116_b : _GEN_6235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6237 = 8'h75 == r_count_30_io_out ? io_r_117_b : _GEN_6236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6238 = 8'h76 == r_count_30_io_out ? io_r_118_b : _GEN_6237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6239 = 8'h77 == r_count_30_io_out ? io_r_119_b : _GEN_6238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6240 = 8'h78 == r_count_30_io_out ? io_r_120_b : _GEN_6239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6241 = 8'h79 == r_count_30_io_out ? io_r_121_b : _GEN_6240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6242 = 8'h7a == r_count_30_io_out ? io_r_122_b : _GEN_6241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6243 = 8'h7b == r_count_30_io_out ? io_r_123_b : _GEN_6242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6244 = 8'h7c == r_count_30_io_out ? io_r_124_b : _GEN_6243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6245 = 8'h7d == r_count_30_io_out ? io_r_125_b : _GEN_6244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6246 = 8'h7e == r_count_30_io_out ? io_r_126_b : _GEN_6245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6247 = 8'h7f == r_count_30_io_out ? io_r_127_b : _GEN_6246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6248 = 8'h80 == r_count_30_io_out ? io_r_128_b : _GEN_6247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6249 = 8'h81 == r_count_30_io_out ? io_r_129_b : _GEN_6248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6250 = 8'h82 == r_count_30_io_out ? io_r_130_b : _GEN_6249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6251 = 8'h83 == r_count_30_io_out ? io_r_131_b : _GEN_6250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6252 = 8'h84 == r_count_30_io_out ? io_r_132_b : _GEN_6251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6253 = 8'h85 == r_count_30_io_out ? io_r_133_b : _GEN_6252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6254 = 8'h86 == r_count_30_io_out ? io_r_134_b : _GEN_6253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6255 = 8'h87 == r_count_30_io_out ? io_r_135_b : _GEN_6254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6256 = 8'h88 == r_count_30_io_out ? io_r_136_b : _GEN_6255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6257 = 8'h89 == r_count_30_io_out ? io_r_137_b : _GEN_6256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6258 = 8'h8a == r_count_30_io_out ? io_r_138_b : _GEN_6257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6259 = 8'h8b == r_count_30_io_out ? io_r_139_b : _GEN_6258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6260 = 8'h8c == r_count_30_io_out ? io_r_140_b : _GEN_6259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6261 = 8'h8d == r_count_30_io_out ? io_r_141_b : _GEN_6260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6262 = 8'h8e == r_count_30_io_out ? io_r_142_b : _GEN_6261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6263 = 8'h8f == r_count_30_io_out ? io_r_143_b : _GEN_6262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6264 = 8'h90 == r_count_30_io_out ? io_r_144_b : _GEN_6263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6265 = 8'h91 == r_count_30_io_out ? io_r_145_b : _GEN_6264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6266 = 8'h92 == r_count_30_io_out ? io_r_146_b : _GEN_6265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6267 = 8'h93 == r_count_30_io_out ? io_r_147_b : _GEN_6266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6268 = 8'h94 == r_count_30_io_out ? io_r_148_b : _GEN_6267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6269 = 8'h95 == r_count_30_io_out ? io_r_149_b : _GEN_6268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6270 = 8'h96 == r_count_30_io_out ? io_r_150_b : _GEN_6269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6271 = 8'h97 == r_count_30_io_out ? io_r_151_b : _GEN_6270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6272 = 8'h98 == r_count_30_io_out ? io_r_152_b : _GEN_6271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6273 = 8'h99 == r_count_30_io_out ? io_r_153_b : _GEN_6272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6274 = 8'h9a == r_count_30_io_out ? io_r_154_b : _GEN_6273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6275 = 8'h9b == r_count_30_io_out ? io_r_155_b : _GEN_6274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6276 = 8'h9c == r_count_30_io_out ? io_r_156_b : _GEN_6275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6277 = 8'h9d == r_count_30_io_out ? io_r_157_b : _GEN_6276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6278 = 8'h9e == r_count_30_io_out ? io_r_158_b : _GEN_6277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6279 = 8'h9f == r_count_30_io_out ? io_r_159_b : _GEN_6278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6280 = 8'ha0 == r_count_30_io_out ? io_r_160_b : _GEN_6279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6281 = 8'ha1 == r_count_30_io_out ? io_r_161_b : _GEN_6280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6282 = 8'ha2 == r_count_30_io_out ? io_r_162_b : _GEN_6281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6283 = 8'ha3 == r_count_30_io_out ? io_r_163_b : _GEN_6282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6284 = 8'ha4 == r_count_30_io_out ? io_r_164_b : _GEN_6283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6285 = 8'ha5 == r_count_30_io_out ? io_r_165_b : _GEN_6284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6286 = 8'ha6 == r_count_30_io_out ? io_r_166_b : _GEN_6285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6287 = 8'ha7 == r_count_30_io_out ? io_r_167_b : _GEN_6286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6288 = 8'ha8 == r_count_30_io_out ? io_r_168_b : _GEN_6287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6289 = 8'ha9 == r_count_30_io_out ? io_r_169_b : _GEN_6288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6290 = 8'haa == r_count_30_io_out ? io_r_170_b : _GEN_6289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6291 = 8'hab == r_count_30_io_out ? io_r_171_b : _GEN_6290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6292 = 8'hac == r_count_30_io_out ? io_r_172_b : _GEN_6291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6293 = 8'had == r_count_30_io_out ? io_r_173_b : _GEN_6292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6294 = 8'hae == r_count_30_io_out ? io_r_174_b : _GEN_6293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6295 = 8'haf == r_count_30_io_out ? io_r_175_b : _GEN_6294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6296 = 8'hb0 == r_count_30_io_out ? io_r_176_b : _GEN_6295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6297 = 8'hb1 == r_count_30_io_out ? io_r_177_b : _GEN_6296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6298 = 8'hb2 == r_count_30_io_out ? io_r_178_b : _GEN_6297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6299 = 8'hb3 == r_count_30_io_out ? io_r_179_b : _GEN_6298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6300 = 8'hb4 == r_count_30_io_out ? io_r_180_b : _GEN_6299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6301 = 8'hb5 == r_count_30_io_out ? io_r_181_b : _GEN_6300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6302 = 8'hb6 == r_count_30_io_out ? io_r_182_b : _GEN_6301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6303 = 8'hb7 == r_count_30_io_out ? io_r_183_b : _GEN_6302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6304 = 8'hb8 == r_count_30_io_out ? io_r_184_b : _GEN_6303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6305 = 8'hb9 == r_count_30_io_out ? io_r_185_b : _GEN_6304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6306 = 8'hba == r_count_30_io_out ? io_r_186_b : _GEN_6305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6307 = 8'hbb == r_count_30_io_out ? io_r_187_b : _GEN_6306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6308 = 8'hbc == r_count_30_io_out ? io_r_188_b : _GEN_6307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6309 = 8'hbd == r_count_30_io_out ? io_r_189_b : _GEN_6308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6310 = 8'hbe == r_count_30_io_out ? io_r_190_b : _GEN_6309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6311 = 8'hbf == r_count_30_io_out ? io_r_191_b : _GEN_6310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6312 = 8'hc0 == r_count_30_io_out ? io_r_192_b : _GEN_6311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6313 = 8'hc1 == r_count_30_io_out ? io_r_193_b : _GEN_6312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6314 = 8'hc2 == r_count_30_io_out ? io_r_194_b : _GEN_6313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6315 = 8'hc3 == r_count_30_io_out ? io_r_195_b : _GEN_6314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6316 = 8'hc4 == r_count_30_io_out ? io_r_196_b : _GEN_6315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6317 = 8'hc5 == r_count_30_io_out ? io_r_197_b : _GEN_6316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6318 = 8'hc6 == r_count_30_io_out ? io_r_198_b : _GEN_6317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6321 = 8'h1 == r_count_31_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6322 = 8'h2 == r_count_31_io_out ? io_r_2_b : _GEN_6321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6323 = 8'h3 == r_count_31_io_out ? io_r_3_b : _GEN_6322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6324 = 8'h4 == r_count_31_io_out ? io_r_4_b : _GEN_6323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6325 = 8'h5 == r_count_31_io_out ? io_r_5_b : _GEN_6324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6326 = 8'h6 == r_count_31_io_out ? io_r_6_b : _GEN_6325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6327 = 8'h7 == r_count_31_io_out ? io_r_7_b : _GEN_6326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6328 = 8'h8 == r_count_31_io_out ? io_r_8_b : _GEN_6327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6329 = 8'h9 == r_count_31_io_out ? io_r_9_b : _GEN_6328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6330 = 8'ha == r_count_31_io_out ? io_r_10_b : _GEN_6329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6331 = 8'hb == r_count_31_io_out ? io_r_11_b : _GEN_6330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6332 = 8'hc == r_count_31_io_out ? io_r_12_b : _GEN_6331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6333 = 8'hd == r_count_31_io_out ? io_r_13_b : _GEN_6332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6334 = 8'he == r_count_31_io_out ? io_r_14_b : _GEN_6333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6335 = 8'hf == r_count_31_io_out ? io_r_15_b : _GEN_6334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6336 = 8'h10 == r_count_31_io_out ? io_r_16_b : _GEN_6335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6337 = 8'h11 == r_count_31_io_out ? io_r_17_b : _GEN_6336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6338 = 8'h12 == r_count_31_io_out ? io_r_18_b : _GEN_6337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6339 = 8'h13 == r_count_31_io_out ? io_r_19_b : _GEN_6338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6340 = 8'h14 == r_count_31_io_out ? io_r_20_b : _GEN_6339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6341 = 8'h15 == r_count_31_io_out ? io_r_21_b : _GEN_6340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6342 = 8'h16 == r_count_31_io_out ? io_r_22_b : _GEN_6341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6343 = 8'h17 == r_count_31_io_out ? io_r_23_b : _GEN_6342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6344 = 8'h18 == r_count_31_io_out ? io_r_24_b : _GEN_6343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6345 = 8'h19 == r_count_31_io_out ? io_r_25_b : _GEN_6344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6346 = 8'h1a == r_count_31_io_out ? io_r_26_b : _GEN_6345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6347 = 8'h1b == r_count_31_io_out ? io_r_27_b : _GEN_6346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6348 = 8'h1c == r_count_31_io_out ? io_r_28_b : _GEN_6347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6349 = 8'h1d == r_count_31_io_out ? io_r_29_b : _GEN_6348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6350 = 8'h1e == r_count_31_io_out ? io_r_30_b : _GEN_6349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6351 = 8'h1f == r_count_31_io_out ? io_r_31_b : _GEN_6350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6352 = 8'h20 == r_count_31_io_out ? io_r_32_b : _GEN_6351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6353 = 8'h21 == r_count_31_io_out ? io_r_33_b : _GEN_6352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6354 = 8'h22 == r_count_31_io_out ? io_r_34_b : _GEN_6353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6355 = 8'h23 == r_count_31_io_out ? io_r_35_b : _GEN_6354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6356 = 8'h24 == r_count_31_io_out ? io_r_36_b : _GEN_6355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6357 = 8'h25 == r_count_31_io_out ? io_r_37_b : _GEN_6356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6358 = 8'h26 == r_count_31_io_out ? io_r_38_b : _GEN_6357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6359 = 8'h27 == r_count_31_io_out ? io_r_39_b : _GEN_6358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6360 = 8'h28 == r_count_31_io_out ? io_r_40_b : _GEN_6359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6361 = 8'h29 == r_count_31_io_out ? io_r_41_b : _GEN_6360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6362 = 8'h2a == r_count_31_io_out ? io_r_42_b : _GEN_6361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6363 = 8'h2b == r_count_31_io_out ? io_r_43_b : _GEN_6362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6364 = 8'h2c == r_count_31_io_out ? io_r_44_b : _GEN_6363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6365 = 8'h2d == r_count_31_io_out ? io_r_45_b : _GEN_6364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6366 = 8'h2e == r_count_31_io_out ? io_r_46_b : _GEN_6365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6367 = 8'h2f == r_count_31_io_out ? io_r_47_b : _GEN_6366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6368 = 8'h30 == r_count_31_io_out ? io_r_48_b : _GEN_6367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6369 = 8'h31 == r_count_31_io_out ? io_r_49_b : _GEN_6368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6370 = 8'h32 == r_count_31_io_out ? io_r_50_b : _GEN_6369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6371 = 8'h33 == r_count_31_io_out ? io_r_51_b : _GEN_6370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6372 = 8'h34 == r_count_31_io_out ? io_r_52_b : _GEN_6371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6373 = 8'h35 == r_count_31_io_out ? io_r_53_b : _GEN_6372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6374 = 8'h36 == r_count_31_io_out ? io_r_54_b : _GEN_6373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6375 = 8'h37 == r_count_31_io_out ? io_r_55_b : _GEN_6374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6376 = 8'h38 == r_count_31_io_out ? io_r_56_b : _GEN_6375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6377 = 8'h39 == r_count_31_io_out ? io_r_57_b : _GEN_6376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6378 = 8'h3a == r_count_31_io_out ? io_r_58_b : _GEN_6377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6379 = 8'h3b == r_count_31_io_out ? io_r_59_b : _GEN_6378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6380 = 8'h3c == r_count_31_io_out ? io_r_60_b : _GEN_6379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6381 = 8'h3d == r_count_31_io_out ? io_r_61_b : _GEN_6380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6382 = 8'h3e == r_count_31_io_out ? io_r_62_b : _GEN_6381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6383 = 8'h3f == r_count_31_io_out ? io_r_63_b : _GEN_6382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6384 = 8'h40 == r_count_31_io_out ? io_r_64_b : _GEN_6383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6385 = 8'h41 == r_count_31_io_out ? io_r_65_b : _GEN_6384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6386 = 8'h42 == r_count_31_io_out ? io_r_66_b : _GEN_6385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6387 = 8'h43 == r_count_31_io_out ? io_r_67_b : _GEN_6386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6388 = 8'h44 == r_count_31_io_out ? io_r_68_b : _GEN_6387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6389 = 8'h45 == r_count_31_io_out ? io_r_69_b : _GEN_6388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6390 = 8'h46 == r_count_31_io_out ? io_r_70_b : _GEN_6389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6391 = 8'h47 == r_count_31_io_out ? io_r_71_b : _GEN_6390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6392 = 8'h48 == r_count_31_io_out ? io_r_72_b : _GEN_6391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6393 = 8'h49 == r_count_31_io_out ? io_r_73_b : _GEN_6392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6394 = 8'h4a == r_count_31_io_out ? io_r_74_b : _GEN_6393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6395 = 8'h4b == r_count_31_io_out ? io_r_75_b : _GEN_6394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6396 = 8'h4c == r_count_31_io_out ? io_r_76_b : _GEN_6395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6397 = 8'h4d == r_count_31_io_out ? io_r_77_b : _GEN_6396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6398 = 8'h4e == r_count_31_io_out ? io_r_78_b : _GEN_6397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6399 = 8'h4f == r_count_31_io_out ? io_r_79_b : _GEN_6398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6400 = 8'h50 == r_count_31_io_out ? io_r_80_b : _GEN_6399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6401 = 8'h51 == r_count_31_io_out ? io_r_81_b : _GEN_6400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6402 = 8'h52 == r_count_31_io_out ? io_r_82_b : _GEN_6401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6403 = 8'h53 == r_count_31_io_out ? io_r_83_b : _GEN_6402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6404 = 8'h54 == r_count_31_io_out ? io_r_84_b : _GEN_6403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6405 = 8'h55 == r_count_31_io_out ? io_r_85_b : _GEN_6404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6406 = 8'h56 == r_count_31_io_out ? io_r_86_b : _GEN_6405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6407 = 8'h57 == r_count_31_io_out ? io_r_87_b : _GEN_6406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6408 = 8'h58 == r_count_31_io_out ? io_r_88_b : _GEN_6407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6409 = 8'h59 == r_count_31_io_out ? io_r_89_b : _GEN_6408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6410 = 8'h5a == r_count_31_io_out ? io_r_90_b : _GEN_6409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6411 = 8'h5b == r_count_31_io_out ? io_r_91_b : _GEN_6410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6412 = 8'h5c == r_count_31_io_out ? io_r_92_b : _GEN_6411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6413 = 8'h5d == r_count_31_io_out ? io_r_93_b : _GEN_6412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6414 = 8'h5e == r_count_31_io_out ? io_r_94_b : _GEN_6413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6415 = 8'h5f == r_count_31_io_out ? io_r_95_b : _GEN_6414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6416 = 8'h60 == r_count_31_io_out ? io_r_96_b : _GEN_6415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6417 = 8'h61 == r_count_31_io_out ? io_r_97_b : _GEN_6416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6418 = 8'h62 == r_count_31_io_out ? io_r_98_b : _GEN_6417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6419 = 8'h63 == r_count_31_io_out ? io_r_99_b : _GEN_6418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6420 = 8'h64 == r_count_31_io_out ? io_r_100_b : _GEN_6419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6421 = 8'h65 == r_count_31_io_out ? io_r_101_b : _GEN_6420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6422 = 8'h66 == r_count_31_io_out ? io_r_102_b : _GEN_6421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6423 = 8'h67 == r_count_31_io_out ? io_r_103_b : _GEN_6422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6424 = 8'h68 == r_count_31_io_out ? io_r_104_b : _GEN_6423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6425 = 8'h69 == r_count_31_io_out ? io_r_105_b : _GEN_6424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6426 = 8'h6a == r_count_31_io_out ? io_r_106_b : _GEN_6425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6427 = 8'h6b == r_count_31_io_out ? io_r_107_b : _GEN_6426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6428 = 8'h6c == r_count_31_io_out ? io_r_108_b : _GEN_6427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6429 = 8'h6d == r_count_31_io_out ? io_r_109_b : _GEN_6428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6430 = 8'h6e == r_count_31_io_out ? io_r_110_b : _GEN_6429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6431 = 8'h6f == r_count_31_io_out ? io_r_111_b : _GEN_6430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6432 = 8'h70 == r_count_31_io_out ? io_r_112_b : _GEN_6431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6433 = 8'h71 == r_count_31_io_out ? io_r_113_b : _GEN_6432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6434 = 8'h72 == r_count_31_io_out ? io_r_114_b : _GEN_6433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6435 = 8'h73 == r_count_31_io_out ? io_r_115_b : _GEN_6434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6436 = 8'h74 == r_count_31_io_out ? io_r_116_b : _GEN_6435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6437 = 8'h75 == r_count_31_io_out ? io_r_117_b : _GEN_6436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6438 = 8'h76 == r_count_31_io_out ? io_r_118_b : _GEN_6437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6439 = 8'h77 == r_count_31_io_out ? io_r_119_b : _GEN_6438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6440 = 8'h78 == r_count_31_io_out ? io_r_120_b : _GEN_6439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6441 = 8'h79 == r_count_31_io_out ? io_r_121_b : _GEN_6440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6442 = 8'h7a == r_count_31_io_out ? io_r_122_b : _GEN_6441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6443 = 8'h7b == r_count_31_io_out ? io_r_123_b : _GEN_6442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6444 = 8'h7c == r_count_31_io_out ? io_r_124_b : _GEN_6443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6445 = 8'h7d == r_count_31_io_out ? io_r_125_b : _GEN_6444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6446 = 8'h7e == r_count_31_io_out ? io_r_126_b : _GEN_6445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6447 = 8'h7f == r_count_31_io_out ? io_r_127_b : _GEN_6446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6448 = 8'h80 == r_count_31_io_out ? io_r_128_b : _GEN_6447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6449 = 8'h81 == r_count_31_io_out ? io_r_129_b : _GEN_6448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6450 = 8'h82 == r_count_31_io_out ? io_r_130_b : _GEN_6449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6451 = 8'h83 == r_count_31_io_out ? io_r_131_b : _GEN_6450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6452 = 8'h84 == r_count_31_io_out ? io_r_132_b : _GEN_6451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6453 = 8'h85 == r_count_31_io_out ? io_r_133_b : _GEN_6452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6454 = 8'h86 == r_count_31_io_out ? io_r_134_b : _GEN_6453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6455 = 8'h87 == r_count_31_io_out ? io_r_135_b : _GEN_6454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6456 = 8'h88 == r_count_31_io_out ? io_r_136_b : _GEN_6455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6457 = 8'h89 == r_count_31_io_out ? io_r_137_b : _GEN_6456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6458 = 8'h8a == r_count_31_io_out ? io_r_138_b : _GEN_6457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6459 = 8'h8b == r_count_31_io_out ? io_r_139_b : _GEN_6458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6460 = 8'h8c == r_count_31_io_out ? io_r_140_b : _GEN_6459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6461 = 8'h8d == r_count_31_io_out ? io_r_141_b : _GEN_6460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6462 = 8'h8e == r_count_31_io_out ? io_r_142_b : _GEN_6461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6463 = 8'h8f == r_count_31_io_out ? io_r_143_b : _GEN_6462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6464 = 8'h90 == r_count_31_io_out ? io_r_144_b : _GEN_6463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6465 = 8'h91 == r_count_31_io_out ? io_r_145_b : _GEN_6464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6466 = 8'h92 == r_count_31_io_out ? io_r_146_b : _GEN_6465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6467 = 8'h93 == r_count_31_io_out ? io_r_147_b : _GEN_6466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6468 = 8'h94 == r_count_31_io_out ? io_r_148_b : _GEN_6467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6469 = 8'h95 == r_count_31_io_out ? io_r_149_b : _GEN_6468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6470 = 8'h96 == r_count_31_io_out ? io_r_150_b : _GEN_6469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6471 = 8'h97 == r_count_31_io_out ? io_r_151_b : _GEN_6470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6472 = 8'h98 == r_count_31_io_out ? io_r_152_b : _GEN_6471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6473 = 8'h99 == r_count_31_io_out ? io_r_153_b : _GEN_6472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6474 = 8'h9a == r_count_31_io_out ? io_r_154_b : _GEN_6473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6475 = 8'h9b == r_count_31_io_out ? io_r_155_b : _GEN_6474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6476 = 8'h9c == r_count_31_io_out ? io_r_156_b : _GEN_6475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6477 = 8'h9d == r_count_31_io_out ? io_r_157_b : _GEN_6476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6478 = 8'h9e == r_count_31_io_out ? io_r_158_b : _GEN_6477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6479 = 8'h9f == r_count_31_io_out ? io_r_159_b : _GEN_6478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6480 = 8'ha0 == r_count_31_io_out ? io_r_160_b : _GEN_6479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6481 = 8'ha1 == r_count_31_io_out ? io_r_161_b : _GEN_6480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6482 = 8'ha2 == r_count_31_io_out ? io_r_162_b : _GEN_6481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6483 = 8'ha3 == r_count_31_io_out ? io_r_163_b : _GEN_6482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6484 = 8'ha4 == r_count_31_io_out ? io_r_164_b : _GEN_6483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6485 = 8'ha5 == r_count_31_io_out ? io_r_165_b : _GEN_6484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6486 = 8'ha6 == r_count_31_io_out ? io_r_166_b : _GEN_6485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6487 = 8'ha7 == r_count_31_io_out ? io_r_167_b : _GEN_6486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6488 = 8'ha8 == r_count_31_io_out ? io_r_168_b : _GEN_6487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6489 = 8'ha9 == r_count_31_io_out ? io_r_169_b : _GEN_6488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6490 = 8'haa == r_count_31_io_out ? io_r_170_b : _GEN_6489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6491 = 8'hab == r_count_31_io_out ? io_r_171_b : _GEN_6490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6492 = 8'hac == r_count_31_io_out ? io_r_172_b : _GEN_6491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6493 = 8'had == r_count_31_io_out ? io_r_173_b : _GEN_6492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6494 = 8'hae == r_count_31_io_out ? io_r_174_b : _GEN_6493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6495 = 8'haf == r_count_31_io_out ? io_r_175_b : _GEN_6494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6496 = 8'hb0 == r_count_31_io_out ? io_r_176_b : _GEN_6495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6497 = 8'hb1 == r_count_31_io_out ? io_r_177_b : _GEN_6496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6498 = 8'hb2 == r_count_31_io_out ? io_r_178_b : _GEN_6497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6499 = 8'hb3 == r_count_31_io_out ? io_r_179_b : _GEN_6498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6500 = 8'hb4 == r_count_31_io_out ? io_r_180_b : _GEN_6499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6501 = 8'hb5 == r_count_31_io_out ? io_r_181_b : _GEN_6500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6502 = 8'hb6 == r_count_31_io_out ? io_r_182_b : _GEN_6501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6503 = 8'hb7 == r_count_31_io_out ? io_r_183_b : _GEN_6502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6504 = 8'hb8 == r_count_31_io_out ? io_r_184_b : _GEN_6503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6505 = 8'hb9 == r_count_31_io_out ? io_r_185_b : _GEN_6504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6506 = 8'hba == r_count_31_io_out ? io_r_186_b : _GEN_6505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6507 = 8'hbb == r_count_31_io_out ? io_r_187_b : _GEN_6506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6508 = 8'hbc == r_count_31_io_out ? io_r_188_b : _GEN_6507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6509 = 8'hbd == r_count_31_io_out ? io_r_189_b : _GEN_6508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6510 = 8'hbe == r_count_31_io_out ? io_r_190_b : _GEN_6509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6511 = 8'hbf == r_count_31_io_out ? io_r_191_b : _GEN_6510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6512 = 8'hc0 == r_count_31_io_out ? io_r_192_b : _GEN_6511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6513 = 8'hc1 == r_count_31_io_out ? io_r_193_b : _GEN_6512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6514 = 8'hc2 == r_count_31_io_out ? io_r_194_b : _GEN_6513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6515 = 8'hc3 == r_count_31_io_out ? io_r_195_b : _GEN_6514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6516 = 8'hc4 == r_count_31_io_out ? io_r_196_b : _GEN_6515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6517 = 8'hc5 == r_count_31_io_out ? io_r_197_b : _GEN_6516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6518 = 8'hc6 == r_count_31_io_out ? io_r_198_b : _GEN_6517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6521 = 8'h1 == r_count_32_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6522 = 8'h2 == r_count_32_io_out ? io_r_2_b : _GEN_6521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6523 = 8'h3 == r_count_32_io_out ? io_r_3_b : _GEN_6522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6524 = 8'h4 == r_count_32_io_out ? io_r_4_b : _GEN_6523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6525 = 8'h5 == r_count_32_io_out ? io_r_5_b : _GEN_6524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6526 = 8'h6 == r_count_32_io_out ? io_r_6_b : _GEN_6525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6527 = 8'h7 == r_count_32_io_out ? io_r_7_b : _GEN_6526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6528 = 8'h8 == r_count_32_io_out ? io_r_8_b : _GEN_6527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6529 = 8'h9 == r_count_32_io_out ? io_r_9_b : _GEN_6528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6530 = 8'ha == r_count_32_io_out ? io_r_10_b : _GEN_6529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6531 = 8'hb == r_count_32_io_out ? io_r_11_b : _GEN_6530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6532 = 8'hc == r_count_32_io_out ? io_r_12_b : _GEN_6531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6533 = 8'hd == r_count_32_io_out ? io_r_13_b : _GEN_6532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6534 = 8'he == r_count_32_io_out ? io_r_14_b : _GEN_6533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6535 = 8'hf == r_count_32_io_out ? io_r_15_b : _GEN_6534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6536 = 8'h10 == r_count_32_io_out ? io_r_16_b : _GEN_6535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6537 = 8'h11 == r_count_32_io_out ? io_r_17_b : _GEN_6536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6538 = 8'h12 == r_count_32_io_out ? io_r_18_b : _GEN_6537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6539 = 8'h13 == r_count_32_io_out ? io_r_19_b : _GEN_6538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6540 = 8'h14 == r_count_32_io_out ? io_r_20_b : _GEN_6539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6541 = 8'h15 == r_count_32_io_out ? io_r_21_b : _GEN_6540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6542 = 8'h16 == r_count_32_io_out ? io_r_22_b : _GEN_6541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6543 = 8'h17 == r_count_32_io_out ? io_r_23_b : _GEN_6542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6544 = 8'h18 == r_count_32_io_out ? io_r_24_b : _GEN_6543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6545 = 8'h19 == r_count_32_io_out ? io_r_25_b : _GEN_6544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6546 = 8'h1a == r_count_32_io_out ? io_r_26_b : _GEN_6545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6547 = 8'h1b == r_count_32_io_out ? io_r_27_b : _GEN_6546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6548 = 8'h1c == r_count_32_io_out ? io_r_28_b : _GEN_6547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6549 = 8'h1d == r_count_32_io_out ? io_r_29_b : _GEN_6548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6550 = 8'h1e == r_count_32_io_out ? io_r_30_b : _GEN_6549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6551 = 8'h1f == r_count_32_io_out ? io_r_31_b : _GEN_6550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6552 = 8'h20 == r_count_32_io_out ? io_r_32_b : _GEN_6551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6553 = 8'h21 == r_count_32_io_out ? io_r_33_b : _GEN_6552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6554 = 8'h22 == r_count_32_io_out ? io_r_34_b : _GEN_6553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6555 = 8'h23 == r_count_32_io_out ? io_r_35_b : _GEN_6554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6556 = 8'h24 == r_count_32_io_out ? io_r_36_b : _GEN_6555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6557 = 8'h25 == r_count_32_io_out ? io_r_37_b : _GEN_6556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6558 = 8'h26 == r_count_32_io_out ? io_r_38_b : _GEN_6557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6559 = 8'h27 == r_count_32_io_out ? io_r_39_b : _GEN_6558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6560 = 8'h28 == r_count_32_io_out ? io_r_40_b : _GEN_6559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6561 = 8'h29 == r_count_32_io_out ? io_r_41_b : _GEN_6560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6562 = 8'h2a == r_count_32_io_out ? io_r_42_b : _GEN_6561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6563 = 8'h2b == r_count_32_io_out ? io_r_43_b : _GEN_6562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6564 = 8'h2c == r_count_32_io_out ? io_r_44_b : _GEN_6563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6565 = 8'h2d == r_count_32_io_out ? io_r_45_b : _GEN_6564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6566 = 8'h2e == r_count_32_io_out ? io_r_46_b : _GEN_6565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6567 = 8'h2f == r_count_32_io_out ? io_r_47_b : _GEN_6566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6568 = 8'h30 == r_count_32_io_out ? io_r_48_b : _GEN_6567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6569 = 8'h31 == r_count_32_io_out ? io_r_49_b : _GEN_6568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6570 = 8'h32 == r_count_32_io_out ? io_r_50_b : _GEN_6569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6571 = 8'h33 == r_count_32_io_out ? io_r_51_b : _GEN_6570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6572 = 8'h34 == r_count_32_io_out ? io_r_52_b : _GEN_6571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6573 = 8'h35 == r_count_32_io_out ? io_r_53_b : _GEN_6572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6574 = 8'h36 == r_count_32_io_out ? io_r_54_b : _GEN_6573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6575 = 8'h37 == r_count_32_io_out ? io_r_55_b : _GEN_6574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6576 = 8'h38 == r_count_32_io_out ? io_r_56_b : _GEN_6575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6577 = 8'h39 == r_count_32_io_out ? io_r_57_b : _GEN_6576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6578 = 8'h3a == r_count_32_io_out ? io_r_58_b : _GEN_6577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6579 = 8'h3b == r_count_32_io_out ? io_r_59_b : _GEN_6578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6580 = 8'h3c == r_count_32_io_out ? io_r_60_b : _GEN_6579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6581 = 8'h3d == r_count_32_io_out ? io_r_61_b : _GEN_6580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6582 = 8'h3e == r_count_32_io_out ? io_r_62_b : _GEN_6581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6583 = 8'h3f == r_count_32_io_out ? io_r_63_b : _GEN_6582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6584 = 8'h40 == r_count_32_io_out ? io_r_64_b : _GEN_6583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6585 = 8'h41 == r_count_32_io_out ? io_r_65_b : _GEN_6584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6586 = 8'h42 == r_count_32_io_out ? io_r_66_b : _GEN_6585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6587 = 8'h43 == r_count_32_io_out ? io_r_67_b : _GEN_6586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6588 = 8'h44 == r_count_32_io_out ? io_r_68_b : _GEN_6587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6589 = 8'h45 == r_count_32_io_out ? io_r_69_b : _GEN_6588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6590 = 8'h46 == r_count_32_io_out ? io_r_70_b : _GEN_6589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6591 = 8'h47 == r_count_32_io_out ? io_r_71_b : _GEN_6590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6592 = 8'h48 == r_count_32_io_out ? io_r_72_b : _GEN_6591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6593 = 8'h49 == r_count_32_io_out ? io_r_73_b : _GEN_6592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6594 = 8'h4a == r_count_32_io_out ? io_r_74_b : _GEN_6593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6595 = 8'h4b == r_count_32_io_out ? io_r_75_b : _GEN_6594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6596 = 8'h4c == r_count_32_io_out ? io_r_76_b : _GEN_6595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6597 = 8'h4d == r_count_32_io_out ? io_r_77_b : _GEN_6596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6598 = 8'h4e == r_count_32_io_out ? io_r_78_b : _GEN_6597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6599 = 8'h4f == r_count_32_io_out ? io_r_79_b : _GEN_6598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6600 = 8'h50 == r_count_32_io_out ? io_r_80_b : _GEN_6599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6601 = 8'h51 == r_count_32_io_out ? io_r_81_b : _GEN_6600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6602 = 8'h52 == r_count_32_io_out ? io_r_82_b : _GEN_6601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6603 = 8'h53 == r_count_32_io_out ? io_r_83_b : _GEN_6602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6604 = 8'h54 == r_count_32_io_out ? io_r_84_b : _GEN_6603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6605 = 8'h55 == r_count_32_io_out ? io_r_85_b : _GEN_6604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6606 = 8'h56 == r_count_32_io_out ? io_r_86_b : _GEN_6605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6607 = 8'h57 == r_count_32_io_out ? io_r_87_b : _GEN_6606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6608 = 8'h58 == r_count_32_io_out ? io_r_88_b : _GEN_6607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6609 = 8'h59 == r_count_32_io_out ? io_r_89_b : _GEN_6608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6610 = 8'h5a == r_count_32_io_out ? io_r_90_b : _GEN_6609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6611 = 8'h5b == r_count_32_io_out ? io_r_91_b : _GEN_6610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6612 = 8'h5c == r_count_32_io_out ? io_r_92_b : _GEN_6611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6613 = 8'h5d == r_count_32_io_out ? io_r_93_b : _GEN_6612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6614 = 8'h5e == r_count_32_io_out ? io_r_94_b : _GEN_6613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6615 = 8'h5f == r_count_32_io_out ? io_r_95_b : _GEN_6614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6616 = 8'h60 == r_count_32_io_out ? io_r_96_b : _GEN_6615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6617 = 8'h61 == r_count_32_io_out ? io_r_97_b : _GEN_6616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6618 = 8'h62 == r_count_32_io_out ? io_r_98_b : _GEN_6617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6619 = 8'h63 == r_count_32_io_out ? io_r_99_b : _GEN_6618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6620 = 8'h64 == r_count_32_io_out ? io_r_100_b : _GEN_6619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6621 = 8'h65 == r_count_32_io_out ? io_r_101_b : _GEN_6620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6622 = 8'h66 == r_count_32_io_out ? io_r_102_b : _GEN_6621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6623 = 8'h67 == r_count_32_io_out ? io_r_103_b : _GEN_6622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6624 = 8'h68 == r_count_32_io_out ? io_r_104_b : _GEN_6623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6625 = 8'h69 == r_count_32_io_out ? io_r_105_b : _GEN_6624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6626 = 8'h6a == r_count_32_io_out ? io_r_106_b : _GEN_6625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6627 = 8'h6b == r_count_32_io_out ? io_r_107_b : _GEN_6626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6628 = 8'h6c == r_count_32_io_out ? io_r_108_b : _GEN_6627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6629 = 8'h6d == r_count_32_io_out ? io_r_109_b : _GEN_6628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6630 = 8'h6e == r_count_32_io_out ? io_r_110_b : _GEN_6629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6631 = 8'h6f == r_count_32_io_out ? io_r_111_b : _GEN_6630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6632 = 8'h70 == r_count_32_io_out ? io_r_112_b : _GEN_6631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6633 = 8'h71 == r_count_32_io_out ? io_r_113_b : _GEN_6632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6634 = 8'h72 == r_count_32_io_out ? io_r_114_b : _GEN_6633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6635 = 8'h73 == r_count_32_io_out ? io_r_115_b : _GEN_6634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6636 = 8'h74 == r_count_32_io_out ? io_r_116_b : _GEN_6635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6637 = 8'h75 == r_count_32_io_out ? io_r_117_b : _GEN_6636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6638 = 8'h76 == r_count_32_io_out ? io_r_118_b : _GEN_6637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6639 = 8'h77 == r_count_32_io_out ? io_r_119_b : _GEN_6638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6640 = 8'h78 == r_count_32_io_out ? io_r_120_b : _GEN_6639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6641 = 8'h79 == r_count_32_io_out ? io_r_121_b : _GEN_6640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6642 = 8'h7a == r_count_32_io_out ? io_r_122_b : _GEN_6641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6643 = 8'h7b == r_count_32_io_out ? io_r_123_b : _GEN_6642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6644 = 8'h7c == r_count_32_io_out ? io_r_124_b : _GEN_6643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6645 = 8'h7d == r_count_32_io_out ? io_r_125_b : _GEN_6644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6646 = 8'h7e == r_count_32_io_out ? io_r_126_b : _GEN_6645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6647 = 8'h7f == r_count_32_io_out ? io_r_127_b : _GEN_6646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6648 = 8'h80 == r_count_32_io_out ? io_r_128_b : _GEN_6647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6649 = 8'h81 == r_count_32_io_out ? io_r_129_b : _GEN_6648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6650 = 8'h82 == r_count_32_io_out ? io_r_130_b : _GEN_6649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6651 = 8'h83 == r_count_32_io_out ? io_r_131_b : _GEN_6650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6652 = 8'h84 == r_count_32_io_out ? io_r_132_b : _GEN_6651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6653 = 8'h85 == r_count_32_io_out ? io_r_133_b : _GEN_6652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6654 = 8'h86 == r_count_32_io_out ? io_r_134_b : _GEN_6653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6655 = 8'h87 == r_count_32_io_out ? io_r_135_b : _GEN_6654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6656 = 8'h88 == r_count_32_io_out ? io_r_136_b : _GEN_6655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6657 = 8'h89 == r_count_32_io_out ? io_r_137_b : _GEN_6656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6658 = 8'h8a == r_count_32_io_out ? io_r_138_b : _GEN_6657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6659 = 8'h8b == r_count_32_io_out ? io_r_139_b : _GEN_6658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6660 = 8'h8c == r_count_32_io_out ? io_r_140_b : _GEN_6659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6661 = 8'h8d == r_count_32_io_out ? io_r_141_b : _GEN_6660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6662 = 8'h8e == r_count_32_io_out ? io_r_142_b : _GEN_6661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6663 = 8'h8f == r_count_32_io_out ? io_r_143_b : _GEN_6662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6664 = 8'h90 == r_count_32_io_out ? io_r_144_b : _GEN_6663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6665 = 8'h91 == r_count_32_io_out ? io_r_145_b : _GEN_6664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6666 = 8'h92 == r_count_32_io_out ? io_r_146_b : _GEN_6665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6667 = 8'h93 == r_count_32_io_out ? io_r_147_b : _GEN_6666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6668 = 8'h94 == r_count_32_io_out ? io_r_148_b : _GEN_6667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6669 = 8'h95 == r_count_32_io_out ? io_r_149_b : _GEN_6668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6670 = 8'h96 == r_count_32_io_out ? io_r_150_b : _GEN_6669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6671 = 8'h97 == r_count_32_io_out ? io_r_151_b : _GEN_6670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6672 = 8'h98 == r_count_32_io_out ? io_r_152_b : _GEN_6671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6673 = 8'h99 == r_count_32_io_out ? io_r_153_b : _GEN_6672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6674 = 8'h9a == r_count_32_io_out ? io_r_154_b : _GEN_6673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6675 = 8'h9b == r_count_32_io_out ? io_r_155_b : _GEN_6674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6676 = 8'h9c == r_count_32_io_out ? io_r_156_b : _GEN_6675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6677 = 8'h9d == r_count_32_io_out ? io_r_157_b : _GEN_6676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6678 = 8'h9e == r_count_32_io_out ? io_r_158_b : _GEN_6677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6679 = 8'h9f == r_count_32_io_out ? io_r_159_b : _GEN_6678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6680 = 8'ha0 == r_count_32_io_out ? io_r_160_b : _GEN_6679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6681 = 8'ha1 == r_count_32_io_out ? io_r_161_b : _GEN_6680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6682 = 8'ha2 == r_count_32_io_out ? io_r_162_b : _GEN_6681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6683 = 8'ha3 == r_count_32_io_out ? io_r_163_b : _GEN_6682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6684 = 8'ha4 == r_count_32_io_out ? io_r_164_b : _GEN_6683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6685 = 8'ha5 == r_count_32_io_out ? io_r_165_b : _GEN_6684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6686 = 8'ha6 == r_count_32_io_out ? io_r_166_b : _GEN_6685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6687 = 8'ha7 == r_count_32_io_out ? io_r_167_b : _GEN_6686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6688 = 8'ha8 == r_count_32_io_out ? io_r_168_b : _GEN_6687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6689 = 8'ha9 == r_count_32_io_out ? io_r_169_b : _GEN_6688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6690 = 8'haa == r_count_32_io_out ? io_r_170_b : _GEN_6689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6691 = 8'hab == r_count_32_io_out ? io_r_171_b : _GEN_6690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6692 = 8'hac == r_count_32_io_out ? io_r_172_b : _GEN_6691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6693 = 8'had == r_count_32_io_out ? io_r_173_b : _GEN_6692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6694 = 8'hae == r_count_32_io_out ? io_r_174_b : _GEN_6693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6695 = 8'haf == r_count_32_io_out ? io_r_175_b : _GEN_6694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6696 = 8'hb0 == r_count_32_io_out ? io_r_176_b : _GEN_6695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6697 = 8'hb1 == r_count_32_io_out ? io_r_177_b : _GEN_6696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6698 = 8'hb2 == r_count_32_io_out ? io_r_178_b : _GEN_6697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6699 = 8'hb3 == r_count_32_io_out ? io_r_179_b : _GEN_6698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6700 = 8'hb4 == r_count_32_io_out ? io_r_180_b : _GEN_6699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6701 = 8'hb5 == r_count_32_io_out ? io_r_181_b : _GEN_6700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6702 = 8'hb6 == r_count_32_io_out ? io_r_182_b : _GEN_6701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6703 = 8'hb7 == r_count_32_io_out ? io_r_183_b : _GEN_6702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6704 = 8'hb8 == r_count_32_io_out ? io_r_184_b : _GEN_6703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6705 = 8'hb9 == r_count_32_io_out ? io_r_185_b : _GEN_6704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6706 = 8'hba == r_count_32_io_out ? io_r_186_b : _GEN_6705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6707 = 8'hbb == r_count_32_io_out ? io_r_187_b : _GEN_6706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6708 = 8'hbc == r_count_32_io_out ? io_r_188_b : _GEN_6707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6709 = 8'hbd == r_count_32_io_out ? io_r_189_b : _GEN_6708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6710 = 8'hbe == r_count_32_io_out ? io_r_190_b : _GEN_6709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6711 = 8'hbf == r_count_32_io_out ? io_r_191_b : _GEN_6710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6712 = 8'hc0 == r_count_32_io_out ? io_r_192_b : _GEN_6711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6713 = 8'hc1 == r_count_32_io_out ? io_r_193_b : _GEN_6712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6714 = 8'hc2 == r_count_32_io_out ? io_r_194_b : _GEN_6713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6715 = 8'hc3 == r_count_32_io_out ? io_r_195_b : _GEN_6714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6716 = 8'hc4 == r_count_32_io_out ? io_r_196_b : _GEN_6715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6717 = 8'hc5 == r_count_32_io_out ? io_r_197_b : _GEN_6716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6718 = 8'hc6 == r_count_32_io_out ? io_r_198_b : _GEN_6717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6721 = 8'h1 == r_count_33_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6722 = 8'h2 == r_count_33_io_out ? io_r_2_b : _GEN_6721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6723 = 8'h3 == r_count_33_io_out ? io_r_3_b : _GEN_6722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6724 = 8'h4 == r_count_33_io_out ? io_r_4_b : _GEN_6723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6725 = 8'h5 == r_count_33_io_out ? io_r_5_b : _GEN_6724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6726 = 8'h6 == r_count_33_io_out ? io_r_6_b : _GEN_6725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6727 = 8'h7 == r_count_33_io_out ? io_r_7_b : _GEN_6726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6728 = 8'h8 == r_count_33_io_out ? io_r_8_b : _GEN_6727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6729 = 8'h9 == r_count_33_io_out ? io_r_9_b : _GEN_6728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6730 = 8'ha == r_count_33_io_out ? io_r_10_b : _GEN_6729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6731 = 8'hb == r_count_33_io_out ? io_r_11_b : _GEN_6730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6732 = 8'hc == r_count_33_io_out ? io_r_12_b : _GEN_6731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6733 = 8'hd == r_count_33_io_out ? io_r_13_b : _GEN_6732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6734 = 8'he == r_count_33_io_out ? io_r_14_b : _GEN_6733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6735 = 8'hf == r_count_33_io_out ? io_r_15_b : _GEN_6734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6736 = 8'h10 == r_count_33_io_out ? io_r_16_b : _GEN_6735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6737 = 8'h11 == r_count_33_io_out ? io_r_17_b : _GEN_6736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6738 = 8'h12 == r_count_33_io_out ? io_r_18_b : _GEN_6737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6739 = 8'h13 == r_count_33_io_out ? io_r_19_b : _GEN_6738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6740 = 8'h14 == r_count_33_io_out ? io_r_20_b : _GEN_6739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6741 = 8'h15 == r_count_33_io_out ? io_r_21_b : _GEN_6740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6742 = 8'h16 == r_count_33_io_out ? io_r_22_b : _GEN_6741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6743 = 8'h17 == r_count_33_io_out ? io_r_23_b : _GEN_6742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6744 = 8'h18 == r_count_33_io_out ? io_r_24_b : _GEN_6743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6745 = 8'h19 == r_count_33_io_out ? io_r_25_b : _GEN_6744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6746 = 8'h1a == r_count_33_io_out ? io_r_26_b : _GEN_6745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6747 = 8'h1b == r_count_33_io_out ? io_r_27_b : _GEN_6746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6748 = 8'h1c == r_count_33_io_out ? io_r_28_b : _GEN_6747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6749 = 8'h1d == r_count_33_io_out ? io_r_29_b : _GEN_6748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6750 = 8'h1e == r_count_33_io_out ? io_r_30_b : _GEN_6749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6751 = 8'h1f == r_count_33_io_out ? io_r_31_b : _GEN_6750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6752 = 8'h20 == r_count_33_io_out ? io_r_32_b : _GEN_6751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6753 = 8'h21 == r_count_33_io_out ? io_r_33_b : _GEN_6752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6754 = 8'h22 == r_count_33_io_out ? io_r_34_b : _GEN_6753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6755 = 8'h23 == r_count_33_io_out ? io_r_35_b : _GEN_6754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6756 = 8'h24 == r_count_33_io_out ? io_r_36_b : _GEN_6755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6757 = 8'h25 == r_count_33_io_out ? io_r_37_b : _GEN_6756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6758 = 8'h26 == r_count_33_io_out ? io_r_38_b : _GEN_6757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6759 = 8'h27 == r_count_33_io_out ? io_r_39_b : _GEN_6758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6760 = 8'h28 == r_count_33_io_out ? io_r_40_b : _GEN_6759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6761 = 8'h29 == r_count_33_io_out ? io_r_41_b : _GEN_6760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6762 = 8'h2a == r_count_33_io_out ? io_r_42_b : _GEN_6761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6763 = 8'h2b == r_count_33_io_out ? io_r_43_b : _GEN_6762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6764 = 8'h2c == r_count_33_io_out ? io_r_44_b : _GEN_6763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6765 = 8'h2d == r_count_33_io_out ? io_r_45_b : _GEN_6764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6766 = 8'h2e == r_count_33_io_out ? io_r_46_b : _GEN_6765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6767 = 8'h2f == r_count_33_io_out ? io_r_47_b : _GEN_6766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6768 = 8'h30 == r_count_33_io_out ? io_r_48_b : _GEN_6767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6769 = 8'h31 == r_count_33_io_out ? io_r_49_b : _GEN_6768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6770 = 8'h32 == r_count_33_io_out ? io_r_50_b : _GEN_6769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6771 = 8'h33 == r_count_33_io_out ? io_r_51_b : _GEN_6770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6772 = 8'h34 == r_count_33_io_out ? io_r_52_b : _GEN_6771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6773 = 8'h35 == r_count_33_io_out ? io_r_53_b : _GEN_6772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6774 = 8'h36 == r_count_33_io_out ? io_r_54_b : _GEN_6773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6775 = 8'h37 == r_count_33_io_out ? io_r_55_b : _GEN_6774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6776 = 8'h38 == r_count_33_io_out ? io_r_56_b : _GEN_6775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6777 = 8'h39 == r_count_33_io_out ? io_r_57_b : _GEN_6776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6778 = 8'h3a == r_count_33_io_out ? io_r_58_b : _GEN_6777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6779 = 8'h3b == r_count_33_io_out ? io_r_59_b : _GEN_6778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6780 = 8'h3c == r_count_33_io_out ? io_r_60_b : _GEN_6779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6781 = 8'h3d == r_count_33_io_out ? io_r_61_b : _GEN_6780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6782 = 8'h3e == r_count_33_io_out ? io_r_62_b : _GEN_6781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6783 = 8'h3f == r_count_33_io_out ? io_r_63_b : _GEN_6782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6784 = 8'h40 == r_count_33_io_out ? io_r_64_b : _GEN_6783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6785 = 8'h41 == r_count_33_io_out ? io_r_65_b : _GEN_6784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6786 = 8'h42 == r_count_33_io_out ? io_r_66_b : _GEN_6785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6787 = 8'h43 == r_count_33_io_out ? io_r_67_b : _GEN_6786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6788 = 8'h44 == r_count_33_io_out ? io_r_68_b : _GEN_6787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6789 = 8'h45 == r_count_33_io_out ? io_r_69_b : _GEN_6788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6790 = 8'h46 == r_count_33_io_out ? io_r_70_b : _GEN_6789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6791 = 8'h47 == r_count_33_io_out ? io_r_71_b : _GEN_6790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6792 = 8'h48 == r_count_33_io_out ? io_r_72_b : _GEN_6791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6793 = 8'h49 == r_count_33_io_out ? io_r_73_b : _GEN_6792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6794 = 8'h4a == r_count_33_io_out ? io_r_74_b : _GEN_6793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6795 = 8'h4b == r_count_33_io_out ? io_r_75_b : _GEN_6794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6796 = 8'h4c == r_count_33_io_out ? io_r_76_b : _GEN_6795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6797 = 8'h4d == r_count_33_io_out ? io_r_77_b : _GEN_6796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6798 = 8'h4e == r_count_33_io_out ? io_r_78_b : _GEN_6797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6799 = 8'h4f == r_count_33_io_out ? io_r_79_b : _GEN_6798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6800 = 8'h50 == r_count_33_io_out ? io_r_80_b : _GEN_6799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6801 = 8'h51 == r_count_33_io_out ? io_r_81_b : _GEN_6800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6802 = 8'h52 == r_count_33_io_out ? io_r_82_b : _GEN_6801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6803 = 8'h53 == r_count_33_io_out ? io_r_83_b : _GEN_6802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6804 = 8'h54 == r_count_33_io_out ? io_r_84_b : _GEN_6803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6805 = 8'h55 == r_count_33_io_out ? io_r_85_b : _GEN_6804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6806 = 8'h56 == r_count_33_io_out ? io_r_86_b : _GEN_6805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6807 = 8'h57 == r_count_33_io_out ? io_r_87_b : _GEN_6806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6808 = 8'h58 == r_count_33_io_out ? io_r_88_b : _GEN_6807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6809 = 8'h59 == r_count_33_io_out ? io_r_89_b : _GEN_6808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6810 = 8'h5a == r_count_33_io_out ? io_r_90_b : _GEN_6809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6811 = 8'h5b == r_count_33_io_out ? io_r_91_b : _GEN_6810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6812 = 8'h5c == r_count_33_io_out ? io_r_92_b : _GEN_6811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6813 = 8'h5d == r_count_33_io_out ? io_r_93_b : _GEN_6812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6814 = 8'h5e == r_count_33_io_out ? io_r_94_b : _GEN_6813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6815 = 8'h5f == r_count_33_io_out ? io_r_95_b : _GEN_6814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6816 = 8'h60 == r_count_33_io_out ? io_r_96_b : _GEN_6815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6817 = 8'h61 == r_count_33_io_out ? io_r_97_b : _GEN_6816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6818 = 8'h62 == r_count_33_io_out ? io_r_98_b : _GEN_6817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6819 = 8'h63 == r_count_33_io_out ? io_r_99_b : _GEN_6818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6820 = 8'h64 == r_count_33_io_out ? io_r_100_b : _GEN_6819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6821 = 8'h65 == r_count_33_io_out ? io_r_101_b : _GEN_6820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6822 = 8'h66 == r_count_33_io_out ? io_r_102_b : _GEN_6821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6823 = 8'h67 == r_count_33_io_out ? io_r_103_b : _GEN_6822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6824 = 8'h68 == r_count_33_io_out ? io_r_104_b : _GEN_6823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6825 = 8'h69 == r_count_33_io_out ? io_r_105_b : _GEN_6824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6826 = 8'h6a == r_count_33_io_out ? io_r_106_b : _GEN_6825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6827 = 8'h6b == r_count_33_io_out ? io_r_107_b : _GEN_6826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6828 = 8'h6c == r_count_33_io_out ? io_r_108_b : _GEN_6827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6829 = 8'h6d == r_count_33_io_out ? io_r_109_b : _GEN_6828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6830 = 8'h6e == r_count_33_io_out ? io_r_110_b : _GEN_6829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6831 = 8'h6f == r_count_33_io_out ? io_r_111_b : _GEN_6830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6832 = 8'h70 == r_count_33_io_out ? io_r_112_b : _GEN_6831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6833 = 8'h71 == r_count_33_io_out ? io_r_113_b : _GEN_6832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6834 = 8'h72 == r_count_33_io_out ? io_r_114_b : _GEN_6833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6835 = 8'h73 == r_count_33_io_out ? io_r_115_b : _GEN_6834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6836 = 8'h74 == r_count_33_io_out ? io_r_116_b : _GEN_6835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6837 = 8'h75 == r_count_33_io_out ? io_r_117_b : _GEN_6836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6838 = 8'h76 == r_count_33_io_out ? io_r_118_b : _GEN_6837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6839 = 8'h77 == r_count_33_io_out ? io_r_119_b : _GEN_6838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6840 = 8'h78 == r_count_33_io_out ? io_r_120_b : _GEN_6839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6841 = 8'h79 == r_count_33_io_out ? io_r_121_b : _GEN_6840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6842 = 8'h7a == r_count_33_io_out ? io_r_122_b : _GEN_6841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6843 = 8'h7b == r_count_33_io_out ? io_r_123_b : _GEN_6842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6844 = 8'h7c == r_count_33_io_out ? io_r_124_b : _GEN_6843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6845 = 8'h7d == r_count_33_io_out ? io_r_125_b : _GEN_6844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6846 = 8'h7e == r_count_33_io_out ? io_r_126_b : _GEN_6845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6847 = 8'h7f == r_count_33_io_out ? io_r_127_b : _GEN_6846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6848 = 8'h80 == r_count_33_io_out ? io_r_128_b : _GEN_6847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6849 = 8'h81 == r_count_33_io_out ? io_r_129_b : _GEN_6848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6850 = 8'h82 == r_count_33_io_out ? io_r_130_b : _GEN_6849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6851 = 8'h83 == r_count_33_io_out ? io_r_131_b : _GEN_6850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6852 = 8'h84 == r_count_33_io_out ? io_r_132_b : _GEN_6851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6853 = 8'h85 == r_count_33_io_out ? io_r_133_b : _GEN_6852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6854 = 8'h86 == r_count_33_io_out ? io_r_134_b : _GEN_6853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6855 = 8'h87 == r_count_33_io_out ? io_r_135_b : _GEN_6854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6856 = 8'h88 == r_count_33_io_out ? io_r_136_b : _GEN_6855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6857 = 8'h89 == r_count_33_io_out ? io_r_137_b : _GEN_6856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6858 = 8'h8a == r_count_33_io_out ? io_r_138_b : _GEN_6857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6859 = 8'h8b == r_count_33_io_out ? io_r_139_b : _GEN_6858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6860 = 8'h8c == r_count_33_io_out ? io_r_140_b : _GEN_6859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6861 = 8'h8d == r_count_33_io_out ? io_r_141_b : _GEN_6860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6862 = 8'h8e == r_count_33_io_out ? io_r_142_b : _GEN_6861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6863 = 8'h8f == r_count_33_io_out ? io_r_143_b : _GEN_6862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6864 = 8'h90 == r_count_33_io_out ? io_r_144_b : _GEN_6863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6865 = 8'h91 == r_count_33_io_out ? io_r_145_b : _GEN_6864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6866 = 8'h92 == r_count_33_io_out ? io_r_146_b : _GEN_6865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6867 = 8'h93 == r_count_33_io_out ? io_r_147_b : _GEN_6866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6868 = 8'h94 == r_count_33_io_out ? io_r_148_b : _GEN_6867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6869 = 8'h95 == r_count_33_io_out ? io_r_149_b : _GEN_6868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6870 = 8'h96 == r_count_33_io_out ? io_r_150_b : _GEN_6869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6871 = 8'h97 == r_count_33_io_out ? io_r_151_b : _GEN_6870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6872 = 8'h98 == r_count_33_io_out ? io_r_152_b : _GEN_6871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6873 = 8'h99 == r_count_33_io_out ? io_r_153_b : _GEN_6872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6874 = 8'h9a == r_count_33_io_out ? io_r_154_b : _GEN_6873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6875 = 8'h9b == r_count_33_io_out ? io_r_155_b : _GEN_6874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6876 = 8'h9c == r_count_33_io_out ? io_r_156_b : _GEN_6875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6877 = 8'h9d == r_count_33_io_out ? io_r_157_b : _GEN_6876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6878 = 8'h9e == r_count_33_io_out ? io_r_158_b : _GEN_6877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6879 = 8'h9f == r_count_33_io_out ? io_r_159_b : _GEN_6878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6880 = 8'ha0 == r_count_33_io_out ? io_r_160_b : _GEN_6879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6881 = 8'ha1 == r_count_33_io_out ? io_r_161_b : _GEN_6880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6882 = 8'ha2 == r_count_33_io_out ? io_r_162_b : _GEN_6881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6883 = 8'ha3 == r_count_33_io_out ? io_r_163_b : _GEN_6882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6884 = 8'ha4 == r_count_33_io_out ? io_r_164_b : _GEN_6883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6885 = 8'ha5 == r_count_33_io_out ? io_r_165_b : _GEN_6884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6886 = 8'ha6 == r_count_33_io_out ? io_r_166_b : _GEN_6885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6887 = 8'ha7 == r_count_33_io_out ? io_r_167_b : _GEN_6886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6888 = 8'ha8 == r_count_33_io_out ? io_r_168_b : _GEN_6887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6889 = 8'ha9 == r_count_33_io_out ? io_r_169_b : _GEN_6888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6890 = 8'haa == r_count_33_io_out ? io_r_170_b : _GEN_6889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6891 = 8'hab == r_count_33_io_out ? io_r_171_b : _GEN_6890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6892 = 8'hac == r_count_33_io_out ? io_r_172_b : _GEN_6891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6893 = 8'had == r_count_33_io_out ? io_r_173_b : _GEN_6892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6894 = 8'hae == r_count_33_io_out ? io_r_174_b : _GEN_6893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6895 = 8'haf == r_count_33_io_out ? io_r_175_b : _GEN_6894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6896 = 8'hb0 == r_count_33_io_out ? io_r_176_b : _GEN_6895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6897 = 8'hb1 == r_count_33_io_out ? io_r_177_b : _GEN_6896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6898 = 8'hb2 == r_count_33_io_out ? io_r_178_b : _GEN_6897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6899 = 8'hb3 == r_count_33_io_out ? io_r_179_b : _GEN_6898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6900 = 8'hb4 == r_count_33_io_out ? io_r_180_b : _GEN_6899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6901 = 8'hb5 == r_count_33_io_out ? io_r_181_b : _GEN_6900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6902 = 8'hb6 == r_count_33_io_out ? io_r_182_b : _GEN_6901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6903 = 8'hb7 == r_count_33_io_out ? io_r_183_b : _GEN_6902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6904 = 8'hb8 == r_count_33_io_out ? io_r_184_b : _GEN_6903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6905 = 8'hb9 == r_count_33_io_out ? io_r_185_b : _GEN_6904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6906 = 8'hba == r_count_33_io_out ? io_r_186_b : _GEN_6905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6907 = 8'hbb == r_count_33_io_out ? io_r_187_b : _GEN_6906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6908 = 8'hbc == r_count_33_io_out ? io_r_188_b : _GEN_6907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6909 = 8'hbd == r_count_33_io_out ? io_r_189_b : _GEN_6908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6910 = 8'hbe == r_count_33_io_out ? io_r_190_b : _GEN_6909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6911 = 8'hbf == r_count_33_io_out ? io_r_191_b : _GEN_6910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6912 = 8'hc0 == r_count_33_io_out ? io_r_192_b : _GEN_6911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6913 = 8'hc1 == r_count_33_io_out ? io_r_193_b : _GEN_6912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6914 = 8'hc2 == r_count_33_io_out ? io_r_194_b : _GEN_6913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6915 = 8'hc3 == r_count_33_io_out ? io_r_195_b : _GEN_6914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6916 = 8'hc4 == r_count_33_io_out ? io_r_196_b : _GEN_6915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6917 = 8'hc5 == r_count_33_io_out ? io_r_197_b : _GEN_6916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6918 = 8'hc6 == r_count_33_io_out ? io_r_198_b : _GEN_6917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6921 = 8'h1 == r_count_34_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6922 = 8'h2 == r_count_34_io_out ? io_r_2_b : _GEN_6921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6923 = 8'h3 == r_count_34_io_out ? io_r_3_b : _GEN_6922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6924 = 8'h4 == r_count_34_io_out ? io_r_4_b : _GEN_6923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6925 = 8'h5 == r_count_34_io_out ? io_r_5_b : _GEN_6924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6926 = 8'h6 == r_count_34_io_out ? io_r_6_b : _GEN_6925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6927 = 8'h7 == r_count_34_io_out ? io_r_7_b : _GEN_6926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6928 = 8'h8 == r_count_34_io_out ? io_r_8_b : _GEN_6927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6929 = 8'h9 == r_count_34_io_out ? io_r_9_b : _GEN_6928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6930 = 8'ha == r_count_34_io_out ? io_r_10_b : _GEN_6929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6931 = 8'hb == r_count_34_io_out ? io_r_11_b : _GEN_6930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6932 = 8'hc == r_count_34_io_out ? io_r_12_b : _GEN_6931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6933 = 8'hd == r_count_34_io_out ? io_r_13_b : _GEN_6932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6934 = 8'he == r_count_34_io_out ? io_r_14_b : _GEN_6933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6935 = 8'hf == r_count_34_io_out ? io_r_15_b : _GEN_6934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6936 = 8'h10 == r_count_34_io_out ? io_r_16_b : _GEN_6935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6937 = 8'h11 == r_count_34_io_out ? io_r_17_b : _GEN_6936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6938 = 8'h12 == r_count_34_io_out ? io_r_18_b : _GEN_6937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6939 = 8'h13 == r_count_34_io_out ? io_r_19_b : _GEN_6938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6940 = 8'h14 == r_count_34_io_out ? io_r_20_b : _GEN_6939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6941 = 8'h15 == r_count_34_io_out ? io_r_21_b : _GEN_6940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6942 = 8'h16 == r_count_34_io_out ? io_r_22_b : _GEN_6941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6943 = 8'h17 == r_count_34_io_out ? io_r_23_b : _GEN_6942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6944 = 8'h18 == r_count_34_io_out ? io_r_24_b : _GEN_6943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6945 = 8'h19 == r_count_34_io_out ? io_r_25_b : _GEN_6944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6946 = 8'h1a == r_count_34_io_out ? io_r_26_b : _GEN_6945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6947 = 8'h1b == r_count_34_io_out ? io_r_27_b : _GEN_6946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6948 = 8'h1c == r_count_34_io_out ? io_r_28_b : _GEN_6947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6949 = 8'h1d == r_count_34_io_out ? io_r_29_b : _GEN_6948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6950 = 8'h1e == r_count_34_io_out ? io_r_30_b : _GEN_6949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6951 = 8'h1f == r_count_34_io_out ? io_r_31_b : _GEN_6950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6952 = 8'h20 == r_count_34_io_out ? io_r_32_b : _GEN_6951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6953 = 8'h21 == r_count_34_io_out ? io_r_33_b : _GEN_6952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6954 = 8'h22 == r_count_34_io_out ? io_r_34_b : _GEN_6953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6955 = 8'h23 == r_count_34_io_out ? io_r_35_b : _GEN_6954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6956 = 8'h24 == r_count_34_io_out ? io_r_36_b : _GEN_6955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6957 = 8'h25 == r_count_34_io_out ? io_r_37_b : _GEN_6956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6958 = 8'h26 == r_count_34_io_out ? io_r_38_b : _GEN_6957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6959 = 8'h27 == r_count_34_io_out ? io_r_39_b : _GEN_6958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6960 = 8'h28 == r_count_34_io_out ? io_r_40_b : _GEN_6959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6961 = 8'h29 == r_count_34_io_out ? io_r_41_b : _GEN_6960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6962 = 8'h2a == r_count_34_io_out ? io_r_42_b : _GEN_6961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6963 = 8'h2b == r_count_34_io_out ? io_r_43_b : _GEN_6962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6964 = 8'h2c == r_count_34_io_out ? io_r_44_b : _GEN_6963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6965 = 8'h2d == r_count_34_io_out ? io_r_45_b : _GEN_6964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6966 = 8'h2e == r_count_34_io_out ? io_r_46_b : _GEN_6965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6967 = 8'h2f == r_count_34_io_out ? io_r_47_b : _GEN_6966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6968 = 8'h30 == r_count_34_io_out ? io_r_48_b : _GEN_6967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6969 = 8'h31 == r_count_34_io_out ? io_r_49_b : _GEN_6968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6970 = 8'h32 == r_count_34_io_out ? io_r_50_b : _GEN_6969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6971 = 8'h33 == r_count_34_io_out ? io_r_51_b : _GEN_6970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6972 = 8'h34 == r_count_34_io_out ? io_r_52_b : _GEN_6971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6973 = 8'h35 == r_count_34_io_out ? io_r_53_b : _GEN_6972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6974 = 8'h36 == r_count_34_io_out ? io_r_54_b : _GEN_6973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6975 = 8'h37 == r_count_34_io_out ? io_r_55_b : _GEN_6974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6976 = 8'h38 == r_count_34_io_out ? io_r_56_b : _GEN_6975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6977 = 8'h39 == r_count_34_io_out ? io_r_57_b : _GEN_6976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6978 = 8'h3a == r_count_34_io_out ? io_r_58_b : _GEN_6977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6979 = 8'h3b == r_count_34_io_out ? io_r_59_b : _GEN_6978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6980 = 8'h3c == r_count_34_io_out ? io_r_60_b : _GEN_6979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6981 = 8'h3d == r_count_34_io_out ? io_r_61_b : _GEN_6980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6982 = 8'h3e == r_count_34_io_out ? io_r_62_b : _GEN_6981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6983 = 8'h3f == r_count_34_io_out ? io_r_63_b : _GEN_6982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6984 = 8'h40 == r_count_34_io_out ? io_r_64_b : _GEN_6983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6985 = 8'h41 == r_count_34_io_out ? io_r_65_b : _GEN_6984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6986 = 8'h42 == r_count_34_io_out ? io_r_66_b : _GEN_6985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6987 = 8'h43 == r_count_34_io_out ? io_r_67_b : _GEN_6986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6988 = 8'h44 == r_count_34_io_out ? io_r_68_b : _GEN_6987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6989 = 8'h45 == r_count_34_io_out ? io_r_69_b : _GEN_6988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6990 = 8'h46 == r_count_34_io_out ? io_r_70_b : _GEN_6989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6991 = 8'h47 == r_count_34_io_out ? io_r_71_b : _GEN_6990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6992 = 8'h48 == r_count_34_io_out ? io_r_72_b : _GEN_6991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6993 = 8'h49 == r_count_34_io_out ? io_r_73_b : _GEN_6992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6994 = 8'h4a == r_count_34_io_out ? io_r_74_b : _GEN_6993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6995 = 8'h4b == r_count_34_io_out ? io_r_75_b : _GEN_6994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6996 = 8'h4c == r_count_34_io_out ? io_r_76_b : _GEN_6995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6997 = 8'h4d == r_count_34_io_out ? io_r_77_b : _GEN_6996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6998 = 8'h4e == r_count_34_io_out ? io_r_78_b : _GEN_6997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_6999 = 8'h4f == r_count_34_io_out ? io_r_79_b : _GEN_6998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7000 = 8'h50 == r_count_34_io_out ? io_r_80_b : _GEN_6999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7001 = 8'h51 == r_count_34_io_out ? io_r_81_b : _GEN_7000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7002 = 8'h52 == r_count_34_io_out ? io_r_82_b : _GEN_7001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7003 = 8'h53 == r_count_34_io_out ? io_r_83_b : _GEN_7002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7004 = 8'h54 == r_count_34_io_out ? io_r_84_b : _GEN_7003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7005 = 8'h55 == r_count_34_io_out ? io_r_85_b : _GEN_7004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7006 = 8'h56 == r_count_34_io_out ? io_r_86_b : _GEN_7005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7007 = 8'h57 == r_count_34_io_out ? io_r_87_b : _GEN_7006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7008 = 8'h58 == r_count_34_io_out ? io_r_88_b : _GEN_7007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7009 = 8'h59 == r_count_34_io_out ? io_r_89_b : _GEN_7008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7010 = 8'h5a == r_count_34_io_out ? io_r_90_b : _GEN_7009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7011 = 8'h5b == r_count_34_io_out ? io_r_91_b : _GEN_7010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7012 = 8'h5c == r_count_34_io_out ? io_r_92_b : _GEN_7011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7013 = 8'h5d == r_count_34_io_out ? io_r_93_b : _GEN_7012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7014 = 8'h5e == r_count_34_io_out ? io_r_94_b : _GEN_7013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7015 = 8'h5f == r_count_34_io_out ? io_r_95_b : _GEN_7014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7016 = 8'h60 == r_count_34_io_out ? io_r_96_b : _GEN_7015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7017 = 8'h61 == r_count_34_io_out ? io_r_97_b : _GEN_7016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7018 = 8'h62 == r_count_34_io_out ? io_r_98_b : _GEN_7017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7019 = 8'h63 == r_count_34_io_out ? io_r_99_b : _GEN_7018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7020 = 8'h64 == r_count_34_io_out ? io_r_100_b : _GEN_7019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7021 = 8'h65 == r_count_34_io_out ? io_r_101_b : _GEN_7020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7022 = 8'h66 == r_count_34_io_out ? io_r_102_b : _GEN_7021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7023 = 8'h67 == r_count_34_io_out ? io_r_103_b : _GEN_7022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7024 = 8'h68 == r_count_34_io_out ? io_r_104_b : _GEN_7023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7025 = 8'h69 == r_count_34_io_out ? io_r_105_b : _GEN_7024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7026 = 8'h6a == r_count_34_io_out ? io_r_106_b : _GEN_7025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7027 = 8'h6b == r_count_34_io_out ? io_r_107_b : _GEN_7026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7028 = 8'h6c == r_count_34_io_out ? io_r_108_b : _GEN_7027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7029 = 8'h6d == r_count_34_io_out ? io_r_109_b : _GEN_7028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7030 = 8'h6e == r_count_34_io_out ? io_r_110_b : _GEN_7029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7031 = 8'h6f == r_count_34_io_out ? io_r_111_b : _GEN_7030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7032 = 8'h70 == r_count_34_io_out ? io_r_112_b : _GEN_7031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7033 = 8'h71 == r_count_34_io_out ? io_r_113_b : _GEN_7032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7034 = 8'h72 == r_count_34_io_out ? io_r_114_b : _GEN_7033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7035 = 8'h73 == r_count_34_io_out ? io_r_115_b : _GEN_7034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7036 = 8'h74 == r_count_34_io_out ? io_r_116_b : _GEN_7035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7037 = 8'h75 == r_count_34_io_out ? io_r_117_b : _GEN_7036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7038 = 8'h76 == r_count_34_io_out ? io_r_118_b : _GEN_7037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7039 = 8'h77 == r_count_34_io_out ? io_r_119_b : _GEN_7038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7040 = 8'h78 == r_count_34_io_out ? io_r_120_b : _GEN_7039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7041 = 8'h79 == r_count_34_io_out ? io_r_121_b : _GEN_7040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7042 = 8'h7a == r_count_34_io_out ? io_r_122_b : _GEN_7041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7043 = 8'h7b == r_count_34_io_out ? io_r_123_b : _GEN_7042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7044 = 8'h7c == r_count_34_io_out ? io_r_124_b : _GEN_7043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7045 = 8'h7d == r_count_34_io_out ? io_r_125_b : _GEN_7044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7046 = 8'h7e == r_count_34_io_out ? io_r_126_b : _GEN_7045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7047 = 8'h7f == r_count_34_io_out ? io_r_127_b : _GEN_7046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7048 = 8'h80 == r_count_34_io_out ? io_r_128_b : _GEN_7047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7049 = 8'h81 == r_count_34_io_out ? io_r_129_b : _GEN_7048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7050 = 8'h82 == r_count_34_io_out ? io_r_130_b : _GEN_7049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7051 = 8'h83 == r_count_34_io_out ? io_r_131_b : _GEN_7050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7052 = 8'h84 == r_count_34_io_out ? io_r_132_b : _GEN_7051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7053 = 8'h85 == r_count_34_io_out ? io_r_133_b : _GEN_7052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7054 = 8'h86 == r_count_34_io_out ? io_r_134_b : _GEN_7053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7055 = 8'h87 == r_count_34_io_out ? io_r_135_b : _GEN_7054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7056 = 8'h88 == r_count_34_io_out ? io_r_136_b : _GEN_7055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7057 = 8'h89 == r_count_34_io_out ? io_r_137_b : _GEN_7056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7058 = 8'h8a == r_count_34_io_out ? io_r_138_b : _GEN_7057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7059 = 8'h8b == r_count_34_io_out ? io_r_139_b : _GEN_7058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7060 = 8'h8c == r_count_34_io_out ? io_r_140_b : _GEN_7059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7061 = 8'h8d == r_count_34_io_out ? io_r_141_b : _GEN_7060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7062 = 8'h8e == r_count_34_io_out ? io_r_142_b : _GEN_7061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7063 = 8'h8f == r_count_34_io_out ? io_r_143_b : _GEN_7062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7064 = 8'h90 == r_count_34_io_out ? io_r_144_b : _GEN_7063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7065 = 8'h91 == r_count_34_io_out ? io_r_145_b : _GEN_7064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7066 = 8'h92 == r_count_34_io_out ? io_r_146_b : _GEN_7065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7067 = 8'h93 == r_count_34_io_out ? io_r_147_b : _GEN_7066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7068 = 8'h94 == r_count_34_io_out ? io_r_148_b : _GEN_7067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7069 = 8'h95 == r_count_34_io_out ? io_r_149_b : _GEN_7068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7070 = 8'h96 == r_count_34_io_out ? io_r_150_b : _GEN_7069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7071 = 8'h97 == r_count_34_io_out ? io_r_151_b : _GEN_7070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7072 = 8'h98 == r_count_34_io_out ? io_r_152_b : _GEN_7071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7073 = 8'h99 == r_count_34_io_out ? io_r_153_b : _GEN_7072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7074 = 8'h9a == r_count_34_io_out ? io_r_154_b : _GEN_7073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7075 = 8'h9b == r_count_34_io_out ? io_r_155_b : _GEN_7074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7076 = 8'h9c == r_count_34_io_out ? io_r_156_b : _GEN_7075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7077 = 8'h9d == r_count_34_io_out ? io_r_157_b : _GEN_7076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7078 = 8'h9e == r_count_34_io_out ? io_r_158_b : _GEN_7077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7079 = 8'h9f == r_count_34_io_out ? io_r_159_b : _GEN_7078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7080 = 8'ha0 == r_count_34_io_out ? io_r_160_b : _GEN_7079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7081 = 8'ha1 == r_count_34_io_out ? io_r_161_b : _GEN_7080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7082 = 8'ha2 == r_count_34_io_out ? io_r_162_b : _GEN_7081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7083 = 8'ha3 == r_count_34_io_out ? io_r_163_b : _GEN_7082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7084 = 8'ha4 == r_count_34_io_out ? io_r_164_b : _GEN_7083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7085 = 8'ha5 == r_count_34_io_out ? io_r_165_b : _GEN_7084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7086 = 8'ha6 == r_count_34_io_out ? io_r_166_b : _GEN_7085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7087 = 8'ha7 == r_count_34_io_out ? io_r_167_b : _GEN_7086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7088 = 8'ha8 == r_count_34_io_out ? io_r_168_b : _GEN_7087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7089 = 8'ha9 == r_count_34_io_out ? io_r_169_b : _GEN_7088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7090 = 8'haa == r_count_34_io_out ? io_r_170_b : _GEN_7089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7091 = 8'hab == r_count_34_io_out ? io_r_171_b : _GEN_7090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7092 = 8'hac == r_count_34_io_out ? io_r_172_b : _GEN_7091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7093 = 8'had == r_count_34_io_out ? io_r_173_b : _GEN_7092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7094 = 8'hae == r_count_34_io_out ? io_r_174_b : _GEN_7093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7095 = 8'haf == r_count_34_io_out ? io_r_175_b : _GEN_7094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7096 = 8'hb0 == r_count_34_io_out ? io_r_176_b : _GEN_7095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7097 = 8'hb1 == r_count_34_io_out ? io_r_177_b : _GEN_7096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7098 = 8'hb2 == r_count_34_io_out ? io_r_178_b : _GEN_7097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7099 = 8'hb3 == r_count_34_io_out ? io_r_179_b : _GEN_7098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7100 = 8'hb4 == r_count_34_io_out ? io_r_180_b : _GEN_7099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7101 = 8'hb5 == r_count_34_io_out ? io_r_181_b : _GEN_7100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7102 = 8'hb6 == r_count_34_io_out ? io_r_182_b : _GEN_7101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7103 = 8'hb7 == r_count_34_io_out ? io_r_183_b : _GEN_7102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7104 = 8'hb8 == r_count_34_io_out ? io_r_184_b : _GEN_7103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7105 = 8'hb9 == r_count_34_io_out ? io_r_185_b : _GEN_7104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7106 = 8'hba == r_count_34_io_out ? io_r_186_b : _GEN_7105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7107 = 8'hbb == r_count_34_io_out ? io_r_187_b : _GEN_7106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7108 = 8'hbc == r_count_34_io_out ? io_r_188_b : _GEN_7107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7109 = 8'hbd == r_count_34_io_out ? io_r_189_b : _GEN_7108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7110 = 8'hbe == r_count_34_io_out ? io_r_190_b : _GEN_7109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7111 = 8'hbf == r_count_34_io_out ? io_r_191_b : _GEN_7110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7112 = 8'hc0 == r_count_34_io_out ? io_r_192_b : _GEN_7111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7113 = 8'hc1 == r_count_34_io_out ? io_r_193_b : _GEN_7112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7114 = 8'hc2 == r_count_34_io_out ? io_r_194_b : _GEN_7113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7115 = 8'hc3 == r_count_34_io_out ? io_r_195_b : _GEN_7114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7116 = 8'hc4 == r_count_34_io_out ? io_r_196_b : _GEN_7115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7117 = 8'hc5 == r_count_34_io_out ? io_r_197_b : _GEN_7116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7118 = 8'hc6 == r_count_34_io_out ? io_r_198_b : _GEN_7117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7121 = 8'h1 == r_count_35_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7122 = 8'h2 == r_count_35_io_out ? io_r_2_b : _GEN_7121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7123 = 8'h3 == r_count_35_io_out ? io_r_3_b : _GEN_7122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7124 = 8'h4 == r_count_35_io_out ? io_r_4_b : _GEN_7123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7125 = 8'h5 == r_count_35_io_out ? io_r_5_b : _GEN_7124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7126 = 8'h6 == r_count_35_io_out ? io_r_6_b : _GEN_7125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7127 = 8'h7 == r_count_35_io_out ? io_r_7_b : _GEN_7126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7128 = 8'h8 == r_count_35_io_out ? io_r_8_b : _GEN_7127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7129 = 8'h9 == r_count_35_io_out ? io_r_9_b : _GEN_7128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7130 = 8'ha == r_count_35_io_out ? io_r_10_b : _GEN_7129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7131 = 8'hb == r_count_35_io_out ? io_r_11_b : _GEN_7130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7132 = 8'hc == r_count_35_io_out ? io_r_12_b : _GEN_7131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7133 = 8'hd == r_count_35_io_out ? io_r_13_b : _GEN_7132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7134 = 8'he == r_count_35_io_out ? io_r_14_b : _GEN_7133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7135 = 8'hf == r_count_35_io_out ? io_r_15_b : _GEN_7134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7136 = 8'h10 == r_count_35_io_out ? io_r_16_b : _GEN_7135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7137 = 8'h11 == r_count_35_io_out ? io_r_17_b : _GEN_7136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7138 = 8'h12 == r_count_35_io_out ? io_r_18_b : _GEN_7137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7139 = 8'h13 == r_count_35_io_out ? io_r_19_b : _GEN_7138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7140 = 8'h14 == r_count_35_io_out ? io_r_20_b : _GEN_7139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7141 = 8'h15 == r_count_35_io_out ? io_r_21_b : _GEN_7140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7142 = 8'h16 == r_count_35_io_out ? io_r_22_b : _GEN_7141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7143 = 8'h17 == r_count_35_io_out ? io_r_23_b : _GEN_7142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7144 = 8'h18 == r_count_35_io_out ? io_r_24_b : _GEN_7143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7145 = 8'h19 == r_count_35_io_out ? io_r_25_b : _GEN_7144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7146 = 8'h1a == r_count_35_io_out ? io_r_26_b : _GEN_7145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7147 = 8'h1b == r_count_35_io_out ? io_r_27_b : _GEN_7146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7148 = 8'h1c == r_count_35_io_out ? io_r_28_b : _GEN_7147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7149 = 8'h1d == r_count_35_io_out ? io_r_29_b : _GEN_7148; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7150 = 8'h1e == r_count_35_io_out ? io_r_30_b : _GEN_7149; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7151 = 8'h1f == r_count_35_io_out ? io_r_31_b : _GEN_7150; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7152 = 8'h20 == r_count_35_io_out ? io_r_32_b : _GEN_7151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7153 = 8'h21 == r_count_35_io_out ? io_r_33_b : _GEN_7152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7154 = 8'h22 == r_count_35_io_out ? io_r_34_b : _GEN_7153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7155 = 8'h23 == r_count_35_io_out ? io_r_35_b : _GEN_7154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7156 = 8'h24 == r_count_35_io_out ? io_r_36_b : _GEN_7155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7157 = 8'h25 == r_count_35_io_out ? io_r_37_b : _GEN_7156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7158 = 8'h26 == r_count_35_io_out ? io_r_38_b : _GEN_7157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7159 = 8'h27 == r_count_35_io_out ? io_r_39_b : _GEN_7158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7160 = 8'h28 == r_count_35_io_out ? io_r_40_b : _GEN_7159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7161 = 8'h29 == r_count_35_io_out ? io_r_41_b : _GEN_7160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7162 = 8'h2a == r_count_35_io_out ? io_r_42_b : _GEN_7161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7163 = 8'h2b == r_count_35_io_out ? io_r_43_b : _GEN_7162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7164 = 8'h2c == r_count_35_io_out ? io_r_44_b : _GEN_7163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7165 = 8'h2d == r_count_35_io_out ? io_r_45_b : _GEN_7164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7166 = 8'h2e == r_count_35_io_out ? io_r_46_b : _GEN_7165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7167 = 8'h2f == r_count_35_io_out ? io_r_47_b : _GEN_7166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7168 = 8'h30 == r_count_35_io_out ? io_r_48_b : _GEN_7167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7169 = 8'h31 == r_count_35_io_out ? io_r_49_b : _GEN_7168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7170 = 8'h32 == r_count_35_io_out ? io_r_50_b : _GEN_7169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7171 = 8'h33 == r_count_35_io_out ? io_r_51_b : _GEN_7170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7172 = 8'h34 == r_count_35_io_out ? io_r_52_b : _GEN_7171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7173 = 8'h35 == r_count_35_io_out ? io_r_53_b : _GEN_7172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7174 = 8'h36 == r_count_35_io_out ? io_r_54_b : _GEN_7173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7175 = 8'h37 == r_count_35_io_out ? io_r_55_b : _GEN_7174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7176 = 8'h38 == r_count_35_io_out ? io_r_56_b : _GEN_7175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7177 = 8'h39 == r_count_35_io_out ? io_r_57_b : _GEN_7176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7178 = 8'h3a == r_count_35_io_out ? io_r_58_b : _GEN_7177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7179 = 8'h3b == r_count_35_io_out ? io_r_59_b : _GEN_7178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7180 = 8'h3c == r_count_35_io_out ? io_r_60_b : _GEN_7179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7181 = 8'h3d == r_count_35_io_out ? io_r_61_b : _GEN_7180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7182 = 8'h3e == r_count_35_io_out ? io_r_62_b : _GEN_7181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7183 = 8'h3f == r_count_35_io_out ? io_r_63_b : _GEN_7182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7184 = 8'h40 == r_count_35_io_out ? io_r_64_b : _GEN_7183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7185 = 8'h41 == r_count_35_io_out ? io_r_65_b : _GEN_7184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7186 = 8'h42 == r_count_35_io_out ? io_r_66_b : _GEN_7185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7187 = 8'h43 == r_count_35_io_out ? io_r_67_b : _GEN_7186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7188 = 8'h44 == r_count_35_io_out ? io_r_68_b : _GEN_7187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7189 = 8'h45 == r_count_35_io_out ? io_r_69_b : _GEN_7188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7190 = 8'h46 == r_count_35_io_out ? io_r_70_b : _GEN_7189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7191 = 8'h47 == r_count_35_io_out ? io_r_71_b : _GEN_7190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7192 = 8'h48 == r_count_35_io_out ? io_r_72_b : _GEN_7191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7193 = 8'h49 == r_count_35_io_out ? io_r_73_b : _GEN_7192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7194 = 8'h4a == r_count_35_io_out ? io_r_74_b : _GEN_7193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7195 = 8'h4b == r_count_35_io_out ? io_r_75_b : _GEN_7194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7196 = 8'h4c == r_count_35_io_out ? io_r_76_b : _GEN_7195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7197 = 8'h4d == r_count_35_io_out ? io_r_77_b : _GEN_7196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7198 = 8'h4e == r_count_35_io_out ? io_r_78_b : _GEN_7197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7199 = 8'h4f == r_count_35_io_out ? io_r_79_b : _GEN_7198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7200 = 8'h50 == r_count_35_io_out ? io_r_80_b : _GEN_7199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7201 = 8'h51 == r_count_35_io_out ? io_r_81_b : _GEN_7200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7202 = 8'h52 == r_count_35_io_out ? io_r_82_b : _GEN_7201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7203 = 8'h53 == r_count_35_io_out ? io_r_83_b : _GEN_7202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7204 = 8'h54 == r_count_35_io_out ? io_r_84_b : _GEN_7203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7205 = 8'h55 == r_count_35_io_out ? io_r_85_b : _GEN_7204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7206 = 8'h56 == r_count_35_io_out ? io_r_86_b : _GEN_7205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7207 = 8'h57 == r_count_35_io_out ? io_r_87_b : _GEN_7206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7208 = 8'h58 == r_count_35_io_out ? io_r_88_b : _GEN_7207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7209 = 8'h59 == r_count_35_io_out ? io_r_89_b : _GEN_7208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7210 = 8'h5a == r_count_35_io_out ? io_r_90_b : _GEN_7209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7211 = 8'h5b == r_count_35_io_out ? io_r_91_b : _GEN_7210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7212 = 8'h5c == r_count_35_io_out ? io_r_92_b : _GEN_7211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7213 = 8'h5d == r_count_35_io_out ? io_r_93_b : _GEN_7212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7214 = 8'h5e == r_count_35_io_out ? io_r_94_b : _GEN_7213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7215 = 8'h5f == r_count_35_io_out ? io_r_95_b : _GEN_7214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7216 = 8'h60 == r_count_35_io_out ? io_r_96_b : _GEN_7215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7217 = 8'h61 == r_count_35_io_out ? io_r_97_b : _GEN_7216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7218 = 8'h62 == r_count_35_io_out ? io_r_98_b : _GEN_7217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7219 = 8'h63 == r_count_35_io_out ? io_r_99_b : _GEN_7218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7220 = 8'h64 == r_count_35_io_out ? io_r_100_b : _GEN_7219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7221 = 8'h65 == r_count_35_io_out ? io_r_101_b : _GEN_7220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7222 = 8'h66 == r_count_35_io_out ? io_r_102_b : _GEN_7221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7223 = 8'h67 == r_count_35_io_out ? io_r_103_b : _GEN_7222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7224 = 8'h68 == r_count_35_io_out ? io_r_104_b : _GEN_7223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7225 = 8'h69 == r_count_35_io_out ? io_r_105_b : _GEN_7224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7226 = 8'h6a == r_count_35_io_out ? io_r_106_b : _GEN_7225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7227 = 8'h6b == r_count_35_io_out ? io_r_107_b : _GEN_7226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7228 = 8'h6c == r_count_35_io_out ? io_r_108_b : _GEN_7227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7229 = 8'h6d == r_count_35_io_out ? io_r_109_b : _GEN_7228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7230 = 8'h6e == r_count_35_io_out ? io_r_110_b : _GEN_7229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7231 = 8'h6f == r_count_35_io_out ? io_r_111_b : _GEN_7230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7232 = 8'h70 == r_count_35_io_out ? io_r_112_b : _GEN_7231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7233 = 8'h71 == r_count_35_io_out ? io_r_113_b : _GEN_7232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7234 = 8'h72 == r_count_35_io_out ? io_r_114_b : _GEN_7233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7235 = 8'h73 == r_count_35_io_out ? io_r_115_b : _GEN_7234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7236 = 8'h74 == r_count_35_io_out ? io_r_116_b : _GEN_7235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7237 = 8'h75 == r_count_35_io_out ? io_r_117_b : _GEN_7236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7238 = 8'h76 == r_count_35_io_out ? io_r_118_b : _GEN_7237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7239 = 8'h77 == r_count_35_io_out ? io_r_119_b : _GEN_7238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7240 = 8'h78 == r_count_35_io_out ? io_r_120_b : _GEN_7239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7241 = 8'h79 == r_count_35_io_out ? io_r_121_b : _GEN_7240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7242 = 8'h7a == r_count_35_io_out ? io_r_122_b : _GEN_7241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7243 = 8'h7b == r_count_35_io_out ? io_r_123_b : _GEN_7242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7244 = 8'h7c == r_count_35_io_out ? io_r_124_b : _GEN_7243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7245 = 8'h7d == r_count_35_io_out ? io_r_125_b : _GEN_7244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7246 = 8'h7e == r_count_35_io_out ? io_r_126_b : _GEN_7245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7247 = 8'h7f == r_count_35_io_out ? io_r_127_b : _GEN_7246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7248 = 8'h80 == r_count_35_io_out ? io_r_128_b : _GEN_7247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7249 = 8'h81 == r_count_35_io_out ? io_r_129_b : _GEN_7248; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7250 = 8'h82 == r_count_35_io_out ? io_r_130_b : _GEN_7249; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7251 = 8'h83 == r_count_35_io_out ? io_r_131_b : _GEN_7250; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7252 = 8'h84 == r_count_35_io_out ? io_r_132_b : _GEN_7251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7253 = 8'h85 == r_count_35_io_out ? io_r_133_b : _GEN_7252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7254 = 8'h86 == r_count_35_io_out ? io_r_134_b : _GEN_7253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7255 = 8'h87 == r_count_35_io_out ? io_r_135_b : _GEN_7254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7256 = 8'h88 == r_count_35_io_out ? io_r_136_b : _GEN_7255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7257 = 8'h89 == r_count_35_io_out ? io_r_137_b : _GEN_7256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7258 = 8'h8a == r_count_35_io_out ? io_r_138_b : _GEN_7257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7259 = 8'h8b == r_count_35_io_out ? io_r_139_b : _GEN_7258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7260 = 8'h8c == r_count_35_io_out ? io_r_140_b : _GEN_7259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7261 = 8'h8d == r_count_35_io_out ? io_r_141_b : _GEN_7260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7262 = 8'h8e == r_count_35_io_out ? io_r_142_b : _GEN_7261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7263 = 8'h8f == r_count_35_io_out ? io_r_143_b : _GEN_7262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7264 = 8'h90 == r_count_35_io_out ? io_r_144_b : _GEN_7263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7265 = 8'h91 == r_count_35_io_out ? io_r_145_b : _GEN_7264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7266 = 8'h92 == r_count_35_io_out ? io_r_146_b : _GEN_7265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7267 = 8'h93 == r_count_35_io_out ? io_r_147_b : _GEN_7266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7268 = 8'h94 == r_count_35_io_out ? io_r_148_b : _GEN_7267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7269 = 8'h95 == r_count_35_io_out ? io_r_149_b : _GEN_7268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7270 = 8'h96 == r_count_35_io_out ? io_r_150_b : _GEN_7269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7271 = 8'h97 == r_count_35_io_out ? io_r_151_b : _GEN_7270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7272 = 8'h98 == r_count_35_io_out ? io_r_152_b : _GEN_7271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7273 = 8'h99 == r_count_35_io_out ? io_r_153_b : _GEN_7272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7274 = 8'h9a == r_count_35_io_out ? io_r_154_b : _GEN_7273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7275 = 8'h9b == r_count_35_io_out ? io_r_155_b : _GEN_7274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7276 = 8'h9c == r_count_35_io_out ? io_r_156_b : _GEN_7275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7277 = 8'h9d == r_count_35_io_out ? io_r_157_b : _GEN_7276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7278 = 8'h9e == r_count_35_io_out ? io_r_158_b : _GEN_7277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7279 = 8'h9f == r_count_35_io_out ? io_r_159_b : _GEN_7278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7280 = 8'ha0 == r_count_35_io_out ? io_r_160_b : _GEN_7279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7281 = 8'ha1 == r_count_35_io_out ? io_r_161_b : _GEN_7280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7282 = 8'ha2 == r_count_35_io_out ? io_r_162_b : _GEN_7281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7283 = 8'ha3 == r_count_35_io_out ? io_r_163_b : _GEN_7282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7284 = 8'ha4 == r_count_35_io_out ? io_r_164_b : _GEN_7283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7285 = 8'ha5 == r_count_35_io_out ? io_r_165_b : _GEN_7284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7286 = 8'ha6 == r_count_35_io_out ? io_r_166_b : _GEN_7285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7287 = 8'ha7 == r_count_35_io_out ? io_r_167_b : _GEN_7286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7288 = 8'ha8 == r_count_35_io_out ? io_r_168_b : _GEN_7287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7289 = 8'ha9 == r_count_35_io_out ? io_r_169_b : _GEN_7288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7290 = 8'haa == r_count_35_io_out ? io_r_170_b : _GEN_7289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7291 = 8'hab == r_count_35_io_out ? io_r_171_b : _GEN_7290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7292 = 8'hac == r_count_35_io_out ? io_r_172_b : _GEN_7291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7293 = 8'had == r_count_35_io_out ? io_r_173_b : _GEN_7292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7294 = 8'hae == r_count_35_io_out ? io_r_174_b : _GEN_7293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7295 = 8'haf == r_count_35_io_out ? io_r_175_b : _GEN_7294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7296 = 8'hb0 == r_count_35_io_out ? io_r_176_b : _GEN_7295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7297 = 8'hb1 == r_count_35_io_out ? io_r_177_b : _GEN_7296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7298 = 8'hb2 == r_count_35_io_out ? io_r_178_b : _GEN_7297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7299 = 8'hb3 == r_count_35_io_out ? io_r_179_b : _GEN_7298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7300 = 8'hb4 == r_count_35_io_out ? io_r_180_b : _GEN_7299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7301 = 8'hb5 == r_count_35_io_out ? io_r_181_b : _GEN_7300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7302 = 8'hb6 == r_count_35_io_out ? io_r_182_b : _GEN_7301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7303 = 8'hb7 == r_count_35_io_out ? io_r_183_b : _GEN_7302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7304 = 8'hb8 == r_count_35_io_out ? io_r_184_b : _GEN_7303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7305 = 8'hb9 == r_count_35_io_out ? io_r_185_b : _GEN_7304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7306 = 8'hba == r_count_35_io_out ? io_r_186_b : _GEN_7305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7307 = 8'hbb == r_count_35_io_out ? io_r_187_b : _GEN_7306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7308 = 8'hbc == r_count_35_io_out ? io_r_188_b : _GEN_7307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7309 = 8'hbd == r_count_35_io_out ? io_r_189_b : _GEN_7308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7310 = 8'hbe == r_count_35_io_out ? io_r_190_b : _GEN_7309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7311 = 8'hbf == r_count_35_io_out ? io_r_191_b : _GEN_7310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7312 = 8'hc0 == r_count_35_io_out ? io_r_192_b : _GEN_7311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7313 = 8'hc1 == r_count_35_io_out ? io_r_193_b : _GEN_7312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7314 = 8'hc2 == r_count_35_io_out ? io_r_194_b : _GEN_7313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7315 = 8'hc3 == r_count_35_io_out ? io_r_195_b : _GEN_7314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7316 = 8'hc4 == r_count_35_io_out ? io_r_196_b : _GEN_7315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7317 = 8'hc5 == r_count_35_io_out ? io_r_197_b : _GEN_7316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7318 = 8'hc6 == r_count_35_io_out ? io_r_198_b : _GEN_7317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7321 = 8'h1 == r_count_36_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7322 = 8'h2 == r_count_36_io_out ? io_r_2_b : _GEN_7321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7323 = 8'h3 == r_count_36_io_out ? io_r_3_b : _GEN_7322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7324 = 8'h4 == r_count_36_io_out ? io_r_4_b : _GEN_7323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7325 = 8'h5 == r_count_36_io_out ? io_r_5_b : _GEN_7324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7326 = 8'h6 == r_count_36_io_out ? io_r_6_b : _GEN_7325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7327 = 8'h7 == r_count_36_io_out ? io_r_7_b : _GEN_7326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7328 = 8'h8 == r_count_36_io_out ? io_r_8_b : _GEN_7327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7329 = 8'h9 == r_count_36_io_out ? io_r_9_b : _GEN_7328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7330 = 8'ha == r_count_36_io_out ? io_r_10_b : _GEN_7329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7331 = 8'hb == r_count_36_io_out ? io_r_11_b : _GEN_7330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7332 = 8'hc == r_count_36_io_out ? io_r_12_b : _GEN_7331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7333 = 8'hd == r_count_36_io_out ? io_r_13_b : _GEN_7332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7334 = 8'he == r_count_36_io_out ? io_r_14_b : _GEN_7333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7335 = 8'hf == r_count_36_io_out ? io_r_15_b : _GEN_7334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7336 = 8'h10 == r_count_36_io_out ? io_r_16_b : _GEN_7335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7337 = 8'h11 == r_count_36_io_out ? io_r_17_b : _GEN_7336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7338 = 8'h12 == r_count_36_io_out ? io_r_18_b : _GEN_7337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7339 = 8'h13 == r_count_36_io_out ? io_r_19_b : _GEN_7338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7340 = 8'h14 == r_count_36_io_out ? io_r_20_b : _GEN_7339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7341 = 8'h15 == r_count_36_io_out ? io_r_21_b : _GEN_7340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7342 = 8'h16 == r_count_36_io_out ? io_r_22_b : _GEN_7341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7343 = 8'h17 == r_count_36_io_out ? io_r_23_b : _GEN_7342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7344 = 8'h18 == r_count_36_io_out ? io_r_24_b : _GEN_7343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7345 = 8'h19 == r_count_36_io_out ? io_r_25_b : _GEN_7344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7346 = 8'h1a == r_count_36_io_out ? io_r_26_b : _GEN_7345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7347 = 8'h1b == r_count_36_io_out ? io_r_27_b : _GEN_7346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7348 = 8'h1c == r_count_36_io_out ? io_r_28_b : _GEN_7347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7349 = 8'h1d == r_count_36_io_out ? io_r_29_b : _GEN_7348; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7350 = 8'h1e == r_count_36_io_out ? io_r_30_b : _GEN_7349; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7351 = 8'h1f == r_count_36_io_out ? io_r_31_b : _GEN_7350; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7352 = 8'h20 == r_count_36_io_out ? io_r_32_b : _GEN_7351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7353 = 8'h21 == r_count_36_io_out ? io_r_33_b : _GEN_7352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7354 = 8'h22 == r_count_36_io_out ? io_r_34_b : _GEN_7353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7355 = 8'h23 == r_count_36_io_out ? io_r_35_b : _GEN_7354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7356 = 8'h24 == r_count_36_io_out ? io_r_36_b : _GEN_7355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7357 = 8'h25 == r_count_36_io_out ? io_r_37_b : _GEN_7356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7358 = 8'h26 == r_count_36_io_out ? io_r_38_b : _GEN_7357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7359 = 8'h27 == r_count_36_io_out ? io_r_39_b : _GEN_7358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7360 = 8'h28 == r_count_36_io_out ? io_r_40_b : _GEN_7359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7361 = 8'h29 == r_count_36_io_out ? io_r_41_b : _GEN_7360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7362 = 8'h2a == r_count_36_io_out ? io_r_42_b : _GEN_7361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7363 = 8'h2b == r_count_36_io_out ? io_r_43_b : _GEN_7362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7364 = 8'h2c == r_count_36_io_out ? io_r_44_b : _GEN_7363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7365 = 8'h2d == r_count_36_io_out ? io_r_45_b : _GEN_7364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7366 = 8'h2e == r_count_36_io_out ? io_r_46_b : _GEN_7365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7367 = 8'h2f == r_count_36_io_out ? io_r_47_b : _GEN_7366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7368 = 8'h30 == r_count_36_io_out ? io_r_48_b : _GEN_7367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7369 = 8'h31 == r_count_36_io_out ? io_r_49_b : _GEN_7368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7370 = 8'h32 == r_count_36_io_out ? io_r_50_b : _GEN_7369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7371 = 8'h33 == r_count_36_io_out ? io_r_51_b : _GEN_7370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7372 = 8'h34 == r_count_36_io_out ? io_r_52_b : _GEN_7371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7373 = 8'h35 == r_count_36_io_out ? io_r_53_b : _GEN_7372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7374 = 8'h36 == r_count_36_io_out ? io_r_54_b : _GEN_7373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7375 = 8'h37 == r_count_36_io_out ? io_r_55_b : _GEN_7374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7376 = 8'h38 == r_count_36_io_out ? io_r_56_b : _GEN_7375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7377 = 8'h39 == r_count_36_io_out ? io_r_57_b : _GEN_7376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7378 = 8'h3a == r_count_36_io_out ? io_r_58_b : _GEN_7377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7379 = 8'h3b == r_count_36_io_out ? io_r_59_b : _GEN_7378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7380 = 8'h3c == r_count_36_io_out ? io_r_60_b : _GEN_7379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7381 = 8'h3d == r_count_36_io_out ? io_r_61_b : _GEN_7380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7382 = 8'h3e == r_count_36_io_out ? io_r_62_b : _GEN_7381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7383 = 8'h3f == r_count_36_io_out ? io_r_63_b : _GEN_7382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7384 = 8'h40 == r_count_36_io_out ? io_r_64_b : _GEN_7383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7385 = 8'h41 == r_count_36_io_out ? io_r_65_b : _GEN_7384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7386 = 8'h42 == r_count_36_io_out ? io_r_66_b : _GEN_7385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7387 = 8'h43 == r_count_36_io_out ? io_r_67_b : _GEN_7386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7388 = 8'h44 == r_count_36_io_out ? io_r_68_b : _GEN_7387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7389 = 8'h45 == r_count_36_io_out ? io_r_69_b : _GEN_7388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7390 = 8'h46 == r_count_36_io_out ? io_r_70_b : _GEN_7389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7391 = 8'h47 == r_count_36_io_out ? io_r_71_b : _GEN_7390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7392 = 8'h48 == r_count_36_io_out ? io_r_72_b : _GEN_7391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7393 = 8'h49 == r_count_36_io_out ? io_r_73_b : _GEN_7392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7394 = 8'h4a == r_count_36_io_out ? io_r_74_b : _GEN_7393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7395 = 8'h4b == r_count_36_io_out ? io_r_75_b : _GEN_7394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7396 = 8'h4c == r_count_36_io_out ? io_r_76_b : _GEN_7395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7397 = 8'h4d == r_count_36_io_out ? io_r_77_b : _GEN_7396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7398 = 8'h4e == r_count_36_io_out ? io_r_78_b : _GEN_7397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7399 = 8'h4f == r_count_36_io_out ? io_r_79_b : _GEN_7398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7400 = 8'h50 == r_count_36_io_out ? io_r_80_b : _GEN_7399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7401 = 8'h51 == r_count_36_io_out ? io_r_81_b : _GEN_7400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7402 = 8'h52 == r_count_36_io_out ? io_r_82_b : _GEN_7401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7403 = 8'h53 == r_count_36_io_out ? io_r_83_b : _GEN_7402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7404 = 8'h54 == r_count_36_io_out ? io_r_84_b : _GEN_7403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7405 = 8'h55 == r_count_36_io_out ? io_r_85_b : _GEN_7404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7406 = 8'h56 == r_count_36_io_out ? io_r_86_b : _GEN_7405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7407 = 8'h57 == r_count_36_io_out ? io_r_87_b : _GEN_7406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7408 = 8'h58 == r_count_36_io_out ? io_r_88_b : _GEN_7407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7409 = 8'h59 == r_count_36_io_out ? io_r_89_b : _GEN_7408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7410 = 8'h5a == r_count_36_io_out ? io_r_90_b : _GEN_7409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7411 = 8'h5b == r_count_36_io_out ? io_r_91_b : _GEN_7410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7412 = 8'h5c == r_count_36_io_out ? io_r_92_b : _GEN_7411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7413 = 8'h5d == r_count_36_io_out ? io_r_93_b : _GEN_7412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7414 = 8'h5e == r_count_36_io_out ? io_r_94_b : _GEN_7413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7415 = 8'h5f == r_count_36_io_out ? io_r_95_b : _GEN_7414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7416 = 8'h60 == r_count_36_io_out ? io_r_96_b : _GEN_7415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7417 = 8'h61 == r_count_36_io_out ? io_r_97_b : _GEN_7416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7418 = 8'h62 == r_count_36_io_out ? io_r_98_b : _GEN_7417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7419 = 8'h63 == r_count_36_io_out ? io_r_99_b : _GEN_7418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7420 = 8'h64 == r_count_36_io_out ? io_r_100_b : _GEN_7419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7421 = 8'h65 == r_count_36_io_out ? io_r_101_b : _GEN_7420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7422 = 8'h66 == r_count_36_io_out ? io_r_102_b : _GEN_7421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7423 = 8'h67 == r_count_36_io_out ? io_r_103_b : _GEN_7422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7424 = 8'h68 == r_count_36_io_out ? io_r_104_b : _GEN_7423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7425 = 8'h69 == r_count_36_io_out ? io_r_105_b : _GEN_7424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7426 = 8'h6a == r_count_36_io_out ? io_r_106_b : _GEN_7425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7427 = 8'h6b == r_count_36_io_out ? io_r_107_b : _GEN_7426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7428 = 8'h6c == r_count_36_io_out ? io_r_108_b : _GEN_7427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7429 = 8'h6d == r_count_36_io_out ? io_r_109_b : _GEN_7428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7430 = 8'h6e == r_count_36_io_out ? io_r_110_b : _GEN_7429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7431 = 8'h6f == r_count_36_io_out ? io_r_111_b : _GEN_7430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7432 = 8'h70 == r_count_36_io_out ? io_r_112_b : _GEN_7431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7433 = 8'h71 == r_count_36_io_out ? io_r_113_b : _GEN_7432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7434 = 8'h72 == r_count_36_io_out ? io_r_114_b : _GEN_7433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7435 = 8'h73 == r_count_36_io_out ? io_r_115_b : _GEN_7434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7436 = 8'h74 == r_count_36_io_out ? io_r_116_b : _GEN_7435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7437 = 8'h75 == r_count_36_io_out ? io_r_117_b : _GEN_7436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7438 = 8'h76 == r_count_36_io_out ? io_r_118_b : _GEN_7437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7439 = 8'h77 == r_count_36_io_out ? io_r_119_b : _GEN_7438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7440 = 8'h78 == r_count_36_io_out ? io_r_120_b : _GEN_7439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7441 = 8'h79 == r_count_36_io_out ? io_r_121_b : _GEN_7440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7442 = 8'h7a == r_count_36_io_out ? io_r_122_b : _GEN_7441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7443 = 8'h7b == r_count_36_io_out ? io_r_123_b : _GEN_7442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7444 = 8'h7c == r_count_36_io_out ? io_r_124_b : _GEN_7443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7445 = 8'h7d == r_count_36_io_out ? io_r_125_b : _GEN_7444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7446 = 8'h7e == r_count_36_io_out ? io_r_126_b : _GEN_7445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7447 = 8'h7f == r_count_36_io_out ? io_r_127_b : _GEN_7446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7448 = 8'h80 == r_count_36_io_out ? io_r_128_b : _GEN_7447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7449 = 8'h81 == r_count_36_io_out ? io_r_129_b : _GEN_7448; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7450 = 8'h82 == r_count_36_io_out ? io_r_130_b : _GEN_7449; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7451 = 8'h83 == r_count_36_io_out ? io_r_131_b : _GEN_7450; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7452 = 8'h84 == r_count_36_io_out ? io_r_132_b : _GEN_7451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7453 = 8'h85 == r_count_36_io_out ? io_r_133_b : _GEN_7452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7454 = 8'h86 == r_count_36_io_out ? io_r_134_b : _GEN_7453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7455 = 8'h87 == r_count_36_io_out ? io_r_135_b : _GEN_7454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7456 = 8'h88 == r_count_36_io_out ? io_r_136_b : _GEN_7455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7457 = 8'h89 == r_count_36_io_out ? io_r_137_b : _GEN_7456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7458 = 8'h8a == r_count_36_io_out ? io_r_138_b : _GEN_7457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7459 = 8'h8b == r_count_36_io_out ? io_r_139_b : _GEN_7458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7460 = 8'h8c == r_count_36_io_out ? io_r_140_b : _GEN_7459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7461 = 8'h8d == r_count_36_io_out ? io_r_141_b : _GEN_7460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7462 = 8'h8e == r_count_36_io_out ? io_r_142_b : _GEN_7461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7463 = 8'h8f == r_count_36_io_out ? io_r_143_b : _GEN_7462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7464 = 8'h90 == r_count_36_io_out ? io_r_144_b : _GEN_7463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7465 = 8'h91 == r_count_36_io_out ? io_r_145_b : _GEN_7464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7466 = 8'h92 == r_count_36_io_out ? io_r_146_b : _GEN_7465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7467 = 8'h93 == r_count_36_io_out ? io_r_147_b : _GEN_7466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7468 = 8'h94 == r_count_36_io_out ? io_r_148_b : _GEN_7467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7469 = 8'h95 == r_count_36_io_out ? io_r_149_b : _GEN_7468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7470 = 8'h96 == r_count_36_io_out ? io_r_150_b : _GEN_7469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7471 = 8'h97 == r_count_36_io_out ? io_r_151_b : _GEN_7470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7472 = 8'h98 == r_count_36_io_out ? io_r_152_b : _GEN_7471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7473 = 8'h99 == r_count_36_io_out ? io_r_153_b : _GEN_7472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7474 = 8'h9a == r_count_36_io_out ? io_r_154_b : _GEN_7473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7475 = 8'h9b == r_count_36_io_out ? io_r_155_b : _GEN_7474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7476 = 8'h9c == r_count_36_io_out ? io_r_156_b : _GEN_7475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7477 = 8'h9d == r_count_36_io_out ? io_r_157_b : _GEN_7476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7478 = 8'h9e == r_count_36_io_out ? io_r_158_b : _GEN_7477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7479 = 8'h9f == r_count_36_io_out ? io_r_159_b : _GEN_7478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7480 = 8'ha0 == r_count_36_io_out ? io_r_160_b : _GEN_7479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7481 = 8'ha1 == r_count_36_io_out ? io_r_161_b : _GEN_7480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7482 = 8'ha2 == r_count_36_io_out ? io_r_162_b : _GEN_7481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7483 = 8'ha3 == r_count_36_io_out ? io_r_163_b : _GEN_7482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7484 = 8'ha4 == r_count_36_io_out ? io_r_164_b : _GEN_7483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7485 = 8'ha5 == r_count_36_io_out ? io_r_165_b : _GEN_7484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7486 = 8'ha6 == r_count_36_io_out ? io_r_166_b : _GEN_7485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7487 = 8'ha7 == r_count_36_io_out ? io_r_167_b : _GEN_7486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7488 = 8'ha8 == r_count_36_io_out ? io_r_168_b : _GEN_7487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7489 = 8'ha9 == r_count_36_io_out ? io_r_169_b : _GEN_7488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7490 = 8'haa == r_count_36_io_out ? io_r_170_b : _GEN_7489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7491 = 8'hab == r_count_36_io_out ? io_r_171_b : _GEN_7490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7492 = 8'hac == r_count_36_io_out ? io_r_172_b : _GEN_7491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7493 = 8'had == r_count_36_io_out ? io_r_173_b : _GEN_7492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7494 = 8'hae == r_count_36_io_out ? io_r_174_b : _GEN_7493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7495 = 8'haf == r_count_36_io_out ? io_r_175_b : _GEN_7494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7496 = 8'hb0 == r_count_36_io_out ? io_r_176_b : _GEN_7495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7497 = 8'hb1 == r_count_36_io_out ? io_r_177_b : _GEN_7496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7498 = 8'hb2 == r_count_36_io_out ? io_r_178_b : _GEN_7497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7499 = 8'hb3 == r_count_36_io_out ? io_r_179_b : _GEN_7498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7500 = 8'hb4 == r_count_36_io_out ? io_r_180_b : _GEN_7499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7501 = 8'hb5 == r_count_36_io_out ? io_r_181_b : _GEN_7500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7502 = 8'hb6 == r_count_36_io_out ? io_r_182_b : _GEN_7501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7503 = 8'hb7 == r_count_36_io_out ? io_r_183_b : _GEN_7502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7504 = 8'hb8 == r_count_36_io_out ? io_r_184_b : _GEN_7503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7505 = 8'hb9 == r_count_36_io_out ? io_r_185_b : _GEN_7504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7506 = 8'hba == r_count_36_io_out ? io_r_186_b : _GEN_7505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7507 = 8'hbb == r_count_36_io_out ? io_r_187_b : _GEN_7506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7508 = 8'hbc == r_count_36_io_out ? io_r_188_b : _GEN_7507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7509 = 8'hbd == r_count_36_io_out ? io_r_189_b : _GEN_7508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7510 = 8'hbe == r_count_36_io_out ? io_r_190_b : _GEN_7509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7511 = 8'hbf == r_count_36_io_out ? io_r_191_b : _GEN_7510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7512 = 8'hc0 == r_count_36_io_out ? io_r_192_b : _GEN_7511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7513 = 8'hc1 == r_count_36_io_out ? io_r_193_b : _GEN_7512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7514 = 8'hc2 == r_count_36_io_out ? io_r_194_b : _GEN_7513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7515 = 8'hc3 == r_count_36_io_out ? io_r_195_b : _GEN_7514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7516 = 8'hc4 == r_count_36_io_out ? io_r_196_b : _GEN_7515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7517 = 8'hc5 == r_count_36_io_out ? io_r_197_b : _GEN_7516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7518 = 8'hc6 == r_count_36_io_out ? io_r_198_b : _GEN_7517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7521 = 8'h1 == r_count_37_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7522 = 8'h2 == r_count_37_io_out ? io_r_2_b : _GEN_7521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7523 = 8'h3 == r_count_37_io_out ? io_r_3_b : _GEN_7522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7524 = 8'h4 == r_count_37_io_out ? io_r_4_b : _GEN_7523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7525 = 8'h5 == r_count_37_io_out ? io_r_5_b : _GEN_7524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7526 = 8'h6 == r_count_37_io_out ? io_r_6_b : _GEN_7525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7527 = 8'h7 == r_count_37_io_out ? io_r_7_b : _GEN_7526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7528 = 8'h8 == r_count_37_io_out ? io_r_8_b : _GEN_7527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7529 = 8'h9 == r_count_37_io_out ? io_r_9_b : _GEN_7528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7530 = 8'ha == r_count_37_io_out ? io_r_10_b : _GEN_7529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7531 = 8'hb == r_count_37_io_out ? io_r_11_b : _GEN_7530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7532 = 8'hc == r_count_37_io_out ? io_r_12_b : _GEN_7531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7533 = 8'hd == r_count_37_io_out ? io_r_13_b : _GEN_7532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7534 = 8'he == r_count_37_io_out ? io_r_14_b : _GEN_7533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7535 = 8'hf == r_count_37_io_out ? io_r_15_b : _GEN_7534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7536 = 8'h10 == r_count_37_io_out ? io_r_16_b : _GEN_7535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7537 = 8'h11 == r_count_37_io_out ? io_r_17_b : _GEN_7536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7538 = 8'h12 == r_count_37_io_out ? io_r_18_b : _GEN_7537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7539 = 8'h13 == r_count_37_io_out ? io_r_19_b : _GEN_7538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7540 = 8'h14 == r_count_37_io_out ? io_r_20_b : _GEN_7539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7541 = 8'h15 == r_count_37_io_out ? io_r_21_b : _GEN_7540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7542 = 8'h16 == r_count_37_io_out ? io_r_22_b : _GEN_7541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7543 = 8'h17 == r_count_37_io_out ? io_r_23_b : _GEN_7542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7544 = 8'h18 == r_count_37_io_out ? io_r_24_b : _GEN_7543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7545 = 8'h19 == r_count_37_io_out ? io_r_25_b : _GEN_7544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7546 = 8'h1a == r_count_37_io_out ? io_r_26_b : _GEN_7545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7547 = 8'h1b == r_count_37_io_out ? io_r_27_b : _GEN_7546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7548 = 8'h1c == r_count_37_io_out ? io_r_28_b : _GEN_7547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7549 = 8'h1d == r_count_37_io_out ? io_r_29_b : _GEN_7548; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7550 = 8'h1e == r_count_37_io_out ? io_r_30_b : _GEN_7549; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7551 = 8'h1f == r_count_37_io_out ? io_r_31_b : _GEN_7550; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7552 = 8'h20 == r_count_37_io_out ? io_r_32_b : _GEN_7551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7553 = 8'h21 == r_count_37_io_out ? io_r_33_b : _GEN_7552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7554 = 8'h22 == r_count_37_io_out ? io_r_34_b : _GEN_7553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7555 = 8'h23 == r_count_37_io_out ? io_r_35_b : _GEN_7554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7556 = 8'h24 == r_count_37_io_out ? io_r_36_b : _GEN_7555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7557 = 8'h25 == r_count_37_io_out ? io_r_37_b : _GEN_7556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7558 = 8'h26 == r_count_37_io_out ? io_r_38_b : _GEN_7557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7559 = 8'h27 == r_count_37_io_out ? io_r_39_b : _GEN_7558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7560 = 8'h28 == r_count_37_io_out ? io_r_40_b : _GEN_7559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7561 = 8'h29 == r_count_37_io_out ? io_r_41_b : _GEN_7560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7562 = 8'h2a == r_count_37_io_out ? io_r_42_b : _GEN_7561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7563 = 8'h2b == r_count_37_io_out ? io_r_43_b : _GEN_7562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7564 = 8'h2c == r_count_37_io_out ? io_r_44_b : _GEN_7563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7565 = 8'h2d == r_count_37_io_out ? io_r_45_b : _GEN_7564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7566 = 8'h2e == r_count_37_io_out ? io_r_46_b : _GEN_7565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7567 = 8'h2f == r_count_37_io_out ? io_r_47_b : _GEN_7566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7568 = 8'h30 == r_count_37_io_out ? io_r_48_b : _GEN_7567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7569 = 8'h31 == r_count_37_io_out ? io_r_49_b : _GEN_7568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7570 = 8'h32 == r_count_37_io_out ? io_r_50_b : _GEN_7569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7571 = 8'h33 == r_count_37_io_out ? io_r_51_b : _GEN_7570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7572 = 8'h34 == r_count_37_io_out ? io_r_52_b : _GEN_7571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7573 = 8'h35 == r_count_37_io_out ? io_r_53_b : _GEN_7572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7574 = 8'h36 == r_count_37_io_out ? io_r_54_b : _GEN_7573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7575 = 8'h37 == r_count_37_io_out ? io_r_55_b : _GEN_7574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7576 = 8'h38 == r_count_37_io_out ? io_r_56_b : _GEN_7575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7577 = 8'h39 == r_count_37_io_out ? io_r_57_b : _GEN_7576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7578 = 8'h3a == r_count_37_io_out ? io_r_58_b : _GEN_7577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7579 = 8'h3b == r_count_37_io_out ? io_r_59_b : _GEN_7578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7580 = 8'h3c == r_count_37_io_out ? io_r_60_b : _GEN_7579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7581 = 8'h3d == r_count_37_io_out ? io_r_61_b : _GEN_7580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7582 = 8'h3e == r_count_37_io_out ? io_r_62_b : _GEN_7581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7583 = 8'h3f == r_count_37_io_out ? io_r_63_b : _GEN_7582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7584 = 8'h40 == r_count_37_io_out ? io_r_64_b : _GEN_7583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7585 = 8'h41 == r_count_37_io_out ? io_r_65_b : _GEN_7584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7586 = 8'h42 == r_count_37_io_out ? io_r_66_b : _GEN_7585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7587 = 8'h43 == r_count_37_io_out ? io_r_67_b : _GEN_7586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7588 = 8'h44 == r_count_37_io_out ? io_r_68_b : _GEN_7587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7589 = 8'h45 == r_count_37_io_out ? io_r_69_b : _GEN_7588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7590 = 8'h46 == r_count_37_io_out ? io_r_70_b : _GEN_7589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7591 = 8'h47 == r_count_37_io_out ? io_r_71_b : _GEN_7590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7592 = 8'h48 == r_count_37_io_out ? io_r_72_b : _GEN_7591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7593 = 8'h49 == r_count_37_io_out ? io_r_73_b : _GEN_7592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7594 = 8'h4a == r_count_37_io_out ? io_r_74_b : _GEN_7593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7595 = 8'h4b == r_count_37_io_out ? io_r_75_b : _GEN_7594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7596 = 8'h4c == r_count_37_io_out ? io_r_76_b : _GEN_7595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7597 = 8'h4d == r_count_37_io_out ? io_r_77_b : _GEN_7596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7598 = 8'h4e == r_count_37_io_out ? io_r_78_b : _GEN_7597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7599 = 8'h4f == r_count_37_io_out ? io_r_79_b : _GEN_7598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7600 = 8'h50 == r_count_37_io_out ? io_r_80_b : _GEN_7599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7601 = 8'h51 == r_count_37_io_out ? io_r_81_b : _GEN_7600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7602 = 8'h52 == r_count_37_io_out ? io_r_82_b : _GEN_7601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7603 = 8'h53 == r_count_37_io_out ? io_r_83_b : _GEN_7602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7604 = 8'h54 == r_count_37_io_out ? io_r_84_b : _GEN_7603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7605 = 8'h55 == r_count_37_io_out ? io_r_85_b : _GEN_7604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7606 = 8'h56 == r_count_37_io_out ? io_r_86_b : _GEN_7605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7607 = 8'h57 == r_count_37_io_out ? io_r_87_b : _GEN_7606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7608 = 8'h58 == r_count_37_io_out ? io_r_88_b : _GEN_7607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7609 = 8'h59 == r_count_37_io_out ? io_r_89_b : _GEN_7608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7610 = 8'h5a == r_count_37_io_out ? io_r_90_b : _GEN_7609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7611 = 8'h5b == r_count_37_io_out ? io_r_91_b : _GEN_7610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7612 = 8'h5c == r_count_37_io_out ? io_r_92_b : _GEN_7611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7613 = 8'h5d == r_count_37_io_out ? io_r_93_b : _GEN_7612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7614 = 8'h5e == r_count_37_io_out ? io_r_94_b : _GEN_7613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7615 = 8'h5f == r_count_37_io_out ? io_r_95_b : _GEN_7614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7616 = 8'h60 == r_count_37_io_out ? io_r_96_b : _GEN_7615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7617 = 8'h61 == r_count_37_io_out ? io_r_97_b : _GEN_7616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7618 = 8'h62 == r_count_37_io_out ? io_r_98_b : _GEN_7617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7619 = 8'h63 == r_count_37_io_out ? io_r_99_b : _GEN_7618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7620 = 8'h64 == r_count_37_io_out ? io_r_100_b : _GEN_7619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7621 = 8'h65 == r_count_37_io_out ? io_r_101_b : _GEN_7620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7622 = 8'h66 == r_count_37_io_out ? io_r_102_b : _GEN_7621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7623 = 8'h67 == r_count_37_io_out ? io_r_103_b : _GEN_7622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7624 = 8'h68 == r_count_37_io_out ? io_r_104_b : _GEN_7623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7625 = 8'h69 == r_count_37_io_out ? io_r_105_b : _GEN_7624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7626 = 8'h6a == r_count_37_io_out ? io_r_106_b : _GEN_7625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7627 = 8'h6b == r_count_37_io_out ? io_r_107_b : _GEN_7626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7628 = 8'h6c == r_count_37_io_out ? io_r_108_b : _GEN_7627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7629 = 8'h6d == r_count_37_io_out ? io_r_109_b : _GEN_7628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7630 = 8'h6e == r_count_37_io_out ? io_r_110_b : _GEN_7629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7631 = 8'h6f == r_count_37_io_out ? io_r_111_b : _GEN_7630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7632 = 8'h70 == r_count_37_io_out ? io_r_112_b : _GEN_7631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7633 = 8'h71 == r_count_37_io_out ? io_r_113_b : _GEN_7632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7634 = 8'h72 == r_count_37_io_out ? io_r_114_b : _GEN_7633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7635 = 8'h73 == r_count_37_io_out ? io_r_115_b : _GEN_7634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7636 = 8'h74 == r_count_37_io_out ? io_r_116_b : _GEN_7635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7637 = 8'h75 == r_count_37_io_out ? io_r_117_b : _GEN_7636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7638 = 8'h76 == r_count_37_io_out ? io_r_118_b : _GEN_7637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7639 = 8'h77 == r_count_37_io_out ? io_r_119_b : _GEN_7638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7640 = 8'h78 == r_count_37_io_out ? io_r_120_b : _GEN_7639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7641 = 8'h79 == r_count_37_io_out ? io_r_121_b : _GEN_7640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7642 = 8'h7a == r_count_37_io_out ? io_r_122_b : _GEN_7641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7643 = 8'h7b == r_count_37_io_out ? io_r_123_b : _GEN_7642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7644 = 8'h7c == r_count_37_io_out ? io_r_124_b : _GEN_7643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7645 = 8'h7d == r_count_37_io_out ? io_r_125_b : _GEN_7644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7646 = 8'h7e == r_count_37_io_out ? io_r_126_b : _GEN_7645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7647 = 8'h7f == r_count_37_io_out ? io_r_127_b : _GEN_7646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7648 = 8'h80 == r_count_37_io_out ? io_r_128_b : _GEN_7647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7649 = 8'h81 == r_count_37_io_out ? io_r_129_b : _GEN_7648; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7650 = 8'h82 == r_count_37_io_out ? io_r_130_b : _GEN_7649; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7651 = 8'h83 == r_count_37_io_out ? io_r_131_b : _GEN_7650; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7652 = 8'h84 == r_count_37_io_out ? io_r_132_b : _GEN_7651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7653 = 8'h85 == r_count_37_io_out ? io_r_133_b : _GEN_7652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7654 = 8'h86 == r_count_37_io_out ? io_r_134_b : _GEN_7653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7655 = 8'h87 == r_count_37_io_out ? io_r_135_b : _GEN_7654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7656 = 8'h88 == r_count_37_io_out ? io_r_136_b : _GEN_7655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7657 = 8'h89 == r_count_37_io_out ? io_r_137_b : _GEN_7656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7658 = 8'h8a == r_count_37_io_out ? io_r_138_b : _GEN_7657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7659 = 8'h8b == r_count_37_io_out ? io_r_139_b : _GEN_7658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7660 = 8'h8c == r_count_37_io_out ? io_r_140_b : _GEN_7659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7661 = 8'h8d == r_count_37_io_out ? io_r_141_b : _GEN_7660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7662 = 8'h8e == r_count_37_io_out ? io_r_142_b : _GEN_7661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7663 = 8'h8f == r_count_37_io_out ? io_r_143_b : _GEN_7662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7664 = 8'h90 == r_count_37_io_out ? io_r_144_b : _GEN_7663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7665 = 8'h91 == r_count_37_io_out ? io_r_145_b : _GEN_7664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7666 = 8'h92 == r_count_37_io_out ? io_r_146_b : _GEN_7665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7667 = 8'h93 == r_count_37_io_out ? io_r_147_b : _GEN_7666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7668 = 8'h94 == r_count_37_io_out ? io_r_148_b : _GEN_7667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7669 = 8'h95 == r_count_37_io_out ? io_r_149_b : _GEN_7668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7670 = 8'h96 == r_count_37_io_out ? io_r_150_b : _GEN_7669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7671 = 8'h97 == r_count_37_io_out ? io_r_151_b : _GEN_7670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7672 = 8'h98 == r_count_37_io_out ? io_r_152_b : _GEN_7671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7673 = 8'h99 == r_count_37_io_out ? io_r_153_b : _GEN_7672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7674 = 8'h9a == r_count_37_io_out ? io_r_154_b : _GEN_7673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7675 = 8'h9b == r_count_37_io_out ? io_r_155_b : _GEN_7674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7676 = 8'h9c == r_count_37_io_out ? io_r_156_b : _GEN_7675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7677 = 8'h9d == r_count_37_io_out ? io_r_157_b : _GEN_7676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7678 = 8'h9e == r_count_37_io_out ? io_r_158_b : _GEN_7677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7679 = 8'h9f == r_count_37_io_out ? io_r_159_b : _GEN_7678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7680 = 8'ha0 == r_count_37_io_out ? io_r_160_b : _GEN_7679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7681 = 8'ha1 == r_count_37_io_out ? io_r_161_b : _GEN_7680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7682 = 8'ha2 == r_count_37_io_out ? io_r_162_b : _GEN_7681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7683 = 8'ha3 == r_count_37_io_out ? io_r_163_b : _GEN_7682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7684 = 8'ha4 == r_count_37_io_out ? io_r_164_b : _GEN_7683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7685 = 8'ha5 == r_count_37_io_out ? io_r_165_b : _GEN_7684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7686 = 8'ha6 == r_count_37_io_out ? io_r_166_b : _GEN_7685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7687 = 8'ha7 == r_count_37_io_out ? io_r_167_b : _GEN_7686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7688 = 8'ha8 == r_count_37_io_out ? io_r_168_b : _GEN_7687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7689 = 8'ha9 == r_count_37_io_out ? io_r_169_b : _GEN_7688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7690 = 8'haa == r_count_37_io_out ? io_r_170_b : _GEN_7689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7691 = 8'hab == r_count_37_io_out ? io_r_171_b : _GEN_7690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7692 = 8'hac == r_count_37_io_out ? io_r_172_b : _GEN_7691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7693 = 8'had == r_count_37_io_out ? io_r_173_b : _GEN_7692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7694 = 8'hae == r_count_37_io_out ? io_r_174_b : _GEN_7693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7695 = 8'haf == r_count_37_io_out ? io_r_175_b : _GEN_7694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7696 = 8'hb0 == r_count_37_io_out ? io_r_176_b : _GEN_7695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7697 = 8'hb1 == r_count_37_io_out ? io_r_177_b : _GEN_7696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7698 = 8'hb2 == r_count_37_io_out ? io_r_178_b : _GEN_7697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7699 = 8'hb3 == r_count_37_io_out ? io_r_179_b : _GEN_7698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7700 = 8'hb4 == r_count_37_io_out ? io_r_180_b : _GEN_7699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7701 = 8'hb5 == r_count_37_io_out ? io_r_181_b : _GEN_7700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7702 = 8'hb6 == r_count_37_io_out ? io_r_182_b : _GEN_7701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7703 = 8'hb7 == r_count_37_io_out ? io_r_183_b : _GEN_7702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7704 = 8'hb8 == r_count_37_io_out ? io_r_184_b : _GEN_7703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7705 = 8'hb9 == r_count_37_io_out ? io_r_185_b : _GEN_7704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7706 = 8'hba == r_count_37_io_out ? io_r_186_b : _GEN_7705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7707 = 8'hbb == r_count_37_io_out ? io_r_187_b : _GEN_7706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7708 = 8'hbc == r_count_37_io_out ? io_r_188_b : _GEN_7707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7709 = 8'hbd == r_count_37_io_out ? io_r_189_b : _GEN_7708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7710 = 8'hbe == r_count_37_io_out ? io_r_190_b : _GEN_7709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7711 = 8'hbf == r_count_37_io_out ? io_r_191_b : _GEN_7710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7712 = 8'hc0 == r_count_37_io_out ? io_r_192_b : _GEN_7711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7713 = 8'hc1 == r_count_37_io_out ? io_r_193_b : _GEN_7712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7714 = 8'hc2 == r_count_37_io_out ? io_r_194_b : _GEN_7713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7715 = 8'hc3 == r_count_37_io_out ? io_r_195_b : _GEN_7714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7716 = 8'hc4 == r_count_37_io_out ? io_r_196_b : _GEN_7715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7717 = 8'hc5 == r_count_37_io_out ? io_r_197_b : _GEN_7716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7718 = 8'hc6 == r_count_37_io_out ? io_r_198_b : _GEN_7717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7721 = 8'h1 == r_count_38_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7722 = 8'h2 == r_count_38_io_out ? io_r_2_b : _GEN_7721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7723 = 8'h3 == r_count_38_io_out ? io_r_3_b : _GEN_7722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7724 = 8'h4 == r_count_38_io_out ? io_r_4_b : _GEN_7723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7725 = 8'h5 == r_count_38_io_out ? io_r_5_b : _GEN_7724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7726 = 8'h6 == r_count_38_io_out ? io_r_6_b : _GEN_7725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7727 = 8'h7 == r_count_38_io_out ? io_r_7_b : _GEN_7726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7728 = 8'h8 == r_count_38_io_out ? io_r_8_b : _GEN_7727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7729 = 8'h9 == r_count_38_io_out ? io_r_9_b : _GEN_7728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7730 = 8'ha == r_count_38_io_out ? io_r_10_b : _GEN_7729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7731 = 8'hb == r_count_38_io_out ? io_r_11_b : _GEN_7730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7732 = 8'hc == r_count_38_io_out ? io_r_12_b : _GEN_7731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7733 = 8'hd == r_count_38_io_out ? io_r_13_b : _GEN_7732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7734 = 8'he == r_count_38_io_out ? io_r_14_b : _GEN_7733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7735 = 8'hf == r_count_38_io_out ? io_r_15_b : _GEN_7734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7736 = 8'h10 == r_count_38_io_out ? io_r_16_b : _GEN_7735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7737 = 8'h11 == r_count_38_io_out ? io_r_17_b : _GEN_7736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7738 = 8'h12 == r_count_38_io_out ? io_r_18_b : _GEN_7737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7739 = 8'h13 == r_count_38_io_out ? io_r_19_b : _GEN_7738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7740 = 8'h14 == r_count_38_io_out ? io_r_20_b : _GEN_7739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7741 = 8'h15 == r_count_38_io_out ? io_r_21_b : _GEN_7740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7742 = 8'h16 == r_count_38_io_out ? io_r_22_b : _GEN_7741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7743 = 8'h17 == r_count_38_io_out ? io_r_23_b : _GEN_7742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7744 = 8'h18 == r_count_38_io_out ? io_r_24_b : _GEN_7743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7745 = 8'h19 == r_count_38_io_out ? io_r_25_b : _GEN_7744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7746 = 8'h1a == r_count_38_io_out ? io_r_26_b : _GEN_7745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7747 = 8'h1b == r_count_38_io_out ? io_r_27_b : _GEN_7746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7748 = 8'h1c == r_count_38_io_out ? io_r_28_b : _GEN_7747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7749 = 8'h1d == r_count_38_io_out ? io_r_29_b : _GEN_7748; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7750 = 8'h1e == r_count_38_io_out ? io_r_30_b : _GEN_7749; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7751 = 8'h1f == r_count_38_io_out ? io_r_31_b : _GEN_7750; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7752 = 8'h20 == r_count_38_io_out ? io_r_32_b : _GEN_7751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7753 = 8'h21 == r_count_38_io_out ? io_r_33_b : _GEN_7752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7754 = 8'h22 == r_count_38_io_out ? io_r_34_b : _GEN_7753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7755 = 8'h23 == r_count_38_io_out ? io_r_35_b : _GEN_7754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7756 = 8'h24 == r_count_38_io_out ? io_r_36_b : _GEN_7755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7757 = 8'h25 == r_count_38_io_out ? io_r_37_b : _GEN_7756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7758 = 8'h26 == r_count_38_io_out ? io_r_38_b : _GEN_7757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7759 = 8'h27 == r_count_38_io_out ? io_r_39_b : _GEN_7758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7760 = 8'h28 == r_count_38_io_out ? io_r_40_b : _GEN_7759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7761 = 8'h29 == r_count_38_io_out ? io_r_41_b : _GEN_7760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7762 = 8'h2a == r_count_38_io_out ? io_r_42_b : _GEN_7761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7763 = 8'h2b == r_count_38_io_out ? io_r_43_b : _GEN_7762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7764 = 8'h2c == r_count_38_io_out ? io_r_44_b : _GEN_7763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7765 = 8'h2d == r_count_38_io_out ? io_r_45_b : _GEN_7764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7766 = 8'h2e == r_count_38_io_out ? io_r_46_b : _GEN_7765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7767 = 8'h2f == r_count_38_io_out ? io_r_47_b : _GEN_7766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7768 = 8'h30 == r_count_38_io_out ? io_r_48_b : _GEN_7767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7769 = 8'h31 == r_count_38_io_out ? io_r_49_b : _GEN_7768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7770 = 8'h32 == r_count_38_io_out ? io_r_50_b : _GEN_7769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7771 = 8'h33 == r_count_38_io_out ? io_r_51_b : _GEN_7770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7772 = 8'h34 == r_count_38_io_out ? io_r_52_b : _GEN_7771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7773 = 8'h35 == r_count_38_io_out ? io_r_53_b : _GEN_7772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7774 = 8'h36 == r_count_38_io_out ? io_r_54_b : _GEN_7773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7775 = 8'h37 == r_count_38_io_out ? io_r_55_b : _GEN_7774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7776 = 8'h38 == r_count_38_io_out ? io_r_56_b : _GEN_7775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7777 = 8'h39 == r_count_38_io_out ? io_r_57_b : _GEN_7776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7778 = 8'h3a == r_count_38_io_out ? io_r_58_b : _GEN_7777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7779 = 8'h3b == r_count_38_io_out ? io_r_59_b : _GEN_7778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7780 = 8'h3c == r_count_38_io_out ? io_r_60_b : _GEN_7779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7781 = 8'h3d == r_count_38_io_out ? io_r_61_b : _GEN_7780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7782 = 8'h3e == r_count_38_io_out ? io_r_62_b : _GEN_7781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7783 = 8'h3f == r_count_38_io_out ? io_r_63_b : _GEN_7782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7784 = 8'h40 == r_count_38_io_out ? io_r_64_b : _GEN_7783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7785 = 8'h41 == r_count_38_io_out ? io_r_65_b : _GEN_7784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7786 = 8'h42 == r_count_38_io_out ? io_r_66_b : _GEN_7785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7787 = 8'h43 == r_count_38_io_out ? io_r_67_b : _GEN_7786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7788 = 8'h44 == r_count_38_io_out ? io_r_68_b : _GEN_7787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7789 = 8'h45 == r_count_38_io_out ? io_r_69_b : _GEN_7788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7790 = 8'h46 == r_count_38_io_out ? io_r_70_b : _GEN_7789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7791 = 8'h47 == r_count_38_io_out ? io_r_71_b : _GEN_7790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7792 = 8'h48 == r_count_38_io_out ? io_r_72_b : _GEN_7791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7793 = 8'h49 == r_count_38_io_out ? io_r_73_b : _GEN_7792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7794 = 8'h4a == r_count_38_io_out ? io_r_74_b : _GEN_7793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7795 = 8'h4b == r_count_38_io_out ? io_r_75_b : _GEN_7794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7796 = 8'h4c == r_count_38_io_out ? io_r_76_b : _GEN_7795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7797 = 8'h4d == r_count_38_io_out ? io_r_77_b : _GEN_7796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7798 = 8'h4e == r_count_38_io_out ? io_r_78_b : _GEN_7797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7799 = 8'h4f == r_count_38_io_out ? io_r_79_b : _GEN_7798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7800 = 8'h50 == r_count_38_io_out ? io_r_80_b : _GEN_7799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7801 = 8'h51 == r_count_38_io_out ? io_r_81_b : _GEN_7800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7802 = 8'h52 == r_count_38_io_out ? io_r_82_b : _GEN_7801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7803 = 8'h53 == r_count_38_io_out ? io_r_83_b : _GEN_7802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7804 = 8'h54 == r_count_38_io_out ? io_r_84_b : _GEN_7803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7805 = 8'h55 == r_count_38_io_out ? io_r_85_b : _GEN_7804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7806 = 8'h56 == r_count_38_io_out ? io_r_86_b : _GEN_7805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7807 = 8'h57 == r_count_38_io_out ? io_r_87_b : _GEN_7806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7808 = 8'h58 == r_count_38_io_out ? io_r_88_b : _GEN_7807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7809 = 8'h59 == r_count_38_io_out ? io_r_89_b : _GEN_7808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7810 = 8'h5a == r_count_38_io_out ? io_r_90_b : _GEN_7809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7811 = 8'h5b == r_count_38_io_out ? io_r_91_b : _GEN_7810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7812 = 8'h5c == r_count_38_io_out ? io_r_92_b : _GEN_7811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7813 = 8'h5d == r_count_38_io_out ? io_r_93_b : _GEN_7812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7814 = 8'h5e == r_count_38_io_out ? io_r_94_b : _GEN_7813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7815 = 8'h5f == r_count_38_io_out ? io_r_95_b : _GEN_7814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7816 = 8'h60 == r_count_38_io_out ? io_r_96_b : _GEN_7815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7817 = 8'h61 == r_count_38_io_out ? io_r_97_b : _GEN_7816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7818 = 8'h62 == r_count_38_io_out ? io_r_98_b : _GEN_7817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7819 = 8'h63 == r_count_38_io_out ? io_r_99_b : _GEN_7818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7820 = 8'h64 == r_count_38_io_out ? io_r_100_b : _GEN_7819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7821 = 8'h65 == r_count_38_io_out ? io_r_101_b : _GEN_7820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7822 = 8'h66 == r_count_38_io_out ? io_r_102_b : _GEN_7821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7823 = 8'h67 == r_count_38_io_out ? io_r_103_b : _GEN_7822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7824 = 8'h68 == r_count_38_io_out ? io_r_104_b : _GEN_7823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7825 = 8'h69 == r_count_38_io_out ? io_r_105_b : _GEN_7824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7826 = 8'h6a == r_count_38_io_out ? io_r_106_b : _GEN_7825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7827 = 8'h6b == r_count_38_io_out ? io_r_107_b : _GEN_7826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7828 = 8'h6c == r_count_38_io_out ? io_r_108_b : _GEN_7827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7829 = 8'h6d == r_count_38_io_out ? io_r_109_b : _GEN_7828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7830 = 8'h6e == r_count_38_io_out ? io_r_110_b : _GEN_7829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7831 = 8'h6f == r_count_38_io_out ? io_r_111_b : _GEN_7830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7832 = 8'h70 == r_count_38_io_out ? io_r_112_b : _GEN_7831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7833 = 8'h71 == r_count_38_io_out ? io_r_113_b : _GEN_7832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7834 = 8'h72 == r_count_38_io_out ? io_r_114_b : _GEN_7833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7835 = 8'h73 == r_count_38_io_out ? io_r_115_b : _GEN_7834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7836 = 8'h74 == r_count_38_io_out ? io_r_116_b : _GEN_7835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7837 = 8'h75 == r_count_38_io_out ? io_r_117_b : _GEN_7836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7838 = 8'h76 == r_count_38_io_out ? io_r_118_b : _GEN_7837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7839 = 8'h77 == r_count_38_io_out ? io_r_119_b : _GEN_7838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7840 = 8'h78 == r_count_38_io_out ? io_r_120_b : _GEN_7839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7841 = 8'h79 == r_count_38_io_out ? io_r_121_b : _GEN_7840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7842 = 8'h7a == r_count_38_io_out ? io_r_122_b : _GEN_7841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7843 = 8'h7b == r_count_38_io_out ? io_r_123_b : _GEN_7842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7844 = 8'h7c == r_count_38_io_out ? io_r_124_b : _GEN_7843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7845 = 8'h7d == r_count_38_io_out ? io_r_125_b : _GEN_7844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7846 = 8'h7e == r_count_38_io_out ? io_r_126_b : _GEN_7845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7847 = 8'h7f == r_count_38_io_out ? io_r_127_b : _GEN_7846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7848 = 8'h80 == r_count_38_io_out ? io_r_128_b : _GEN_7847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7849 = 8'h81 == r_count_38_io_out ? io_r_129_b : _GEN_7848; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7850 = 8'h82 == r_count_38_io_out ? io_r_130_b : _GEN_7849; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7851 = 8'h83 == r_count_38_io_out ? io_r_131_b : _GEN_7850; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7852 = 8'h84 == r_count_38_io_out ? io_r_132_b : _GEN_7851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7853 = 8'h85 == r_count_38_io_out ? io_r_133_b : _GEN_7852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7854 = 8'h86 == r_count_38_io_out ? io_r_134_b : _GEN_7853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7855 = 8'h87 == r_count_38_io_out ? io_r_135_b : _GEN_7854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7856 = 8'h88 == r_count_38_io_out ? io_r_136_b : _GEN_7855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7857 = 8'h89 == r_count_38_io_out ? io_r_137_b : _GEN_7856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7858 = 8'h8a == r_count_38_io_out ? io_r_138_b : _GEN_7857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7859 = 8'h8b == r_count_38_io_out ? io_r_139_b : _GEN_7858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7860 = 8'h8c == r_count_38_io_out ? io_r_140_b : _GEN_7859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7861 = 8'h8d == r_count_38_io_out ? io_r_141_b : _GEN_7860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7862 = 8'h8e == r_count_38_io_out ? io_r_142_b : _GEN_7861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7863 = 8'h8f == r_count_38_io_out ? io_r_143_b : _GEN_7862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7864 = 8'h90 == r_count_38_io_out ? io_r_144_b : _GEN_7863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7865 = 8'h91 == r_count_38_io_out ? io_r_145_b : _GEN_7864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7866 = 8'h92 == r_count_38_io_out ? io_r_146_b : _GEN_7865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7867 = 8'h93 == r_count_38_io_out ? io_r_147_b : _GEN_7866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7868 = 8'h94 == r_count_38_io_out ? io_r_148_b : _GEN_7867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7869 = 8'h95 == r_count_38_io_out ? io_r_149_b : _GEN_7868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7870 = 8'h96 == r_count_38_io_out ? io_r_150_b : _GEN_7869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7871 = 8'h97 == r_count_38_io_out ? io_r_151_b : _GEN_7870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7872 = 8'h98 == r_count_38_io_out ? io_r_152_b : _GEN_7871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7873 = 8'h99 == r_count_38_io_out ? io_r_153_b : _GEN_7872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7874 = 8'h9a == r_count_38_io_out ? io_r_154_b : _GEN_7873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7875 = 8'h9b == r_count_38_io_out ? io_r_155_b : _GEN_7874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7876 = 8'h9c == r_count_38_io_out ? io_r_156_b : _GEN_7875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7877 = 8'h9d == r_count_38_io_out ? io_r_157_b : _GEN_7876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7878 = 8'h9e == r_count_38_io_out ? io_r_158_b : _GEN_7877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7879 = 8'h9f == r_count_38_io_out ? io_r_159_b : _GEN_7878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7880 = 8'ha0 == r_count_38_io_out ? io_r_160_b : _GEN_7879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7881 = 8'ha1 == r_count_38_io_out ? io_r_161_b : _GEN_7880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7882 = 8'ha2 == r_count_38_io_out ? io_r_162_b : _GEN_7881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7883 = 8'ha3 == r_count_38_io_out ? io_r_163_b : _GEN_7882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7884 = 8'ha4 == r_count_38_io_out ? io_r_164_b : _GEN_7883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7885 = 8'ha5 == r_count_38_io_out ? io_r_165_b : _GEN_7884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7886 = 8'ha6 == r_count_38_io_out ? io_r_166_b : _GEN_7885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7887 = 8'ha7 == r_count_38_io_out ? io_r_167_b : _GEN_7886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7888 = 8'ha8 == r_count_38_io_out ? io_r_168_b : _GEN_7887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7889 = 8'ha9 == r_count_38_io_out ? io_r_169_b : _GEN_7888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7890 = 8'haa == r_count_38_io_out ? io_r_170_b : _GEN_7889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7891 = 8'hab == r_count_38_io_out ? io_r_171_b : _GEN_7890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7892 = 8'hac == r_count_38_io_out ? io_r_172_b : _GEN_7891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7893 = 8'had == r_count_38_io_out ? io_r_173_b : _GEN_7892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7894 = 8'hae == r_count_38_io_out ? io_r_174_b : _GEN_7893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7895 = 8'haf == r_count_38_io_out ? io_r_175_b : _GEN_7894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7896 = 8'hb0 == r_count_38_io_out ? io_r_176_b : _GEN_7895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7897 = 8'hb1 == r_count_38_io_out ? io_r_177_b : _GEN_7896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7898 = 8'hb2 == r_count_38_io_out ? io_r_178_b : _GEN_7897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7899 = 8'hb3 == r_count_38_io_out ? io_r_179_b : _GEN_7898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7900 = 8'hb4 == r_count_38_io_out ? io_r_180_b : _GEN_7899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7901 = 8'hb5 == r_count_38_io_out ? io_r_181_b : _GEN_7900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7902 = 8'hb6 == r_count_38_io_out ? io_r_182_b : _GEN_7901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7903 = 8'hb7 == r_count_38_io_out ? io_r_183_b : _GEN_7902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7904 = 8'hb8 == r_count_38_io_out ? io_r_184_b : _GEN_7903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7905 = 8'hb9 == r_count_38_io_out ? io_r_185_b : _GEN_7904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7906 = 8'hba == r_count_38_io_out ? io_r_186_b : _GEN_7905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7907 = 8'hbb == r_count_38_io_out ? io_r_187_b : _GEN_7906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7908 = 8'hbc == r_count_38_io_out ? io_r_188_b : _GEN_7907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7909 = 8'hbd == r_count_38_io_out ? io_r_189_b : _GEN_7908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7910 = 8'hbe == r_count_38_io_out ? io_r_190_b : _GEN_7909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7911 = 8'hbf == r_count_38_io_out ? io_r_191_b : _GEN_7910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7912 = 8'hc0 == r_count_38_io_out ? io_r_192_b : _GEN_7911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7913 = 8'hc1 == r_count_38_io_out ? io_r_193_b : _GEN_7912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7914 = 8'hc2 == r_count_38_io_out ? io_r_194_b : _GEN_7913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7915 = 8'hc3 == r_count_38_io_out ? io_r_195_b : _GEN_7914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7916 = 8'hc4 == r_count_38_io_out ? io_r_196_b : _GEN_7915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7917 = 8'hc5 == r_count_38_io_out ? io_r_197_b : _GEN_7916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7918 = 8'hc6 == r_count_38_io_out ? io_r_198_b : _GEN_7917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7921 = 8'h1 == r_count_39_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7922 = 8'h2 == r_count_39_io_out ? io_r_2_b : _GEN_7921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7923 = 8'h3 == r_count_39_io_out ? io_r_3_b : _GEN_7922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7924 = 8'h4 == r_count_39_io_out ? io_r_4_b : _GEN_7923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7925 = 8'h5 == r_count_39_io_out ? io_r_5_b : _GEN_7924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7926 = 8'h6 == r_count_39_io_out ? io_r_6_b : _GEN_7925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7927 = 8'h7 == r_count_39_io_out ? io_r_7_b : _GEN_7926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7928 = 8'h8 == r_count_39_io_out ? io_r_8_b : _GEN_7927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7929 = 8'h9 == r_count_39_io_out ? io_r_9_b : _GEN_7928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7930 = 8'ha == r_count_39_io_out ? io_r_10_b : _GEN_7929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7931 = 8'hb == r_count_39_io_out ? io_r_11_b : _GEN_7930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7932 = 8'hc == r_count_39_io_out ? io_r_12_b : _GEN_7931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7933 = 8'hd == r_count_39_io_out ? io_r_13_b : _GEN_7932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7934 = 8'he == r_count_39_io_out ? io_r_14_b : _GEN_7933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7935 = 8'hf == r_count_39_io_out ? io_r_15_b : _GEN_7934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7936 = 8'h10 == r_count_39_io_out ? io_r_16_b : _GEN_7935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7937 = 8'h11 == r_count_39_io_out ? io_r_17_b : _GEN_7936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7938 = 8'h12 == r_count_39_io_out ? io_r_18_b : _GEN_7937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7939 = 8'h13 == r_count_39_io_out ? io_r_19_b : _GEN_7938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7940 = 8'h14 == r_count_39_io_out ? io_r_20_b : _GEN_7939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7941 = 8'h15 == r_count_39_io_out ? io_r_21_b : _GEN_7940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7942 = 8'h16 == r_count_39_io_out ? io_r_22_b : _GEN_7941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7943 = 8'h17 == r_count_39_io_out ? io_r_23_b : _GEN_7942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7944 = 8'h18 == r_count_39_io_out ? io_r_24_b : _GEN_7943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7945 = 8'h19 == r_count_39_io_out ? io_r_25_b : _GEN_7944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7946 = 8'h1a == r_count_39_io_out ? io_r_26_b : _GEN_7945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7947 = 8'h1b == r_count_39_io_out ? io_r_27_b : _GEN_7946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7948 = 8'h1c == r_count_39_io_out ? io_r_28_b : _GEN_7947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7949 = 8'h1d == r_count_39_io_out ? io_r_29_b : _GEN_7948; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7950 = 8'h1e == r_count_39_io_out ? io_r_30_b : _GEN_7949; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7951 = 8'h1f == r_count_39_io_out ? io_r_31_b : _GEN_7950; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7952 = 8'h20 == r_count_39_io_out ? io_r_32_b : _GEN_7951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7953 = 8'h21 == r_count_39_io_out ? io_r_33_b : _GEN_7952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7954 = 8'h22 == r_count_39_io_out ? io_r_34_b : _GEN_7953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7955 = 8'h23 == r_count_39_io_out ? io_r_35_b : _GEN_7954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7956 = 8'h24 == r_count_39_io_out ? io_r_36_b : _GEN_7955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7957 = 8'h25 == r_count_39_io_out ? io_r_37_b : _GEN_7956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7958 = 8'h26 == r_count_39_io_out ? io_r_38_b : _GEN_7957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7959 = 8'h27 == r_count_39_io_out ? io_r_39_b : _GEN_7958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7960 = 8'h28 == r_count_39_io_out ? io_r_40_b : _GEN_7959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7961 = 8'h29 == r_count_39_io_out ? io_r_41_b : _GEN_7960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7962 = 8'h2a == r_count_39_io_out ? io_r_42_b : _GEN_7961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7963 = 8'h2b == r_count_39_io_out ? io_r_43_b : _GEN_7962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7964 = 8'h2c == r_count_39_io_out ? io_r_44_b : _GEN_7963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7965 = 8'h2d == r_count_39_io_out ? io_r_45_b : _GEN_7964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7966 = 8'h2e == r_count_39_io_out ? io_r_46_b : _GEN_7965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7967 = 8'h2f == r_count_39_io_out ? io_r_47_b : _GEN_7966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7968 = 8'h30 == r_count_39_io_out ? io_r_48_b : _GEN_7967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7969 = 8'h31 == r_count_39_io_out ? io_r_49_b : _GEN_7968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7970 = 8'h32 == r_count_39_io_out ? io_r_50_b : _GEN_7969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7971 = 8'h33 == r_count_39_io_out ? io_r_51_b : _GEN_7970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7972 = 8'h34 == r_count_39_io_out ? io_r_52_b : _GEN_7971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7973 = 8'h35 == r_count_39_io_out ? io_r_53_b : _GEN_7972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7974 = 8'h36 == r_count_39_io_out ? io_r_54_b : _GEN_7973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7975 = 8'h37 == r_count_39_io_out ? io_r_55_b : _GEN_7974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7976 = 8'h38 == r_count_39_io_out ? io_r_56_b : _GEN_7975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7977 = 8'h39 == r_count_39_io_out ? io_r_57_b : _GEN_7976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7978 = 8'h3a == r_count_39_io_out ? io_r_58_b : _GEN_7977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7979 = 8'h3b == r_count_39_io_out ? io_r_59_b : _GEN_7978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7980 = 8'h3c == r_count_39_io_out ? io_r_60_b : _GEN_7979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7981 = 8'h3d == r_count_39_io_out ? io_r_61_b : _GEN_7980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7982 = 8'h3e == r_count_39_io_out ? io_r_62_b : _GEN_7981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7983 = 8'h3f == r_count_39_io_out ? io_r_63_b : _GEN_7982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7984 = 8'h40 == r_count_39_io_out ? io_r_64_b : _GEN_7983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7985 = 8'h41 == r_count_39_io_out ? io_r_65_b : _GEN_7984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7986 = 8'h42 == r_count_39_io_out ? io_r_66_b : _GEN_7985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7987 = 8'h43 == r_count_39_io_out ? io_r_67_b : _GEN_7986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7988 = 8'h44 == r_count_39_io_out ? io_r_68_b : _GEN_7987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7989 = 8'h45 == r_count_39_io_out ? io_r_69_b : _GEN_7988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7990 = 8'h46 == r_count_39_io_out ? io_r_70_b : _GEN_7989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7991 = 8'h47 == r_count_39_io_out ? io_r_71_b : _GEN_7990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7992 = 8'h48 == r_count_39_io_out ? io_r_72_b : _GEN_7991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7993 = 8'h49 == r_count_39_io_out ? io_r_73_b : _GEN_7992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7994 = 8'h4a == r_count_39_io_out ? io_r_74_b : _GEN_7993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7995 = 8'h4b == r_count_39_io_out ? io_r_75_b : _GEN_7994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7996 = 8'h4c == r_count_39_io_out ? io_r_76_b : _GEN_7995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7997 = 8'h4d == r_count_39_io_out ? io_r_77_b : _GEN_7996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7998 = 8'h4e == r_count_39_io_out ? io_r_78_b : _GEN_7997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_7999 = 8'h4f == r_count_39_io_out ? io_r_79_b : _GEN_7998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8000 = 8'h50 == r_count_39_io_out ? io_r_80_b : _GEN_7999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8001 = 8'h51 == r_count_39_io_out ? io_r_81_b : _GEN_8000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8002 = 8'h52 == r_count_39_io_out ? io_r_82_b : _GEN_8001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8003 = 8'h53 == r_count_39_io_out ? io_r_83_b : _GEN_8002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8004 = 8'h54 == r_count_39_io_out ? io_r_84_b : _GEN_8003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8005 = 8'h55 == r_count_39_io_out ? io_r_85_b : _GEN_8004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8006 = 8'h56 == r_count_39_io_out ? io_r_86_b : _GEN_8005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8007 = 8'h57 == r_count_39_io_out ? io_r_87_b : _GEN_8006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8008 = 8'h58 == r_count_39_io_out ? io_r_88_b : _GEN_8007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8009 = 8'h59 == r_count_39_io_out ? io_r_89_b : _GEN_8008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8010 = 8'h5a == r_count_39_io_out ? io_r_90_b : _GEN_8009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8011 = 8'h5b == r_count_39_io_out ? io_r_91_b : _GEN_8010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8012 = 8'h5c == r_count_39_io_out ? io_r_92_b : _GEN_8011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8013 = 8'h5d == r_count_39_io_out ? io_r_93_b : _GEN_8012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8014 = 8'h5e == r_count_39_io_out ? io_r_94_b : _GEN_8013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8015 = 8'h5f == r_count_39_io_out ? io_r_95_b : _GEN_8014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8016 = 8'h60 == r_count_39_io_out ? io_r_96_b : _GEN_8015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8017 = 8'h61 == r_count_39_io_out ? io_r_97_b : _GEN_8016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8018 = 8'h62 == r_count_39_io_out ? io_r_98_b : _GEN_8017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8019 = 8'h63 == r_count_39_io_out ? io_r_99_b : _GEN_8018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8020 = 8'h64 == r_count_39_io_out ? io_r_100_b : _GEN_8019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8021 = 8'h65 == r_count_39_io_out ? io_r_101_b : _GEN_8020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8022 = 8'h66 == r_count_39_io_out ? io_r_102_b : _GEN_8021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8023 = 8'h67 == r_count_39_io_out ? io_r_103_b : _GEN_8022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8024 = 8'h68 == r_count_39_io_out ? io_r_104_b : _GEN_8023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8025 = 8'h69 == r_count_39_io_out ? io_r_105_b : _GEN_8024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8026 = 8'h6a == r_count_39_io_out ? io_r_106_b : _GEN_8025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8027 = 8'h6b == r_count_39_io_out ? io_r_107_b : _GEN_8026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8028 = 8'h6c == r_count_39_io_out ? io_r_108_b : _GEN_8027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8029 = 8'h6d == r_count_39_io_out ? io_r_109_b : _GEN_8028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8030 = 8'h6e == r_count_39_io_out ? io_r_110_b : _GEN_8029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8031 = 8'h6f == r_count_39_io_out ? io_r_111_b : _GEN_8030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8032 = 8'h70 == r_count_39_io_out ? io_r_112_b : _GEN_8031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8033 = 8'h71 == r_count_39_io_out ? io_r_113_b : _GEN_8032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8034 = 8'h72 == r_count_39_io_out ? io_r_114_b : _GEN_8033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8035 = 8'h73 == r_count_39_io_out ? io_r_115_b : _GEN_8034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8036 = 8'h74 == r_count_39_io_out ? io_r_116_b : _GEN_8035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8037 = 8'h75 == r_count_39_io_out ? io_r_117_b : _GEN_8036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8038 = 8'h76 == r_count_39_io_out ? io_r_118_b : _GEN_8037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8039 = 8'h77 == r_count_39_io_out ? io_r_119_b : _GEN_8038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8040 = 8'h78 == r_count_39_io_out ? io_r_120_b : _GEN_8039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8041 = 8'h79 == r_count_39_io_out ? io_r_121_b : _GEN_8040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8042 = 8'h7a == r_count_39_io_out ? io_r_122_b : _GEN_8041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8043 = 8'h7b == r_count_39_io_out ? io_r_123_b : _GEN_8042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8044 = 8'h7c == r_count_39_io_out ? io_r_124_b : _GEN_8043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8045 = 8'h7d == r_count_39_io_out ? io_r_125_b : _GEN_8044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8046 = 8'h7e == r_count_39_io_out ? io_r_126_b : _GEN_8045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8047 = 8'h7f == r_count_39_io_out ? io_r_127_b : _GEN_8046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8048 = 8'h80 == r_count_39_io_out ? io_r_128_b : _GEN_8047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8049 = 8'h81 == r_count_39_io_out ? io_r_129_b : _GEN_8048; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8050 = 8'h82 == r_count_39_io_out ? io_r_130_b : _GEN_8049; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8051 = 8'h83 == r_count_39_io_out ? io_r_131_b : _GEN_8050; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8052 = 8'h84 == r_count_39_io_out ? io_r_132_b : _GEN_8051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8053 = 8'h85 == r_count_39_io_out ? io_r_133_b : _GEN_8052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8054 = 8'h86 == r_count_39_io_out ? io_r_134_b : _GEN_8053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8055 = 8'h87 == r_count_39_io_out ? io_r_135_b : _GEN_8054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8056 = 8'h88 == r_count_39_io_out ? io_r_136_b : _GEN_8055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8057 = 8'h89 == r_count_39_io_out ? io_r_137_b : _GEN_8056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8058 = 8'h8a == r_count_39_io_out ? io_r_138_b : _GEN_8057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8059 = 8'h8b == r_count_39_io_out ? io_r_139_b : _GEN_8058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8060 = 8'h8c == r_count_39_io_out ? io_r_140_b : _GEN_8059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8061 = 8'h8d == r_count_39_io_out ? io_r_141_b : _GEN_8060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8062 = 8'h8e == r_count_39_io_out ? io_r_142_b : _GEN_8061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8063 = 8'h8f == r_count_39_io_out ? io_r_143_b : _GEN_8062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8064 = 8'h90 == r_count_39_io_out ? io_r_144_b : _GEN_8063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8065 = 8'h91 == r_count_39_io_out ? io_r_145_b : _GEN_8064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8066 = 8'h92 == r_count_39_io_out ? io_r_146_b : _GEN_8065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8067 = 8'h93 == r_count_39_io_out ? io_r_147_b : _GEN_8066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8068 = 8'h94 == r_count_39_io_out ? io_r_148_b : _GEN_8067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8069 = 8'h95 == r_count_39_io_out ? io_r_149_b : _GEN_8068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8070 = 8'h96 == r_count_39_io_out ? io_r_150_b : _GEN_8069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8071 = 8'h97 == r_count_39_io_out ? io_r_151_b : _GEN_8070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8072 = 8'h98 == r_count_39_io_out ? io_r_152_b : _GEN_8071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8073 = 8'h99 == r_count_39_io_out ? io_r_153_b : _GEN_8072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8074 = 8'h9a == r_count_39_io_out ? io_r_154_b : _GEN_8073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8075 = 8'h9b == r_count_39_io_out ? io_r_155_b : _GEN_8074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8076 = 8'h9c == r_count_39_io_out ? io_r_156_b : _GEN_8075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8077 = 8'h9d == r_count_39_io_out ? io_r_157_b : _GEN_8076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8078 = 8'h9e == r_count_39_io_out ? io_r_158_b : _GEN_8077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8079 = 8'h9f == r_count_39_io_out ? io_r_159_b : _GEN_8078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8080 = 8'ha0 == r_count_39_io_out ? io_r_160_b : _GEN_8079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8081 = 8'ha1 == r_count_39_io_out ? io_r_161_b : _GEN_8080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8082 = 8'ha2 == r_count_39_io_out ? io_r_162_b : _GEN_8081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8083 = 8'ha3 == r_count_39_io_out ? io_r_163_b : _GEN_8082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8084 = 8'ha4 == r_count_39_io_out ? io_r_164_b : _GEN_8083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8085 = 8'ha5 == r_count_39_io_out ? io_r_165_b : _GEN_8084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8086 = 8'ha6 == r_count_39_io_out ? io_r_166_b : _GEN_8085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8087 = 8'ha7 == r_count_39_io_out ? io_r_167_b : _GEN_8086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8088 = 8'ha8 == r_count_39_io_out ? io_r_168_b : _GEN_8087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8089 = 8'ha9 == r_count_39_io_out ? io_r_169_b : _GEN_8088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8090 = 8'haa == r_count_39_io_out ? io_r_170_b : _GEN_8089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8091 = 8'hab == r_count_39_io_out ? io_r_171_b : _GEN_8090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8092 = 8'hac == r_count_39_io_out ? io_r_172_b : _GEN_8091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8093 = 8'had == r_count_39_io_out ? io_r_173_b : _GEN_8092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8094 = 8'hae == r_count_39_io_out ? io_r_174_b : _GEN_8093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8095 = 8'haf == r_count_39_io_out ? io_r_175_b : _GEN_8094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8096 = 8'hb0 == r_count_39_io_out ? io_r_176_b : _GEN_8095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8097 = 8'hb1 == r_count_39_io_out ? io_r_177_b : _GEN_8096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8098 = 8'hb2 == r_count_39_io_out ? io_r_178_b : _GEN_8097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8099 = 8'hb3 == r_count_39_io_out ? io_r_179_b : _GEN_8098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8100 = 8'hb4 == r_count_39_io_out ? io_r_180_b : _GEN_8099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8101 = 8'hb5 == r_count_39_io_out ? io_r_181_b : _GEN_8100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8102 = 8'hb6 == r_count_39_io_out ? io_r_182_b : _GEN_8101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8103 = 8'hb7 == r_count_39_io_out ? io_r_183_b : _GEN_8102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8104 = 8'hb8 == r_count_39_io_out ? io_r_184_b : _GEN_8103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8105 = 8'hb9 == r_count_39_io_out ? io_r_185_b : _GEN_8104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8106 = 8'hba == r_count_39_io_out ? io_r_186_b : _GEN_8105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8107 = 8'hbb == r_count_39_io_out ? io_r_187_b : _GEN_8106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8108 = 8'hbc == r_count_39_io_out ? io_r_188_b : _GEN_8107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8109 = 8'hbd == r_count_39_io_out ? io_r_189_b : _GEN_8108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8110 = 8'hbe == r_count_39_io_out ? io_r_190_b : _GEN_8109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8111 = 8'hbf == r_count_39_io_out ? io_r_191_b : _GEN_8110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8112 = 8'hc0 == r_count_39_io_out ? io_r_192_b : _GEN_8111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8113 = 8'hc1 == r_count_39_io_out ? io_r_193_b : _GEN_8112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8114 = 8'hc2 == r_count_39_io_out ? io_r_194_b : _GEN_8113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8115 = 8'hc3 == r_count_39_io_out ? io_r_195_b : _GEN_8114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8116 = 8'hc4 == r_count_39_io_out ? io_r_196_b : _GEN_8115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8117 = 8'hc5 == r_count_39_io_out ? io_r_197_b : _GEN_8116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_8118 = 8'hc6 == r_count_39_io_out ? io_r_198_b : _GEN_8117; // @[SWChisel.scala 221:{19,19}]
  SWCell array_0 ( // @[SWChisel.scala 170:39]
    .io_q(array_0_io_q),
    .io_r(array_0_io_r),
    .io_e_i(array_0_io_e_i),
    .io_f_i(array_0_io_f_i),
    .io_ve_i(array_0_io_ve_i),
    .io_vf_i(array_0_io_vf_i),
    .io_vv_i(array_0_io_vv_i),
    .io_e_o(array_0_io_e_o),
    .io_f_o(array_0_io_f_o),
    .io_v_o(array_0_io_v_o)
  );
  SWCell array_1 ( // @[SWChisel.scala 170:39]
    .io_q(array_1_io_q),
    .io_r(array_1_io_r),
    .io_e_i(array_1_io_e_i),
    .io_f_i(array_1_io_f_i),
    .io_ve_i(array_1_io_ve_i),
    .io_vf_i(array_1_io_vf_i),
    .io_vv_i(array_1_io_vv_i),
    .io_e_o(array_1_io_e_o),
    .io_f_o(array_1_io_f_o),
    .io_v_o(array_1_io_v_o)
  );
  SWCell array_2 ( // @[SWChisel.scala 170:39]
    .io_q(array_2_io_q),
    .io_r(array_2_io_r),
    .io_e_i(array_2_io_e_i),
    .io_f_i(array_2_io_f_i),
    .io_ve_i(array_2_io_ve_i),
    .io_vf_i(array_2_io_vf_i),
    .io_vv_i(array_2_io_vv_i),
    .io_e_o(array_2_io_e_o),
    .io_f_o(array_2_io_f_o),
    .io_v_o(array_2_io_v_o)
  );
  SWCell array_3 ( // @[SWChisel.scala 170:39]
    .io_q(array_3_io_q),
    .io_r(array_3_io_r),
    .io_e_i(array_3_io_e_i),
    .io_f_i(array_3_io_f_i),
    .io_ve_i(array_3_io_ve_i),
    .io_vf_i(array_3_io_vf_i),
    .io_vv_i(array_3_io_vv_i),
    .io_e_o(array_3_io_e_o),
    .io_f_o(array_3_io_f_o),
    .io_v_o(array_3_io_v_o)
  );
  SWCell array_4 ( // @[SWChisel.scala 170:39]
    .io_q(array_4_io_q),
    .io_r(array_4_io_r),
    .io_e_i(array_4_io_e_i),
    .io_f_i(array_4_io_f_i),
    .io_ve_i(array_4_io_ve_i),
    .io_vf_i(array_4_io_vf_i),
    .io_vv_i(array_4_io_vv_i),
    .io_e_o(array_4_io_e_o),
    .io_f_o(array_4_io_f_o),
    .io_v_o(array_4_io_v_o)
  );
  SWCell array_5 ( // @[SWChisel.scala 170:39]
    .io_q(array_5_io_q),
    .io_r(array_5_io_r),
    .io_e_i(array_5_io_e_i),
    .io_f_i(array_5_io_f_i),
    .io_ve_i(array_5_io_ve_i),
    .io_vf_i(array_5_io_vf_i),
    .io_vv_i(array_5_io_vv_i),
    .io_e_o(array_5_io_e_o),
    .io_f_o(array_5_io_f_o),
    .io_v_o(array_5_io_v_o)
  );
  SWCell array_6 ( // @[SWChisel.scala 170:39]
    .io_q(array_6_io_q),
    .io_r(array_6_io_r),
    .io_e_i(array_6_io_e_i),
    .io_f_i(array_6_io_f_i),
    .io_ve_i(array_6_io_ve_i),
    .io_vf_i(array_6_io_vf_i),
    .io_vv_i(array_6_io_vv_i),
    .io_e_o(array_6_io_e_o),
    .io_f_o(array_6_io_f_o),
    .io_v_o(array_6_io_v_o)
  );
  SWCell array_7 ( // @[SWChisel.scala 170:39]
    .io_q(array_7_io_q),
    .io_r(array_7_io_r),
    .io_e_i(array_7_io_e_i),
    .io_f_i(array_7_io_f_i),
    .io_ve_i(array_7_io_ve_i),
    .io_vf_i(array_7_io_vf_i),
    .io_vv_i(array_7_io_vv_i),
    .io_e_o(array_7_io_e_o),
    .io_f_o(array_7_io_f_o),
    .io_v_o(array_7_io_v_o)
  );
  SWCell array_8 ( // @[SWChisel.scala 170:39]
    .io_q(array_8_io_q),
    .io_r(array_8_io_r),
    .io_e_i(array_8_io_e_i),
    .io_f_i(array_8_io_f_i),
    .io_ve_i(array_8_io_ve_i),
    .io_vf_i(array_8_io_vf_i),
    .io_vv_i(array_8_io_vv_i),
    .io_e_o(array_8_io_e_o),
    .io_f_o(array_8_io_f_o),
    .io_v_o(array_8_io_v_o)
  );
  SWCell array_9 ( // @[SWChisel.scala 170:39]
    .io_q(array_9_io_q),
    .io_r(array_9_io_r),
    .io_e_i(array_9_io_e_i),
    .io_f_i(array_9_io_f_i),
    .io_ve_i(array_9_io_ve_i),
    .io_vf_i(array_9_io_vf_i),
    .io_vv_i(array_9_io_vv_i),
    .io_e_o(array_9_io_e_o),
    .io_f_o(array_9_io_f_o),
    .io_v_o(array_9_io_v_o)
  );
  SWCell array_10 ( // @[SWChisel.scala 170:39]
    .io_q(array_10_io_q),
    .io_r(array_10_io_r),
    .io_e_i(array_10_io_e_i),
    .io_f_i(array_10_io_f_i),
    .io_ve_i(array_10_io_ve_i),
    .io_vf_i(array_10_io_vf_i),
    .io_vv_i(array_10_io_vv_i),
    .io_e_o(array_10_io_e_o),
    .io_f_o(array_10_io_f_o),
    .io_v_o(array_10_io_v_o)
  );
  SWCell array_11 ( // @[SWChisel.scala 170:39]
    .io_q(array_11_io_q),
    .io_r(array_11_io_r),
    .io_e_i(array_11_io_e_i),
    .io_f_i(array_11_io_f_i),
    .io_ve_i(array_11_io_ve_i),
    .io_vf_i(array_11_io_vf_i),
    .io_vv_i(array_11_io_vv_i),
    .io_e_o(array_11_io_e_o),
    .io_f_o(array_11_io_f_o),
    .io_v_o(array_11_io_v_o)
  );
  SWCell array_12 ( // @[SWChisel.scala 170:39]
    .io_q(array_12_io_q),
    .io_r(array_12_io_r),
    .io_e_i(array_12_io_e_i),
    .io_f_i(array_12_io_f_i),
    .io_ve_i(array_12_io_ve_i),
    .io_vf_i(array_12_io_vf_i),
    .io_vv_i(array_12_io_vv_i),
    .io_e_o(array_12_io_e_o),
    .io_f_o(array_12_io_f_o),
    .io_v_o(array_12_io_v_o)
  );
  SWCell array_13 ( // @[SWChisel.scala 170:39]
    .io_q(array_13_io_q),
    .io_r(array_13_io_r),
    .io_e_i(array_13_io_e_i),
    .io_f_i(array_13_io_f_i),
    .io_ve_i(array_13_io_ve_i),
    .io_vf_i(array_13_io_vf_i),
    .io_vv_i(array_13_io_vv_i),
    .io_e_o(array_13_io_e_o),
    .io_f_o(array_13_io_f_o),
    .io_v_o(array_13_io_v_o)
  );
  SWCell array_14 ( // @[SWChisel.scala 170:39]
    .io_q(array_14_io_q),
    .io_r(array_14_io_r),
    .io_e_i(array_14_io_e_i),
    .io_f_i(array_14_io_f_i),
    .io_ve_i(array_14_io_ve_i),
    .io_vf_i(array_14_io_vf_i),
    .io_vv_i(array_14_io_vv_i),
    .io_e_o(array_14_io_e_o),
    .io_f_o(array_14_io_f_o),
    .io_v_o(array_14_io_v_o)
  );
  SWCell array_15 ( // @[SWChisel.scala 170:39]
    .io_q(array_15_io_q),
    .io_r(array_15_io_r),
    .io_e_i(array_15_io_e_i),
    .io_f_i(array_15_io_f_i),
    .io_ve_i(array_15_io_ve_i),
    .io_vf_i(array_15_io_vf_i),
    .io_vv_i(array_15_io_vv_i),
    .io_e_o(array_15_io_e_o),
    .io_f_o(array_15_io_f_o),
    .io_v_o(array_15_io_v_o)
  );
  SWCell array_16 ( // @[SWChisel.scala 170:39]
    .io_q(array_16_io_q),
    .io_r(array_16_io_r),
    .io_e_i(array_16_io_e_i),
    .io_f_i(array_16_io_f_i),
    .io_ve_i(array_16_io_ve_i),
    .io_vf_i(array_16_io_vf_i),
    .io_vv_i(array_16_io_vv_i),
    .io_e_o(array_16_io_e_o),
    .io_f_o(array_16_io_f_o),
    .io_v_o(array_16_io_v_o)
  );
  SWCell array_17 ( // @[SWChisel.scala 170:39]
    .io_q(array_17_io_q),
    .io_r(array_17_io_r),
    .io_e_i(array_17_io_e_i),
    .io_f_i(array_17_io_f_i),
    .io_ve_i(array_17_io_ve_i),
    .io_vf_i(array_17_io_vf_i),
    .io_vv_i(array_17_io_vv_i),
    .io_e_o(array_17_io_e_o),
    .io_f_o(array_17_io_f_o),
    .io_v_o(array_17_io_v_o)
  );
  SWCell array_18 ( // @[SWChisel.scala 170:39]
    .io_q(array_18_io_q),
    .io_r(array_18_io_r),
    .io_e_i(array_18_io_e_i),
    .io_f_i(array_18_io_f_i),
    .io_ve_i(array_18_io_ve_i),
    .io_vf_i(array_18_io_vf_i),
    .io_vv_i(array_18_io_vv_i),
    .io_e_o(array_18_io_e_o),
    .io_f_o(array_18_io_f_o),
    .io_v_o(array_18_io_v_o)
  );
  SWCell array_19 ( // @[SWChisel.scala 170:39]
    .io_q(array_19_io_q),
    .io_r(array_19_io_r),
    .io_e_i(array_19_io_e_i),
    .io_f_i(array_19_io_f_i),
    .io_ve_i(array_19_io_ve_i),
    .io_vf_i(array_19_io_vf_i),
    .io_vv_i(array_19_io_vv_i),
    .io_e_o(array_19_io_e_o),
    .io_f_o(array_19_io_f_o),
    .io_v_o(array_19_io_v_o)
  );
  SWCell array_20 ( // @[SWChisel.scala 170:39]
    .io_q(array_20_io_q),
    .io_r(array_20_io_r),
    .io_e_i(array_20_io_e_i),
    .io_f_i(array_20_io_f_i),
    .io_ve_i(array_20_io_ve_i),
    .io_vf_i(array_20_io_vf_i),
    .io_vv_i(array_20_io_vv_i),
    .io_e_o(array_20_io_e_o),
    .io_f_o(array_20_io_f_o),
    .io_v_o(array_20_io_v_o)
  );
  SWCell array_21 ( // @[SWChisel.scala 170:39]
    .io_q(array_21_io_q),
    .io_r(array_21_io_r),
    .io_e_i(array_21_io_e_i),
    .io_f_i(array_21_io_f_i),
    .io_ve_i(array_21_io_ve_i),
    .io_vf_i(array_21_io_vf_i),
    .io_vv_i(array_21_io_vv_i),
    .io_e_o(array_21_io_e_o),
    .io_f_o(array_21_io_f_o),
    .io_v_o(array_21_io_v_o)
  );
  SWCell array_22 ( // @[SWChisel.scala 170:39]
    .io_q(array_22_io_q),
    .io_r(array_22_io_r),
    .io_e_i(array_22_io_e_i),
    .io_f_i(array_22_io_f_i),
    .io_ve_i(array_22_io_ve_i),
    .io_vf_i(array_22_io_vf_i),
    .io_vv_i(array_22_io_vv_i),
    .io_e_o(array_22_io_e_o),
    .io_f_o(array_22_io_f_o),
    .io_v_o(array_22_io_v_o)
  );
  SWCell array_23 ( // @[SWChisel.scala 170:39]
    .io_q(array_23_io_q),
    .io_r(array_23_io_r),
    .io_e_i(array_23_io_e_i),
    .io_f_i(array_23_io_f_i),
    .io_ve_i(array_23_io_ve_i),
    .io_vf_i(array_23_io_vf_i),
    .io_vv_i(array_23_io_vv_i),
    .io_e_o(array_23_io_e_o),
    .io_f_o(array_23_io_f_o),
    .io_v_o(array_23_io_v_o)
  );
  SWCell array_24 ( // @[SWChisel.scala 170:39]
    .io_q(array_24_io_q),
    .io_r(array_24_io_r),
    .io_e_i(array_24_io_e_i),
    .io_f_i(array_24_io_f_i),
    .io_ve_i(array_24_io_ve_i),
    .io_vf_i(array_24_io_vf_i),
    .io_vv_i(array_24_io_vv_i),
    .io_e_o(array_24_io_e_o),
    .io_f_o(array_24_io_f_o),
    .io_v_o(array_24_io_v_o)
  );
  SWCell array_25 ( // @[SWChisel.scala 170:39]
    .io_q(array_25_io_q),
    .io_r(array_25_io_r),
    .io_e_i(array_25_io_e_i),
    .io_f_i(array_25_io_f_i),
    .io_ve_i(array_25_io_ve_i),
    .io_vf_i(array_25_io_vf_i),
    .io_vv_i(array_25_io_vv_i),
    .io_e_o(array_25_io_e_o),
    .io_f_o(array_25_io_f_o),
    .io_v_o(array_25_io_v_o)
  );
  SWCell array_26 ( // @[SWChisel.scala 170:39]
    .io_q(array_26_io_q),
    .io_r(array_26_io_r),
    .io_e_i(array_26_io_e_i),
    .io_f_i(array_26_io_f_i),
    .io_ve_i(array_26_io_ve_i),
    .io_vf_i(array_26_io_vf_i),
    .io_vv_i(array_26_io_vv_i),
    .io_e_o(array_26_io_e_o),
    .io_f_o(array_26_io_f_o),
    .io_v_o(array_26_io_v_o)
  );
  SWCell array_27 ( // @[SWChisel.scala 170:39]
    .io_q(array_27_io_q),
    .io_r(array_27_io_r),
    .io_e_i(array_27_io_e_i),
    .io_f_i(array_27_io_f_i),
    .io_ve_i(array_27_io_ve_i),
    .io_vf_i(array_27_io_vf_i),
    .io_vv_i(array_27_io_vv_i),
    .io_e_o(array_27_io_e_o),
    .io_f_o(array_27_io_f_o),
    .io_v_o(array_27_io_v_o)
  );
  SWCell array_28 ( // @[SWChisel.scala 170:39]
    .io_q(array_28_io_q),
    .io_r(array_28_io_r),
    .io_e_i(array_28_io_e_i),
    .io_f_i(array_28_io_f_i),
    .io_ve_i(array_28_io_ve_i),
    .io_vf_i(array_28_io_vf_i),
    .io_vv_i(array_28_io_vv_i),
    .io_e_o(array_28_io_e_o),
    .io_f_o(array_28_io_f_o),
    .io_v_o(array_28_io_v_o)
  );
  SWCell array_29 ( // @[SWChisel.scala 170:39]
    .io_q(array_29_io_q),
    .io_r(array_29_io_r),
    .io_e_i(array_29_io_e_i),
    .io_f_i(array_29_io_f_i),
    .io_ve_i(array_29_io_ve_i),
    .io_vf_i(array_29_io_vf_i),
    .io_vv_i(array_29_io_vv_i),
    .io_e_o(array_29_io_e_o),
    .io_f_o(array_29_io_f_o),
    .io_v_o(array_29_io_v_o)
  );
  SWCell array_30 ( // @[SWChisel.scala 170:39]
    .io_q(array_30_io_q),
    .io_r(array_30_io_r),
    .io_e_i(array_30_io_e_i),
    .io_f_i(array_30_io_f_i),
    .io_ve_i(array_30_io_ve_i),
    .io_vf_i(array_30_io_vf_i),
    .io_vv_i(array_30_io_vv_i),
    .io_e_o(array_30_io_e_o),
    .io_f_o(array_30_io_f_o),
    .io_v_o(array_30_io_v_o)
  );
  SWCell array_31 ( // @[SWChisel.scala 170:39]
    .io_q(array_31_io_q),
    .io_r(array_31_io_r),
    .io_e_i(array_31_io_e_i),
    .io_f_i(array_31_io_f_i),
    .io_ve_i(array_31_io_ve_i),
    .io_vf_i(array_31_io_vf_i),
    .io_vv_i(array_31_io_vv_i),
    .io_e_o(array_31_io_e_o),
    .io_f_o(array_31_io_f_o),
    .io_v_o(array_31_io_v_o)
  );
  SWCell array_32 ( // @[SWChisel.scala 170:39]
    .io_q(array_32_io_q),
    .io_r(array_32_io_r),
    .io_e_i(array_32_io_e_i),
    .io_f_i(array_32_io_f_i),
    .io_ve_i(array_32_io_ve_i),
    .io_vf_i(array_32_io_vf_i),
    .io_vv_i(array_32_io_vv_i),
    .io_e_o(array_32_io_e_o),
    .io_f_o(array_32_io_f_o),
    .io_v_o(array_32_io_v_o)
  );
  SWCell array_33 ( // @[SWChisel.scala 170:39]
    .io_q(array_33_io_q),
    .io_r(array_33_io_r),
    .io_e_i(array_33_io_e_i),
    .io_f_i(array_33_io_f_i),
    .io_ve_i(array_33_io_ve_i),
    .io_vf_i(array_33_io_vf_i),
    .io_vv_i(array_33_io_vv_i),
    .io_e_o(array_33_io_e_o),
    .io_f_o(array_33_io_f_o),
    .io_v_o(array_33_io_v_o)
  );
  SWCell array_34 ( // @[SWChisel.scala 170:39]
    .io_q(array_34_io_q),
    .io_r(array_34_io_r),
    .io_e_i(array_34_io_e_i),
    .io_f_i(array_34_io_f_i),
    .io_ve_i(array_34_io_ve_i),
    .io_vf_i(array_34_io_vf_i),
    .io_vv_i(array_34_io_vv_i),
    .io_e_o(array_34_io_e_o),
    .io_f_o(array_34_io_f_o),
    .io_v_o(array_34_io_v_o)
  );
  SWCell array_35 ( // @[SWChisel.scala 170:39]
    .io_q(array_35_io_q),
    .io_r(array_35_io_r),
    .io_e_i(array_35_io_e_i),
    .io_f_i(array_35_io_f_i),
    .io_ve_i(array_35_io_ve_i),
    .io_vf_i(array_35_io_vf_i),
    .io_vv_i(array_35_io_vv_i),
    .io_e_o(array_35_io_e_o),
    .io_f_o(array_35_io_f_o),
    .io_v_o(array_35_io_v_o)
  );
  SWCell array_36 ( // @[SWChisel.scala 170:39]
    .io_q(array_36_io_q),
    .io_r(array_36_io_r),
    .io_e_i(array_36_io_e_i),
    .io_f_i(array_36_io_f_i),
    .io_ve_i(array_36_io_ve_i),
    .io_vf_i(array_36_io_vf_i),
    .io_vv_i(array_36_io_vv_i),
    .io_e_o(array_36_io_e_o),
    .io_f_o(array_36_io_f_o),
    .io_v_o(array_36_io_v_o)
  );
  SWCell array_37 ( // @[SWChisel.scala 170:39]
    .io_q(array_37_io_q),
    .io_r(array_37_io_r),
    .io_e_i(array_37_io_e_i),
    .io_f_i(array_37_io_f_i),
    .io_ve_i(array_37_io_ve_i),
    .io_vf_i(array_37_io_vf_i),
    .io_vv_i(array_37_io_vv_i),
    .io_e_o(array_37_io_e_o),
    .io_f_o(array_37_io_f_o),
    .io_v_o(array_37_io_v_o)
  );
  SWCell array_38 ( // @[SWChisel.scala 170:39]
    .io_q(array_38_io_q),
    .io_r(array_38_io_r),
    .io_e_i(array_38_io_e_i),
    .io_f_i(array_38_io_f_i),
    .io_ve_i(array_38_io_ve_i),
    .io_vf_i(array_38_io_vf_i),
    .io_vv_i(array_38_io_vv_i),
    .io_e_o(array_38_io_e_o),
    .io_f_o(array_38_io_f_o),
    .io_v_o(array_38_io_v_o)
  );
  SWCell array_39 ( // @[SWChisel.scala 170:39]
    .io_q(array_39_io_q),
    .io_r(array_39_io_r),
    .io_e_i(array_39_io_e_i),
    .io_f_i(array_39_io_f_i),
    .io_ve_i(array_39_io_ve_i),
    .io_vf_i(array_39_io_vf_i),
    .io_vv_i(array_39_io_vv_i),
    .io_e_o(array_39_io_e_o),
    .io_f_o(array_39_io_f_o),
    .io_v_o(array_39_io_v_o)
  );
  MyCounter r_count_0 ( // @[SWChisel.scala 171:41]
    .clock(r_count_0_clock),
    .reset(r_count_0_reset),
    .io_en(r_count_0_io_en),
    .io_out(r_count_0_io_out)
  );
  MyCounter r_count_1 ( // @[SWChisel.scala 171:41]
    .clock(r_count_1_clock),
    .reset(r_count_1_reset),
    .io_en(r_count_1_io_en),
    .io_out(r_count_1_io_out)
  );
  MyCounter r_count_2 ( // @[SWChisel.scala 171:41]
    .clock(r_count_2_clock),
    .reset(r_count_2_reset),
    .io_en(r_count_2_io_en),
    .io_out(r_count_2_io_out)
  );
  MyCounter r_count_3 ( // @[SWChisel.scala 171:41]
    .clock(r_count_3_clock),
    .reset(r_count_3_reset),
    .io_en(r_count_3_io_en),
    .io_out(r_count_3_io_out)
  );
  MyCounter r_count_4 ( // @[SWChisel.scala 171:41]
    .clock(r_count_4_clock),
    .reset(r_count_4_reset),
    .io_en(r_count_4_io_en),
    .io_out(r_count_4_io_out)
  );
  MyCounter r_count_5 ( // @[SWChisel.scala 171:41]
    .clock(r_count_5_clock),
    .reset(r_count_5_reset),
    .io_en(r_count_5_io_en),
    .io_out(r_count_5_io_out)
  );
  MyCounter r_count_6 ( // @[SWChisel.scala 171:41]
    .clock(r_count_6_clock),
    .reset(r_count_6_reset),
    .io_en(r_count_6_io_en),
    .io_out(r_count_6_io_out)
  );
  MyCounter r_count_7 ( // @[SWChisel.scala 171:41]
    .clock(r_count_7_clock),
    .reset(r_count_7_reset),
    .io_en(r_count_7_io_en),
    .io_out(r_count_7_io_out)
  );
  MyCounter r_count_8 ( // @[SWChisel.scala 171:41]
    .clock(r_count_8_clock),
    .reset(r_count_8_reset),
    .io_en(r_count_8_io_en),
    .io_out(r_count_8_io_out)
  );
  MyCounter r_count_9 ( // @[SWChisel.scala 171:41]
    .clock(r_count_9_clock),
    .reset(r_count_9_reset),
    .io_en(r_count_9_io_en),
    .io_out(r_count_9_io_out)
  );
  MyCounter r_count_10 ( // @[SWChisel.scala 171:41]
    .clock(r_count_10_clock),
    .reset(r_count_10_reset),
    .io_en(r_count_10_io_en),
    .io_out(r_count_10_io_out)
  );
  MyCounter r_count_11 ( // @[SWChisel.scala 171:41]
    .clock(r_count_11_clock),
    .reset(r_count_11_reset),
    .io_en(r_count_11_io_en),
    .io_out(r_count_11_io_out)
  );
  MyCounter r_count_12 ( // @[SWChisel.scala 171:41]
    .clock(r_count_12_clock),
    .reset(r_count_12_reset),
    .io_en(r_count_12_io_en),
    .io_out(r_count_12_io_out)
  );
  MyCounter r_count_13 ( // @[SWChisel.scala 171:41]
    .clock(r_count_13_clock),
    .reset(r_count_13_reset),
    .io_en(r_count_13_io_en),
    .io_out(r_count_13_io_out)
  );
  MyCounter r_count_14 ( // @[SWChisel.scala 171:41]
    .clock(r_count_14_clock),
    .reset(r_count_14_reset),
    .io_en(r_count_14_io_en),
    .io_out(r_count_14_io_out)
  );
  MyCounter r_count_15 ( // @[SWChisel.scala 171:41]
    .clock(r_count_15_clock),
    .reset(r_count_15_reset),
    .io_en(r_count_15_io_en),
    .io_out(r_count_15_io_out)
  );
  MyCounter r_count_16 ( // @[SWChisel.scala 171:41]
    .clock(r_count_16_clock),
    .reset(r_count_16_reset),
    .io_en(r_count_16_io_en),
    .io_out(r_count_16_io_out)
  );
  MyCounter r_count_17 ( // @[SWChisel.scala 171:41]
    .clock(r_count_17_clock),
    .reset(r_count_17_reset),
    .io_en(r_count_17_io_en),
    .io_out(r_count_17_io_out)
  );
  MyCounter r_count_18 ( // @[SWChisel.scala 171:41]
    .clock(r_count_18_clock),
    .reset(r_count_18_reset),
    .io_en(r_count_18_io_en),
    .io_out(r_count_18_io_out)
  );
  MyCounter r_count_19 ( // @[SWChisel.scala 171:41]
    .clock(r_count_19_clock),
    .reset(r_count_19_reset),
    .io_en(r_count_19_io_en),
    .io_out(r_count_19_io_out)
  );
  MyCounter r_count_20 ( // @[SWChisel.scala 171:41]
    .clock(r_count_20_clock),
    .reset(r_count_20_reset),
    .io_en(r_count_20_io_en),
    .io_out(r_count_20_io_out)
  );
  MyCounter r_count_21 ( // @[SWChisel.scala 171:41]
    .clock(r_count_21_clock),
    .reset(r_count_21_reset),
    .io_en(r_count_21_io_en),
    .io_out(r_count_21_io_out)
  );
  MyCounter r_count_22 ( // @[SWChisel.scala 171:41]
    .clock(r_count_22_clock),
    .reset(r_count_22_reset),
    .io_en(r_count_22_io_en),
    .io_out(r_count_22_io_out)
  );
  MyCounter r_count_23 ( // @[SWChisel.scala 171:41]
    .clock(r_count_23_clock),
    .reset(r_count_23_reset),
    .io_en(r_count_23_io_en),
    .io_out(r_count_23_io_out)
  );
  MyCounter r_count_24 ( // @[SWChisel.scala 171:41]
    .clock(r_count_24_clock),
    .reset(r_count_24_reset),
    .io_en(r_count_24_io_en),
    .io_out(r_count_24_io_out)
  );
  MyCounter r_count_25 ( // @[SWChisel.scala 171:41]
    .clock(r_count_25_clock),
    .reset(r_count_25_reset),
    .io_en(r_count_25_io_en),
    .io_out(r_count_25_io_out)
  );
  MyCounter r_count_26 ( // @[SWChisel.scala 171:41]
    .clock(r_count_26_clock),
    .reset(r_count_26_reset),
    .io_en(r_count_26_io_en),
    .io_out(r_count_26_io_out)
  );
  MyCounter r_count_27 ( // @[SWChisel.scala 171:41]
    .clock(r_count_27_clock),
    .reset(r_count_27_reset),
    .io_en(r_count_27_io_en),
    .io_out(r_count_27_io_out)
  );
  MyCounter r_count_28 ( // @[SWChisel.scala 171:41]
    .clock(r_count_28_clock),
    .reset(r_count_28_reset),
    .io_en(r_count_28_io_en),
    .io_out(r_count_28_io_out)
  );
  MyCounter r_count_29 ( // @[SWChisel.scala 171:41]
    .clock(r_count_29_clock),
    .reset(r_count_29_reset),
    .io_en(r_count_29_io_en),
    .io_out(r_count_29_io_out)
  );
  MyCounter r_count_30 ( // @[SWChisel.scala 171:41]
    .clock(r_count_30_clock),
    .reset(r_count_30_reset),
    .io_en(r_count_30_io_en),
    .io_out(r_count_30_io_out)
  );
  MyCounter r_count_31 ( // @[SWChisel.scala 171:41]
    .clock(r_count_31_clock),
    .reset(r_count_31_reset),
    .io_en(r_count_31_io_en),
    .io_out(r_count_31_io_out)
  );
  MyCounter r_count_32 ( // @[SWChisel.scala 171:41]
    .clock(r_count_32_clock),
    .reset(r_count_32_reset),
    .io_en(r_count_32_io_en),
    .io_out(r_count_32_io_out)
  );
  MyCounter r_count_33 ( // @[SWChisel.scala 171:41]
    .clock(r_count_33_clock),
    .reset(r_count_33_reset),
    .io_en(r_count_33_io_en),
    .io_out(r_count_33_io_out)
  );
  MyCounter r_count_34 ( // @[SWChisel.scala 171:41]
    .clock(r_count_34_clock),
    .reset(r_count_34_reset),
    .io_en(r_count_34_io_en),
    .io_out(r_count_34_io_out)
  );
  MyCounter r_count_35 ( // @[SWChisel.scala 171:41]
    .clock(r_count_35_clock),
    .reset(r_count_35_reset),
    .io_en(r_count_35_io_en),
    .io_out(r_count_35_io_out)
  );
  MyCounter r_count_36 ( // @[SWChisel.scala 171:41]
    .clock(r_count_36_clock),
    .reset(r_count_36_reset),
    .io_en(r_count_36_io_en),
    .io_out(r_count_36_io_out)
  );
  MyCounter r_count_37 ( // @[SWChisel.scala 171:41]
    .clock(r_count_37_clock),
    .reset(r_count_37_reset),
    .io_en(r_count_37_io_en),
    .io_out(r_count_37_io_out)
  );
  MyCounter r_count_38 ( // @[SWChisel.scala 171:41]
    .clock(r_count_38_clock),
    .reset(r_count_38_reset),
    .io_en(r_count_38_io_en),
    .io_out(r_count_38_io_out)
  );
  MyCounter r_count_39 ( // @[SWChisel.scala 171:41]
    .clock(r_count_39_clock),
    .reset(r_count_39_reset),
    .io_en(r_count_39_io_en),
    .io_out(r_count_39_io_out)
  );
  MAX max ( // @[SWChisel.scala 174:19]
    .clock(max_clock),
    .reset(max_reset),
    .io_start(max_io_start),
    .io_in(max_io_in),
    .io_done(max_io_done),
    .io_out(max_io_out)
  );
  assign io_result = max_io_out; // @[SWChisel.scala 181:13]
  assign io_done = max_io_done; // @[SWChisel.scala 182:11]
  assign array_0_io_q = io_q_0_b; // @[SWChisel.scala 220:19]
  assign array_0_io_r = 8'hc7 == r_count_0_io_out ? io_r_199_b : _GEN_318; // @[SWChisel.scala 221:{19,19}]
  assign array_0_io_e_i = E_0; // @[SWChisel.scala 196:21]
  assign array_0_io_f_i = 16'sh0; // @[SWChisel.scala 198:21]
  assign array_0_io_ve_i = V1_1; // @[SWChisel.scala 197:22]
  assign array_0_io_vf_i = V1_0; // @[SWChisel.scala 199:22]
  assign array_0_io_vv_i = V2_0; // @[SWChisel.scala 200:22]
  assign array_1_io_q = io_q_1_b; // @[SWChisel.scala 220:19]
  assign array_1_io_r = 8'hc7 == r_count_1_io_out ? io_r_199_b : _GEN_518; // @[SWChisel.scala 221:{19,19}]
  assign array_1_io_e_i = E_1; // @[SWChisel.scala 196:21]
  assign array_1_io_f_i = F_1; // @[SWChisel.scala 198:21]
  assign array_1_io_ve_i = V1_2; // @[SWChisel.scala 197:22]
  assign array_1_io_vf_i = V1_1; // @[SWChisel.scala 199:22]
  assign array_1_io_vv_i = V2_1; // @[SWChisel.scala 200:22]
  assign array_2_io_q = io_q_2_b; // @[SWChisel.scala 220:19]
  assign array_2_io_r = 8'hc7 == r_count_2_io_out ? io_r_199_b : _GEN_718; // @[SWChisel.scala 221:{19,19}]
  assign array_2_io_e_i = E_2; // @[SWChisel.scala 196:21]
  assign array_2_io_f_i = F_2; // @[SWChisel.scala 198:21]
  assign array_2_io_ve_i = V1_3; // @[SWChisel.scala 197:22]
  assign array_2_io_vf_i = V1_2; // @[SWChisel.scala 199:22]
  assign array_2_io_vv_i = V2_2; // @[SWChisel.scala 200:22]
  assign array_3_io_q = io_q_3_b; // @[SWChisel.scala 220:19]
  assign array_3_io_r = 8'hc7 == r_count_3_io_out ? io_r_199_b : _GEN_918; // @[SWChisel.scala 221:{19,19}]
  assign array_3_io_e_i = E_3; // @[SWChisel.scala 196:21]
  assign array_3_io_f_i = F_3; // @[SWChisel.scala 198:21]
  assign array_3_io_ve_i = V1_4; // @[SWChisel.scala 197:22]
  assign array_3_io_vf_i = V1_3; // @[SWChisel.scala 199:22]
  assign array_3_io_vv_i = V2_3; // @[SWChisel.scala 200:22]
  assign array_4_io_q = io_q_4_b; // @[SWChisel.scala 220:19]
  assign array_4_io_r = 8'hc7 == r_count_4_io_out ? io_r_199_b : _GEN_1118; // @[SWChisel.scala 221:{19,19}]
  assign array_4_io_e_i = E_4; // @[SWChisel.scala 196:21]
  assign array_4_io_f_i = F_4; // @[SWChisel.scala 198:21]
  assign array_4_io_ve_i = V1_5; // @[SWChisel.scala 197:22]
  assign array_4_io_vf_i = V1_4; // @[SWChisel.scala 199:22]
  assign array_4_io_vv_i = V2_4; // @[SWChisel.scala 200:22]
  assign array_5_io_q = io_q_5_b; // @[SWChisel.scala 220:19]
  assign array_5_io_r = 8'hc7 == r_count_5_io_out ? io_r_199_b : _GEN_1318; // @[SWChisel.scala 221:{19,19}]
  assign array_5_io_e_i = E_5; // @[SWChisel.scala 196:21]
  assign array_5_io_f_i = F_5; // @[SWChisel.scala 198:21]
  assign array_5_io_ve_i = V1_6; // @[SWChisel.scala 197:22]
  assign array_5_io_vf_i = V1_5; // @[SWChisel.scala 199:22]
  assign array_5_io_vv_i = V2_5; // @[SWChisel.scala 200:22]
  assign array_6_io_q = io_q_6_b; // @[SWChisel.scala 220:19]
  assign array_6_io_r = 8'hc7 == r_count_6_io_out ? io_r_199_b : _GEN_1518; // @[SWChisel.scala 221:{19,19}]
  assign array_6_io_e_i = E_6; // @[SWChisel.scala 196:21]
  assign array_6_io_f_i = F_6; // @[SWChisel.scala 198:21]
  assign array_6_io_ve_i = V1_7; // @[SWChisel.scala 197:22]
  assign array_6_io_vf_i = V1_6; // @[SWChisel.scala 199:22]
  assign array_6_io_vv_i = V2_6; // @[SWChisel.scala 200:22]
  assign array_7_io_q = io_q_7_b; // @[SWChisel.scala 220:19]
  assign array_7_io_r = 8'hc7 == r_count_7_io_out ? io_r_199_b : _GEN_1718; // @[SWChisel.scala 221:{19,19}]
  assign array_7_io_e_i = E_7; // @[SWChisel.scala 196:21]
  assign array_7_io_f_i = F_7; // @[SWChisel.scala 198:21]
  assign array_7_io_ve_i = V1_8; // @[SWChisel.scala 197:22]
  assign array_7_io_vf_i = V1_7; // @[SWChisel.scala 199:22]
  assign array_7_io_vv_i = V2_7; // @[SWChisel.scala 200:22]
  assign array_8_io_q = io_q_8_b; // @[SWChisel.scala 220:19]
  assign array_8_io_r = 8'hc7 == r_count_8_io_out ? io_r_199_b : _GEN_1918; // @[SWChisel.scala 221:{19,19}]
  assign array_8_io_e_i = E_8; // @[SWChisel.scala 196:21]
  assign array_8_io_f_i = F_8; // @[SWChisel.scala 198:21]
  assign array_8_io_ve_i = V1_9; // @[SWChisel.scala 197:22]
  assign array_8_io_vf_i = V1_8; // @[SWChisel.scala 199:22]
  assign array_8_io_vv_i = V2_8; // @[SWChisel.scala 200:22]
  assign array_9_io_q = io_q_9_b; // @[SWChisel.scala 220:19]
  assign array_9_io_r = 8'hc7 == r_count_9_io_out ? io_r_199_b : _GEN_2118; // @[SWChisel.scala 221:{19,19}]
  assign array_9_io_e_i = E_9; // @[SWChisel.scala 196:21]
  assign array_9_io_f_i = F_9; // @[SWChisel.scala 198:21]
  assign array_9_io_ve_i = V1_10; // @[SWChisel.scala 197:22]
  assign array_9_io_vf_i = V1_9; // @[SWChisel.scala 199:22]
  assign array_9_io_vv_i = V2_9; // @[SWChisel.scala 200:22]
  assign array_10_io_q = io_q_10_b; // @[SWChisel.scala 220:19]
  assign array_10_io_r = 8'hc7 == r_count_10_io_out ? io_r_199_b : _GEN_2318; // @[SWChisel.scala 221:{19,19}]
  assign array_10_io_e_i = E_10; // @[SWChisel.scala 196:21]
  assign array_10_io_f_i = F_10; // @[SWChisel.scala 198:21]
  assign array_10_io_ve_i = V1_11; // @[SWChisel.scala 197:22]
  assign array_10_io_vf_i = V1_10; // @[SWChisel.scala 199:22]
  assign array_10_io_vv_i = V2_10; // @[SWChisel.scala 200:22]
  assign array_11_io_q = io_q_11_b; // @[SWChisel.scala 220:19]
  assign array_11_io_r = 8'hc7 == r_count_11_io_out ? io_r_199_b : _GEN_2518; // @[SWChisel.scala 221:{19,19}]
  assign array_11_io_e_i = E_11; // @[SWChisel.scala 196:21]
  assign array_11_io_f_i = F_11; // @[SWChisel.scala 198:21]
  assign array_11_io_ve_i = V1_12; // @[SWChisel.scala 197:22]
  assign array_11_io_vf_i = V1_11; // @[SWChisel.scala 199:22]
  assign array_11_io_vv_i = V2_11; // @[SWChisel.scala 200:22]
  assign array_12_io_q = io_q_12_b; // @[SWChisel.scala 220:19]
  assign array_12_io_r = 8'hc7 == r_count_12_io_out ? io_r_199_b : _GEN_2718; // @[SWChisel.scala 221:{19,19}]
  assign array_12_io_e_i = E_12; // @[SWChisel.scala 196:21]
  assign array_12_io_f_i = F_12; // @[SWChisel.scala 198:21]
  assign array_12_io_ve_i = V1_13; // @[SWChisel.scala 197:22]
  assign array_12_io_vf_i = V1_12; // @[SWChisel.scala 199:22]
  assign array_12_io_vv_i = V2_12; // @[SWChisel.scala 200:22]
  assign array_13_io_q = io_q_13_b; // @[SWChisel.scala 220:19]
  assign array_13_io_r = 8'hc7 == r_count_13_io_out ? io_r_199_b : _GEN_2918; // @[SWChisel.scala 221:{19,19}]
  assign array_13_io_e_i = E_13; // @[SWChisel.scala 196:21]
  assign array_13_io_f_i = F_13; // @[SWChisel.scala 198:21]
  assign array_13_io_ve_i = V1_14; // @[SWChisel.scala 197:22]
  assign array_13_io_vf_i = V1_13; // @[SWChisel.scala 199:22]
  assign array_13_io_vv_i = V2_13; // @[SWChisel.scala 200:22]
  assign array_14_io_q = io_q_14_b; // @[SWChisel.scala 220:19]
  assign array_14_io_r = 8'hc7 == r_count_14_io_out ? io_r_199_b : _GEN_3118; // @[SWChisel.scala 221:{19,19}]
  assign array_14_io_e_i = E_14; // @[SWChisel.scala 196:21]
  assign array_14_io_f_i = F_14; // @[SWChisel.scala 198:21]
  assign array_14_io_ve_i = V1_15; // @[SWChisel.scala 197:22]
  assign array_14_io_vf_i = V1_14; // @[SWChisel.scala 199:22]
  assign array_14_io_vv_i = V2_14; // @[SWChisel.scala 200:22]
  assign array_15_io_q = io_q_15_b; // @[SWChisel.scala 220:19]
  assign array_15_io_r = 8'hc7 == r_count_15_io_out ? io_r_199_b : _GEN_3318; // @[SWChisel.scala 221:{19,19}]
  assign array_15_io_e_i = E_15; // @[SWChisel.scala 196:21]
  assign array_15_io_f_i = F_15; // @[SWChisel.scala 198:21]
  assign array_15_io_ve_i = V1_16; // @[SWChisel.scala 197:22]
  assign array_15_io_vf_i = V1_15; // @[SWChisel.scala 199:22]
  assign array_15_io_vv_i = V2_15; // @[SWChisel.scala 200:22]
  assign array_16_io_q = io_q_16_b; // @[SWChisel.scala 220:19]
  assign array_16_io_r = 8'hc7 == r_count_16_io_out ? io_r_199_b : _GEN_3518; // @[SWChisel.scala 221:{19,19}]
  assign array_16_io_e_i = E_16; // @[SWChisel.scala 196:21]
  assign array_16_io_f_i = F_16; // @[SWChisel.scala 198:21]
  assign array_16_io_ve_i = V1_17; // @[SWChisel.scala 197:22]
  assign array_16_io_vf_i = V1_16; // @[SWChisel.scala 199:22]
  assign array_16_io_vv_i = V2_16; // @[SWChisel.scala 200:22]
  assign array_17_io_q = io_q_17_b; // @[SWChisel.scala 220:19]
  assign array_17_io_r = 8'hc7 == r_count_17_io_out ? io_r_199_b : _GEN_3718; // @[SWChisel.scala 221:{19,19}]
  assign array_17_io_e_i = E_17; // @[SWChisel.scala 196:21]
  assign array_17_io_f_i = F_17; // @[SWChisel.scala 198:21]
  assign array_17_io_ve_i = V1_18; // @[SWChisel.scala 197:22]
  assign array_17_io_vf_i = V1_17; // @[SWChisel.scala 199:22]
  assign array_17_io_vv_i = V2_17; // @[SWChisel.scala 200:22]
  assign array_18_io_q = io_q_18_b; // @[SWChisel.scala 220:19]
  assign array_18_io_r = 8'hc7 == r_count_18_io_out ? io_r_199_b : _GEN_3918; // @[SWChisel.scala 221:{19,19}]
  assign array_18_io_e_i = E_18; // @[SWChisel.scala 196:21]
  assign array_18_io_f_i = F_18; // @[SWChisel.scala 198:21]
  assign array_18_io_ve_i = V1_19; // @[SWChisel.scala 197:22]
  assign array_18_io_vf_i = V1_18; // @[SWChisel.scala 199:22]
  assign array_18_io_vv_i = V2_18; // @[SWChisel.scala 200:22]
  assign array_19_io_q = io_q_19_b; // @[SWChisel.scala 220:19]
  assign array_19_io_r = 8'hc7 == r_count_19_io_out ? io_r_199_b : _GEN_4118; // @[SWChisel.scala 221:{19,19}]
  assign array_19_io_e_i = E_19; // @[SWChisel.scala 196:21]
  assign array_19_io_f_i = F_19; // @[SWChisel.scala 198:21]
  assign array_19_io_ve_i = V1_20; // @[SWChisel.scala 197:22]
  assign array_19_io_vf_i = V1_19; // @[SWChisel.scala 199:22]
  assign array_19_io_vv_i = V2_19; // @[SWChisel.scala 200:22]
  assign array_20_io_q = io_q_20_b; // @[SWChisel.scala 220:19]
  assign array_20_io_r = 8'hc7 == r_count_20_io_out ? io_r_199_b : _GEN_4318; // @[SWChisel.scala 221:{19,19}]
  assign array_20_io_e_i = E_20; // @[SWChisel.scala 196:21]
  assign array_20_io_f_i = F_20; // @[SWChisel.scala 198:21]
  assign array_20_io_ve_i = V1_21; // @[SWChisel.scala 197:22]
  assign array_20_io_vf_i = V1_20; // @[SWChisel.scala 199:22]
  assign array_20_io_vv_i = V2_20; // @[SWChisel.scala 200:22]
  assign array_21_io_q = io_q_21_b; // @[SWChisel.scala 220:19]
  assign array_21_io_r = 8'hc7 == r_count_21_io_out ? io_r_199_b : _GEN_4518; // @[SWChisel.scala 221:{19,19}]
  assign array_21_io_e_i = E_21; // @[SWChisel.scala 196:21]
  assign array_21_io_f_i = F_21; // @[SWChisel.scala 198:21]
  assign array_21_io_ve_i = V1_22; // @[SWChisel.scala 197:22]
  assign array_21_io_vf_i = V1_21; // @[SWChisel.scala 199:22]
  assign array_21_io_vv_i = V2_21; // @[SWChisel.scala 200:22]
  assign array_22_io_q = io_q_22_b; // @[SWChisel.scala 220:19]
  assign array_22_io_r = 8'hc7 == r_count_22_io_out ? io_r_199_b : _GEN_4718; // @[SWChisel.scala 221:{19,19}]
  assign array_22_io_e_i = E_22; // @[SWChisel.scala 196:21]
  assign array_22_io_f_i = F_22; // @[SWChisel.scala 198:21]
  assign array_22_io_ve_i = V1_23; // @[SWChisel.scala 197:22]
  assign array_22_io_vf_i = V1_22; // @[SWChisel.scala 199:22]
  assign array_22_io_vv_i = V2_22; // @[SWChisel.scala 200:22]
  assign array_23_io_q = io_q_23_b; // @[SWChisel.scala 220:19]
  assign array_23_io_r = 8'hc7 == r_count_23_io_out ? io_r_199_b : _GEN_4918; // @[SWChisel.scala 221:{19,19}]
  assign array_23_io_e_i = E_23; // @[SWChisel.scala 196:21]
  assign array_23_io_f_i = F_23; // @[SWChisel.scala 198:21]
  assign array_23_io_ve_i = V1_24; // @[SWChisel.scala 197:22]
  assign array_23_io_vf_i = V1_23; // @[SWChisel.scala 199:22]
  assign array_23_io_vv_i = V2_23; // @[SWChisel.scala 200:22]
  assign array_24_io_q = io_q_24_b; // @[SWChisel.scala 220:19]
  assign array_24_io_r = 8'hc7 == r_count_24_io_out ? io_r_199_b : _GEN_5118; // @[SWChisel.scala 221:{19,19}]
  assign array_24_io_e_i = E_24; // @[SWChisel.scala 196:21]
  assign array_24_io_f_i = F_24; // @[SWChisel.scala 198:21]
  assign array_24_io_ve_i = V1_25; // @[SWChisel.scala 197:22]
  assign array_24_io_vf_i = V1_24; // @[SWChisel.scala 199:22]
  assign array_24_io_vv_i = V2_24; // @[SWChisel.scala 200:22]
  assign array_25_io_q = io_q_25_b; // @[SWChisel.scala 220:19]
  assign array_25_io_r = 8'hc7 == r_count_25_io_out ? io_r_199_b : _GEN_5318; // @[SWChisel.scala 221:{19,19}]
  assign array_25_io_e_i = E_25; // @[SWChisel.scala 196:21]
  assign array_25_io_f_i = F_25; // @[SWChisel.scala 198:21]
  assign array_25_io_ve_i = V1_26; // @[SWChisel.scala 197:22]
  assign array_25_io_vf_i = V1_25; // @[SWChisel.scala 199:22]
  assign array_25_io_vv_i = V2_25; // @[SWChisel.scala 200:22]
  assign array_26_io_q = io_q_26_b; // @[SWChisel.scala 220:19]
  assign array_26_io_r = 8'hc7 == r_count_26_io_out ? io_r_199_b : _GEN_5518; // @[SWChisel.scala 221:{19,19}]
  assign array_26_io_e_i = E_26; // @[SWChisel.scala 196:21]
  assign array_26_io_f_i = F_26; // @[SWChisel.scala 198:21]
  assign array_26_io_ve_i = V1_27; // @[SWChisel.scala 197:22]
  assign array_26_io_vf_i = V1_26; // @[SWChisel.scala 199:22]
  assign array_26_io_vv_i = V2_26; // @[SWChisel.scala 200:22]
  assign array_27_io_q = io_q_27_b; // @[SWChisel.scala 220:19]
  assign array_27_io_r = 8'hc7 == r_count_27_io_out ? io_r_199_b : _GEN_5718; // @[SWChisel.scala 221:{19,19}]
  assign array_27_io_e_i = E_27; // @[SWChisel.scala 196:21]
  assign array_27_io_f_i = F_27; // @[SWChisel.scala 198:21]
  assign array_27_io_ve_i = V1_28; // @[SWChisel.scala 197:22]
  assign array_27_io_vf_i = V1_27; // @[SWChisel.scala 199:22]
  assign array_27_io_vv_i = V2_27; // @[SWChisel.scala 200:22]
  assign array_28_io_q = io_q_28_b; // @[SWChisel.scala 220:19]
  assign array_28_io_r = 8'hc7 == r_count_28_io_out ? io_r_199_b : _GEN_5918; // @[SWChisel.scala 221:{19,19}]
  assign array_28_io_e_i = E_28; // @[SWChisel.scala 196:21]
  assign array_28_io_f_i = F_28; // @[SWChisel.scala 198:21]
  assign array_28_io_ve_i = V1_29; // @[SWChisel.scala 197:22]
  assign array_28_io_vf_i = V1_28; // @[SWChisel.scala 199:22]
  assign array_28_io_vv_i = V2_28; // @[SWChisel.scala 200:22]
  assign array_29_io_q = io_q_29_b; // @[SWChisel.scala 220:19]
  assign array_29_io_r = 8'hc7 == r_count_29_io_out ? io_r_199_b : _GEN_6118; // @[SWChisel.scala 221:{19,19}]
  assign array_29_io_e_i = E_29; // @[SWChisel.scala 196:21]
  assign array_29_io_f_i = F_29; // @[SWChisel.scala 198:21]
  assign array_29_io_ve_i = V1_30; // @[SWChisel.scala 197:22]
  assign array_29_io_vf_i = V1_29; // @[SWChisel.scala 199:22]
  assign array_29_io_vv_i = V2_29; // @[SWChisel.scala 200:22]
  assign array_30_io_q = io_q_30_b; // @[SWChisel.scala 220:19]
  assign array_30_io_r = 8'hc7 == r_count_30_io_out ? io_r_199_b : _GEN_6318; // @[SWChisel.scala 221:{19,19}]
  assign array_30_io_e_i = E_30; // @[SWChisel.scala 196:21]
  assign array_30_io_f_i = F_30; // @[SWChisel.scala 198:21]
  assign array_30_io_ve_i = V1_31; // @[SWChisel.scala 197:22]
  assign array_30_io_vf_i = V1_30; // @[SWChisel.scala 199:22]
  assign array_30_io_vv_i = V2_30; // @[SWChisel.scala 200:22]
  assign array_31_io_q = io_q_31_b; // @[SWChisel.scala 220:19]
  assign array_31_io_r = 8'hc7 == r_count_31_io_out ? io_r_199_b : _GEN_6518; // @[SWChisel.scala 221:{19,19}]
  assign array_31_io_e_i = E_31; // @[SWChisel.scala 196:21]
  assign array_31_io_f_i = F_31; // @[SWChisel.scala 198:21]
  assign array_31_io_ve_i = V1_32; // @[SWChisel.scala 197:22]
  assign array_31_io_vf_i = V1_31; // @[SWChisel.scala 199:22]
  assign array_31_io_vv_i = V2_31; // @[SWChisel.scala 200:22]
  assign array_32_io_q = io_q_32_b; // @[SWChisel.scala 220:19]
  assign array_32_io_r = 8'hc7 == r_count_32_io_out ? io_r_199_b : _GEN_6718; // @[SWChisel.scala 221:{19,19}]
  assign array_32_io_e_i = E_32; // @[SWChisel.scala 196:21]
  assign array_32_io_f_i = F_32; // @[SWChisel.scala 198:21]
  assign array_32_io_ve_i = V1_33; // @[SWChisel.scala 197:22]
  assign array_32_io_vf_i = V1_32; // @[SWChisel.scala 199:22]
  assign array_32_io_vv_i = V2_32; // @[SWChisel.scala 200:22]
  assign array_33_io_q = io_q_33_b; // @[SWChisel.scala 220:19]
  assign array_33_io_r = 8'hc7 == r_count_33_io_out ? io_r_199_b : _GEN_6918; // @[SWChisel.scala 221:{19,19}]
  assign array_33_io_e_i = E_33; // @[SWChisel.scala 196:21]
  assign array_33_io_f_i = F_33; // @[SWChisel.scala 198:21]
  assign array_33_io_ve_i = V1_34; // @[SWChisel.scala 197:22]
  assign array_33_io_vf_i = V1_33; // @[SWChisel.scala 199:22]
  assign array_33_io_vv_i = V2_33; // @[SWChisel.scala 200:22]
  assign array_34_io_q = io_q_34_b; // @[SWChisel.scala 220:19]
  assign array_34_io_r = 8'hc7 == r_count_34_io_out ? io_r_199_b : _GEN_7118; // @[SWChisel.scala 221:{19,19}]
  assign array_34_io_e_i = E_34; // @[SWChisel.scala 196:21]
  assign array_34_io_f_i = F_34; // @[SWChisel.scala 198:21]
  assign array_34_io_ve_i = V1_35; // @[SWChisel.scala 197:22]
  assign array_34_io_vf_i = V1_34; // @[SWChisel.scala 199:22]
  assign array_34_io_vv_i = V2_34; // @[SWChisel.scala 200:22]
  assign array_35_io_q = io_q_35_b; // @[SWChisel.scala 220:19]
  assign array_35_io_r = 8'hc7 == r_count_35_io_out ? io_r_199_b : _GEN_7318; // @[SWChisel.scala 221:{19,19}]
  assign array_35_io_e_i = E_35; // @[SWChisel.scala 196:21]
  assign array_35_io_f_i = F_35; // @[SWChisel.scala 198:21]
  assign array_35_io_ve_i = V1_36; // @[SWChisel.scala 197:22]
  assign array_35_io_vf_i = V1_35; // @[SWChisel.scala 199:22]
  assign array_35_io_vv_i = V2_35; // @[SWChisel.scala 200:22]
  assign array_36_io_q = io_q_36_b; // @[SWChisel.scala 220:19]
  assign array_36_io_r = 8'hc7 == r_count_36_io_out ? io_r_199_b : _GEN_7518; // @[SWChisel.scala 221:{19,19}]
  assign array_36_io_e_i = E_36; // @[SWChisel.scala 196:21]
  assign array_36_io_f_i = F_36; // @[SWChisel.scala 198:21]
  assign array_36_io_ve_i = V1_37; // @[SWChisel.scala 197:22]
  assign array_36_io_vf_i = V1_36; // @[SWChisel.scala 199:22]
  assign array_36_io_vv_i = V2_36; // @[SWChisel.scala 200:22]
  assign array_37_io_q = io_q_37_b; // @[SWChisel.scala 220:19]
  assign array_37_io_r = 8'hc7 == r_count_37_io_out ? io_r_199_b : _GEN_7718; // @[SWChisel.scala 221:{19,19}]
  assign array_37_io_e_i = E_37; // @[SWChisel.scala 196:21]
  assign array_37_io_f_i = F_37; // @[SWChisel.scala 198:21]
  assign array_37_io_ve_i = V1_38; // @[SWChisel.scala 197:22]
  assign array_37_io_vf_i = V1_37; // @[SWChisel.scala 199:22]
  assign array_37_io_vv_i = V2_37; // @[SWChisel.scala 200:22]
  assign array_38_io_q = io_q_38_b; // @[SWChisel.scala 220:19]
  assign array_38_io_r = 8'hc7 == r_count_38_io_out ? io_r_199_b : _GEN_7918; // @[SWChisel.scala 221:{19,19}]
  assign array_38_io_e_i = E_38; // @[SWChisel.scala 196:21]
  assign array_38_io_f_i = F_38; // @[SWChisel.scala 198:21]
  assign array_38_io_ve_i = V1_39; // @[SWChisel.scala 197:22]
  assign array_38_io_vf_i = V1_38; // @[SWChisel.scala 199:22]
  assign array_38_io_vv_i = V2_38; // @[SWChisel.scala 200:22]
  assign array_39_io_q = io_q_39_b; // @[SWChisel.scala 220:19]
  assign array_39_io_r = 8'hc7 == r_count_39_io_out ? io_r_199_b : _GEN_8118; // @[SWChisel.scala 221:{19,19}]
  assign array_39_io_e_i = E_39; // @[SWChisel.scala 196:21]
  assign array_39_io_f_i = F_39; // @[SWChisel.scala 198:21]
  assign array_39_io_ve_i = V1_40; // @[SWChisel.scala 197:22]
  assign array_39_io_vf_i = V1_39; // @[SWChisel.scala 199:22]
  assign array_39_io_vv_i = V2_39; // @[SWChisel.scala 200:22]
  assign r_count_0_clock = clock;
  assign r_count_0_reset = reset;
  assign r_count_0_io_en = start_reg_0; // @[SWChisel.scala 192:22]
  assign r_count_1_clock = clock;
  assign r_count_1_reset = reset;
  assign r_count_1_io_en = start_reg_1; // @[SWChisel.scala 192:22]
  assign r_count_2_clock = clock;
  assign r_count_2_reset = reset;
  assign r_count_2_io_en = start_reg_2; // @[SWChisel.scala 192:22]
  assign r_count_3_clock = clock;
  assign r_count_3_reset = reset;
  assign r_count_3_io_en = start_reg_3; // @[SWChisel.scala 192:22]
  assign r_count_4_clock = clock;
  assign r_count_4_reset = reset;
  assign r_count_4_io_en = start_reg_4; // @[SWChisel.scala 192:22]
  assign r_count_5_clock = clock;
  assign r_count_5_reset = reset;
  assign r_count_5_io_en = start_reg_5; // @[SWChisel.scala 192:22]
  assign r_count_6_clock = clock;
  assign r_count_6_reset = reset;
  assign r_count_6_io_en = start_reg_6; // @[SWChisel.scala 192:22]
  assign r_count_7_clock = clock;
  assign r_count_7_reset = reset;
  assign r_count_7_io_en = start_reg_7; // @[SWChisel.scala 192:22]
  assign r_count_8_clock = clock;
  assign r_count_8_reset = reset;
  assign r_count_8_io_en = start_reg_8; // @[SWChisel.scala 192:22]
  assign r_count_9_clock = clock;
  assign r_count_9_reset = reset;
  assign r_count_9_io_en = start_reg_9; // @[SWChisel.scala 192:22]
  assign r_count_10_clock = clock;
  assign r_count_10_reset = reset;
  assign r_count_10_io_en = start_reg_10; // @[SWChisel.scala 192:22]
  assign r_count_11_clock = clock;
  assign r_count_11_reset = reset;
  assign r_count_11_io_en = start_reg_11; // @[SWChisel.scala 192:22]
  assign r_count_12_clock = clock;
  assign r_count_12_reset = reset;
  assign r_count_12_io_en = start_reg_12; // @[SWChisel.scala 192:22]
  assign r_count_13_clock = clock;
  assign r_count_13_reset = reset;
  assign r_count_13_io_en = start_reg_13; // @[SWChisel.scala 192:22]
  assign r_count_14_clock = clock;
  assign r_count_14_reset = reset;
  assign r_count_14_io_en = start_reg_14; // @[SWChisel.scala 192:22]
  assign r_count_15_clock = clock;
  assign r_count_15_reset = reset;
  assign r_count_15_io_en = start_reg_15; // @[SWChisel.scala 192:22]
  assign r_count_16_clock = clock;
  assign r_count_16_reset = reset;
  assign r_count_16_io_en = start_reg_16; // @[SWChisel.scala 192:22]
  assign r_count_17_clock = clock;
  assign r_count_17_reset = reset;
  assign r_count_17_io_en = start_reg_17; // @[SWChisel.scala 192:22]
  assign r_count_18_clock = clock;
  assign r_count_18_reset = reset;
  assign r_count_18_io_en = start_reg_18; // @[SWChisel.scala 192:22]
  assign r_count_19_clock = clock;
  assign r_count_19_reset = reset;
  assign r_count_19_io_en = start_reg_19; // @[SWChisel.scala 192:22]
  assign r_count_20_clock = clock;
  assign r_count_20_reset = reset;
  assign r_count_20_io_en = start_reg_20; // @[SWChisel.scala 192:22]
  assign r_count_21_clock = clock;
  assign r_count_21_reset = reset;
  assign r_count_21_io_en = start_reg_21; // @[SWChisel.scala 192:22]
  assign r_count_22_clock = clock;
  assign r_count_22_reset = reset;
  assign r_count_22_io_en = start_reg_22; // @[SWChisel.scala 192:22]
  assign r_count_23_clock = clock;
  assign r_count_23_reset = reset;
  assign r_count_23_io_en = start_reg_23; // @[SWChisel.scala 192:22]
  assign r_count_24_clock = clock;
  assign r_count_24_reset = reset;
  assign r_count_24_io_en = start_reg_24; // @[SWChisel.scala 192:22]
  assign r_count_25_clock = clock;
  assign r_count_25_reset = reset;
  assign r_count_25_io_en = start_reg_25; // @[SWChisel.scala 192:22]
  assign r_count_26_clock = clock;
  assign r_count_26_reset = reset;
  assign r_count_26_io_en = start_reg_26; // @[SWChisel.scala 192:22]
  assign r_count_27_clock = clock;
  assign r_count_27_reset = reset;
  assign r_count_27_io_en = start_reg_27; // @[SWChisel.scala 192:22]
  assign r_count_28_clock = clock;
  assign r_count_28_reset = reset;
  assign r_count_28_io_en = start_reg_28; // @[SWChisel.scala 192:22]
  assign r_count_29_clock = clock;
  assign r_count_29_reset = reset;
  assign r_count_29_io_en = start_reg_29; // @[SWChisel.scala 192:22]
  assign r_count_30_clock = clock;
  assign r_count_30_reset = reset;
  assign r_count_30_io_en = start_reg_30; // @[SWChisel.scala 192:22]
  assign r_count_31_clock = clock;
  assign r_count_31_reset = reset;
  assign r_count_31_io_en = start_reg_31; // @[SWChisel.scala 192:22]
  assign r_count_32_clock = clock;
  assign r_count_32_reset = reset;
  assign r_count_32_io_en = start_reg_32; // @[SWChisel.scala 192:22]
  assign r_count_33_clock = clock;
  assign r_count_33_reset = reset;
  assign r_count_33_io_en = start_reg_33; // @[SWChisel.scala 192:22]
  assign r_count_34_clock = clock;
  assign r_count_34_reset = reset;
  assign r_count_34_io_en = start_reg_34; // @[SWChisel.scala 192:22]
  assign r_count_35_clock = clock;
  assign r_count_35_reset = reset;
  assign r_count_35_io_en = start_reg_35; // @[SWChisel.scala 192:22]
  assign r_count_36_clock = clock;
  assign r_count_36_reset = reset;
  assign r_count_36_io_en = start_reg_36; // @[SWChisel.scala 192:22]
  assign r_count_37_clock = clock;
  assign r_count_37_reset = reset;
  assign r_count_37_io_en = start_reg_37; // @[SWChisel.scala 192:22]
  assign r_count_38_clock = clock;
  assign r_count_38_reset = reset;
  assign r_count_38_io_en = start_reg_38; // @[SWChisel.scala 192:22]
  assign r_count_39_clock = clock;
  assign r_count_39_reset = reset;
  assign r_count_39_io_en = start_reg_39; // @[SWChisel.scala 192:22]
  assign max_clock = clock;
  assign max_reset = reset;
  assign max_io_start = start_reg_39; // @[SWChisel.scala 178:16]
  assign max_io_in = V1_40; // @[SWChisel.scala 177:13]
  always @(posedge clock) begin
    if (reset) begin // @[SWChisel.scala 162:18]
      E_0 <= -16'sh2; // @[SWChisel.scala 162:18]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      E_0 <= array_0_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_1 <= -16'sh3; // @[SWChisel.scala 162:18]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      E_1 <= array_1_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_2 <= -16'sh4; // @[SWChisel.scala 162:18]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      E_2 <= array_2_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_3 <= -16'sh5; // @[SWChisel.scala 162:18]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      E_3 <= array_3_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_4 <= -16'sh6; // @[SWChisel.scala 162:18]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      E_4 <= array_4_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_5 <= -16'sh7; // @[SWChisel.scala 162:18]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      E_5 <= array_5_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_6 <= -16'sh8; // @[SWChisel.scala 162:18]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      E_6 <= array_6_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_7 <= -16'sh9; // @[SWChisel.scala 162:18]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      E_7 <= array_7_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_8 <= -16'sha; // @[SWChisel.scala 162:18]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      E_8 <= array_8_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_9 <= -16'shb; // @[SWChisel.scala 162:18]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      E_9 <= array_9_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_10 <= -16'shc; // @[SWChisel.scala 162:18]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      E_10 <= array_10_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_11 <= -16'shd; // @[SWChisel.scala 162:18]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      E_11 <= array_11_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_12 <= -16'she; // @[SWChisel.scala 162:18]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      E_12 <= array_12_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_13 <= -16'shf; // @[SWChisel.scala 162:18]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      E_13 <= array_13_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_14 <= -16'sh10; // @[SWChisel.scala 162:18]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      E_14 <= array_14_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_15 <= -16'sh11; // @[SWChisel.scala 162:18]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      E_15 <= array_15_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_16 <= -16'sh12; // @[SWChisel.scala 162:18]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      E_16 <= array_16_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_17 <= -16'sh13; // @[SWChisel.scala 162:18]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      E_17 <= array_17_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_18 <= -16'sh14; // @[SWChisel.scala 162:18]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      E_18 <= array_18_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_19 <= -16'sh15; // @[SWChisel.scala 162:18]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      E_19 <= array_19_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_20 <= -16'sh16; // @[SWChisel.scala 162:18]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      E_20 <= array_20_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_21 <= -16'sh17; // @[SWChisel.scala 162:18]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      E_21 <= array_21_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_22 <= -16'sh18; // @[SWChisel.scala 162:18]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      E_22 <= array_22_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_23 <= -16'sh19; // @[SWChisel.scala 162:18]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      E_23 <= array_23_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_24 <= -16'sh1a; // @[SWChisel.scala 162:18]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      E_24 <= array_24_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_25 <= -16'sh1b; // @[SWChisel.scala 162:18]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      E_25 <= array_25_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_26 <= -16'sh1c; // @[SWChisel.scala 162:18]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      E_26 <= array_26_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_27 <= -16'sh1d; // @[SWChisel.scala 162:18]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      E_27 <= array_27_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_28 <= -16'sh1e; // @[SWChisel.scala 162:18]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      E_28 <= array_28_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_29 <= -16'sh1f; // @[SWChisel.scala 162:18]
    end else if (start_reg_29) begin // @[SWChisel.scala 207:25]
      E_29 <= array_29_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_30 <= -16'sh20; // @[SWChisel.scala 162:18]
    end else if (start_reg_30) begin // @[SWChisel.scala 207:25]
      E_30 <= array_30_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_31 <= -16'sh21; // @[SWChisel.scala 162:18]
    end else if (start_reg_31) begin // @[SWChisel.scala 207:25]
      E_31 <= array_31_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_32 <= -16'sh22; // @[SWChisel.scala 162:18]
    end else if (start_reg_32) begin // @[SWChisel.scala 207:25]
      E_32 <= array_32_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_33 <= -16'sh23; // @[SWChisel.scala 162:18]
    end else if (start_reg_33) begin // @[SWChisel.scala 207:25]
      E_33 <= array_33_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_34 <= -16'sh24; // @[SWChisel.scala 162:18]
    end else if (start_reg_34) begin // @[SWChisel.scala 207:25]
      E_34 <= array_34_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_35 <= -16'sh25; // @[SWChisel.scala 162:18]
    end else if (start_reg_35) begin // @[SWChisel.scala 207:25]
      E_35 <= array_35_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_36 <= -16'sh26; // @[SWChisel.scala 162:18]
    end else if (start_reg_36) begin // @[SWChisel.scala 207:25]
      E_36 <= array_36_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_37 <= -16'sh27; // @[SWChisel.scala 162:18]
    end else if (start_reg_37) begin // @[SWChisel.scala 207:25]
      E_37 <= array_37_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_38 <= -16'sh28; // @[SWChisel.scala 162:18]
    end else if (start_reg_38) begin // @[SWChisel.scala 207:25]
      E_38 <= array_38_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_39 <= -16'sh29; // @[SWChisel.scala 162:18]
    end else if (start_reg_39) begin // @[SWChisel.scala 207:25]
      E_39 <= array_39_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_1 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      F_1 <= array_0_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_2 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      F_2 <= array_1_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_3 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      F_3 <= array_2_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_4 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      F_4 <= array_3_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_5 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      F_5 <= array_4_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_6 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      F_6 <= array_5_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_7 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      F_7 <= array_6_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_8 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      F_8 <= array_7_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_9 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      F_9 <= array_8_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_10 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      F_10 <= array_9_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_11 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      F_11 <= array_10_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_12 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      F_12 <= array_11_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_13 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      F_13 <= array_12_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_14 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      F_14 <= array_13_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_15 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      F_15 <= array_14_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_16 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      F_16 <= array_15_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_17 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      F_17 <= array_16_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_18 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      F_18 <= array_17_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_19 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      F_19 <= array_18_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_20 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      F_20 <= array_19_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_21 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      F_21 <= array_20_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_22 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      F_22 <= array_21_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_23 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      F_23 <= array_22_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_24 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      F_24 <= array_23_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_25 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      F_25 <= array_24_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_26 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      F_26 <= array_25_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_27 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      F_27 <= array_26_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_28 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      F_28 <= array_27_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_29 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      F_29 <= array_28_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_30 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_29) begin // @[SWChisel.scala 207:25]
      F_30 <= array_29_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_31 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_30) begin // @[SWChisel.scala 207:25]
      F_31 <= array_30_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_32 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_31) begin // @[SWChisel.scala 207:25]
      F_32 <= array_31_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_33 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_32) begin // @[SWChisel.scala 207:25]
      F_33 <= array_32_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_34 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_33) begin // @[SWChisel.scala 207:25]
      F_34 <= array_33_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_35 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_34) begin // @[SWChisel.scala 207:25]
      F_35 <= array_34_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_36 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_35) begin // @[SWChisel.scala 207:25]
      F_36 <= array_35_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_37 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_36) begin // @[SWChisel.scala 207:25]
      F_37 <= array_36_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_38 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_37) begin // @[SWChisel.scala 207:25]
      F_38 <= array_37_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_39 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_38) begin // @[SWChisel.scala 207:25]
      F_39 <= array_38_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_0 <= -16'sh1; // @[SWChisel.scala 164:19]
    end else begin
      V1_0 <= 16'sh0; // @[SWChisel.scala 165:9]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_1 <= -16'sh2; // @[SWChisel.scala 164:19]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      V1_1 <= array_0_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_2 <= -16'sh3; // @[SWChisel.scala 164:19]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      V1_2 <= array_1_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_3 <= -16'sh4; // @[SWChisel.scala 164:19]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      V1_3 <= array_2_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_4 <= -16'sh5; // @[SWChisel.scala 164:19]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      V1_4 <= array_3_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_5 <= -16'sh6; // @[SWChisel.scala 164:19]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      V1_5 <= array_4_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_6 <= -16'sh7; // @[SWChisel.scala 164:19]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      V1_6 <= array_5_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_7 <= -16'sh8; // @[SWChisel.scala 164:19]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      V1_7 <= array_6_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_8 <= -16'sh9; // @[SWChisel.scala 164:19]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      V1_8 <= array_7_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_9 <= -16'sha; // @[SWChisel.scala 164:19]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      V1_9 <= array_8_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_10 <= -16'shb; // @[SWChisel.scala 164:19]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      V1_10 <= array_9_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_11 <= -16'shc; // @[SWChisel.scala 164:19]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      V1_11 <= array_10_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_12 <= -16'shd; // @[SWChisel.scala 164:19]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      V1_12 <= array_11_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_13 <= -16'she; // @[SWChisel.scala 164:19]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      V1_13 <= array_12_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_14 <= -16'shf; // @[SWChisel.scala 164:19]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      V1_14 <= array_13_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_15 <= -16'sh10; // @[SWChisel.scala 164:19]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      V1_15 <= array_14_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_16 <= -16'sh11; // @[SWChisel.scala 164:19]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      V1_16 <= array_15_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_17 <= -16'sh12; // @[SWChisel.scala 164:19]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      V1_17 <= array_16_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_18 <= -16'sh13; // @[SWChisel.scala 164:19]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      V1_18 <= array_17_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_19 <= -16'sh14; // @[SWChisel.scala 164:19]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      V1_19 <= array_18_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_20 <= -16'sh15; // @[SWChisel.scala 164:19]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      V1_20 <= array_19_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_21 <= -16'sh16; // @[SWChisel.scala 164:19]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      V1_21 <= array_20_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_22 <= -16'sh17; // @[SWChisel.scala 164:19]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      V1_22 <= array_21_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_23 <= -16'sh18; // @[SWChisel.scala 164:19]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      V1_23 <= array_22_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_24 <= -16'sh19; // @[SWChisel.scala 164:19]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      V1_24 <= array_23_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_25 <= -16'sh1a; // @[SWChisel.scala 164:19]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      V1_25 <= array_24_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_26 <= -16'sh1b; // @[SWChisel.scala 164:19]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      V1_26 <= array_25_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_27 <= -16'sh1c; // @[SWChisel.scala 164:19]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      V1_27 <= array_26_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_28 <= -16'sh1d; // @[SWChisel.scala 164:19]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      V1_28 <= array_27_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_29 <= -16'sh1e; // @[SWChisel.scala 164:19]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      V1_29 <= array_28_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_30 <= -16'sh1f; // @[SWChisel.scala 164:19]
    end else if (start_reg_29) begin // @[SWChisel.scala 207:25]
      V1_30 <= array_29_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_31 <= -16'sh20; // @[SWChisel.scala 164:19]
    end else if (start_reg_30) begin // @[SWChisel.scala 207:25]
      V1_31 <= array_30_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_32 <= -16'sh21; // @[SWChisel.scala 164:19]
    end else if (start_reg_31) begin // @[SWChisel.scala 207:25]
      V1_32 <= array_31_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_33 <= -16'sh22; // @[SWChisel.scala 164:19]
    end else if (start_reg_32) begin // @[SWChisel.scala 207:25]
      V1_33 <= array_32_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_34 <= -16'sh23; // @[SWChisel.scala 164:19]
    end else if (start_reg_33) begin // @[SWChisel.scala 207:25]
      V1_34 <= array_33_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_35 <= -16'sh24; // @[SWChisel.scala 164:19]
    end else if (start_reg_34) begin // @[SWChisel.scala 207:25]
      V1_35 <= array_34_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_36 <= -16'sh25; // @[SWChisel.scala 164:19]
    end else if (start_reg_35) begin // @[SWChisel.scala 207:25]
      V1_36 <= array_35_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_37 <= -16'sh26; // @[SWChisel.scala 164:19]
    end else if (start_reg_36) begin // @[SWChisel.scala 207:25]
      V1_37 <= array_36_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_38 <= -16'sh27; // @[SWChisel.scala 164:19]
    end else if (start_reg_37) begin // @[SWChisel.scala 207:25]
      V1_38 <= array_37_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_39 <= -16'sh28; // @[SWChisel.scala 164:19]
    end else if (start_reg_38) begin // @[SWChisel.scala 207:25]
      V1_39 <= array_38_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_40 <= -16'sh29; // @[SWChisel.scala 164:19]
    end else if (start_reg_39) begin // @[SWChisel.scala 207:25]
      V1_40 <= array_39_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_0 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_0 <= V1_0; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_1 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_1 <= V1_1; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_2 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_2 <= V1_2; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_3 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_3 <= V1_3; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_4 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_4 <= V1_4; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_5 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_5 <= V1_5; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_6 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_6 <= V1_6; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_7 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_7 <= V1_7; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_8 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_8 <= V1_8; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_9 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_9 <= V1_9; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_10 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_10 <= V1_10; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_11 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_11 <= V1_11; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_12 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_12 <= V1_12; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_13 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_13 <= V1_13; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_14 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_14 <= V1_14; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_15 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_15 <= V1_15; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_16 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_16 <= V1_16; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_17 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_17 <= V1_17; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_18 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_18 <= V1_18; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_19 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_19 <= V1_19; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_20 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_20 <= V1_20; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_21 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_21 <= V1_21; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_22 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_22 <= V1_22; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_23 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_23 <= V1_23; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_24 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_24 <= V1_24; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_25 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_25 <= V1_25; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_26 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_26 <= V1_26; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_27 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_27 <= V1_27; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_28 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_28 <= V1_28; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_29 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_29 <= V1_29; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_30 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_30 <= V1_30; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_31 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_31 <= V1_31; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_32 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_32 <= V1_32; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_33 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_33 <= V1_33; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_34 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_34 <= V1_34; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_35 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_35 <= V1_35; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_36 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_36 <= V1_36; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_37 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_37 <= V1_37; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_38 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_38 <= V1_38; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_39 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_39 <= V1_39; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_0 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_0 <= io_start; // @[SWChisel.scala 185:16]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_1 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_1 <= start_reg_0; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_2 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_2 <= start_reg_1; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_3 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_3 <= start_reg_2; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_4 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_4 <= start_reg_3; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_5 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_5 <= start_reg_4; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_6 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_6 <= start_reg_5; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_7 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_7 <= start_reg_6; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_8 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_8 <= start_reg_7; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_9 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_9 <= start_reg_8; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_10 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_10 <= start_reg_9; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_11 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_11 <= start_reg_10; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_12 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_12 <= start_reg_11; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_13 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_13 <= start_reg_12; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_14 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_14 <= start_reg_13; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_15 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_15 <= start_reg_14; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_16 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_16 <= start_reg_15; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_17 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_17 <= start_reg_16; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_18 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_18 <= start_reg_17; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_19 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_19 <= start_reg_18; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_20 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_20 <= start_reg_19; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_21 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_21 <= start_reg_20; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_22 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_22 <= start_reg_21; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_23 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_23 <= start_reg_22; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_24 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_24 <= start_reg_23; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_25 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_25 <= start_reg_24; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_26 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_26 <= start_reg_25; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_27 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_27 <= start_reg_26; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_28 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_28 <= start_reg_27; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_29 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_29 <= start_reg_28; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_30 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_30 <= start_reg_29; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_31 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_31 <= start_reg_30; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_32 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_32 <= start_reg_31; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_33 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_33 <= start_reg_32; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_34 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_34 <= start_reg_33; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_35 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_35 <= start_reg_34; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_36 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_36 <= start_reg_35; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_37 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_37 <= start_reg_36; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_38 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_38 <= start_reg_37; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_39 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_39 <= start_reg_38; // @[SWChisel.scala 187:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  E_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  E_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  E_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  E_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  E_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  E_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  E_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  E_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  E_8 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  E_9 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  E_10 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  E_11 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  E_12 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  E_13 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  E_14 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  E_15 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  E_16 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  E_17 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  E_18 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  E_19 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  E_20 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  E_21 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  E_22 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  E_23 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  E_24 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  E_25 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  E_26 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  E_27 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  E_28 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  E_29 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  E_30 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  E_31 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  E_32 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  E_33 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  E_34 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  E_35 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  E_36 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  E_37 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  E_38 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  E_39 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  F_1 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  F_2 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  F_3 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  F_4 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  F_5 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  F_6 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  F_7 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  F_8 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  F_9 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  F_10 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  F_11 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  F_12 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  F_13 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  F_14 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  F_15 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  F_16 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  F_17 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  F_18 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  F_19 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  F_20 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  F_21 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  F_22 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  F_23 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  F_24 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  F_25 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  F_26 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  F_27 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  F_28 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  F_29 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  F_30 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  F_31 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  F_32 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  F_33 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  F_34 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  F_35 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  F_36 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  F_37 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  F_38 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  F_39 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  V1_0 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  V1_1 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  V1_2 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  V1_3 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  V1_4 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  V1_5 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  V1_6 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  V1_7 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  V1_8 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  V1_9 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  V1_10 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  V1_11 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  V1_12 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  V1_13 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  V1_14 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  V1_15 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  V1_16 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  V1_17 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  V1_18 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  V1_19 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  V1_20 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  V1_21 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  V1_22 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  V1_23 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  V1_24 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  V1_25 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  V1_26 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  V1_27 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  V1_28 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  V1_29 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  V1_30 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  V1_31 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  V1_32 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  V1_33 = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  V1_34 = _RAND_113[15:0];
  _RAND_114 = {1{`RANDOM}};
  V1_35 = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  V1_36 = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  V1_37 = _RAND_116[15:0];
  _RAND_117 = {1{`RANDOM}};
  V1_38 = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  V1_39 = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  V1_40 = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  V2_0 = _RAND_120[15:0];
  _RAND_121 = {1{`RANDOM}};
  V2_1 = _RAND_121[15:0];
  _RAND_122 = {1{`RANDOM}};
  V2_2 = _RAND_122[15:0];
  _RAND_123 = {1{`RANDOM}};
  V2_3 = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  V2_4 = _RAND_124[15:0];
  _RAND_125 = {1{`RANDOM}};
  V2_5 = _RAND_125[15:0];
  _RAND_126 = {1{`RANDOM}};
  V2_6 = _RAND_126[15:0];
  _RAND_127 = {1{`RANDOM}};
  V2_7 = _RAND_127[15:0];
  _RAND_128 = {1{`RANDOM}};
  V2_8 = _RAND_128[15:0];
  _RAND_129 = {1{`RANDOM}};
  V2_9 = _RAND_129[15:0];
  _RAND_130 = {1{`RANDOM}};
  V2_10 = _RAND_130[15:0];
  _RAND_131 = {1{`RANDOM}};
  V2_11 = _RAND_131[15:0];
  _RAND_132 = {1{`RANDOM}};
  V2_12 = _RAND_132[15:0];
  _RAND_133 = {1{`RANDOM}};
  V2_13 = _RAND_133[15:0];
  _RAND_134 = {1{`RANDOM}};
  V2_14 = _RAND_134[15:0];
  _RAND_135 = {1{`RANDOM}};
  V2_15 = _RAND_135[15:0];
  _RAND_136 = {1{`RANDOM}};
  V2_16 = _RAND_136[15:0];
  _RAND_137 = {1{`RANDOM}};
  V2_17 = _RAND_137[15:0];
  _RAND_138 = {1{`RANDOM}};
  V2_18 = _RAND_138[15:0];
  _RAND_139 = {1{`RANDOM}};
  V2_19 = _RAND_139[15:0];
  _RAND_140 = {1{`RANDOM}};
  V2_20 = _RAND_140[15:0];
  _RAND_141 = {1{`RANDOM}};
  V2_21 = _RAND_141[15:0];
  _RAND_142 = {1{`RANDOM}};
  V2_22 = _RAND_142[15:0];
  _RAND_143 = {1{`RANDOM}};
  V2_23 = _RAND_143[15:0];
  _RAND_144 = {1{`RANDOM}};
  V2_24 = _RAND_144[15:0];
  _RAND_145 = {1{`RANDOM}};
  V2_25 = _RAND_145[15:0];
  _RAND_146 = {1{`RANDOM}};
  V2_26 = _RAND_146[15:0];
  _RAND_147 = {1{`RANDOM}};
  V2_27 = _RAND_147[15:0];
  _RAND_148 = {1{`RANDOM}};
  V2_28 = _RAND_148[15:0];
  _RAND_149 = {1{`RANDOM}};
  V2_29 = _RAND_149[15:0];
  _RAND_150 = {1{`RANDOM}};
  V2_30 = _RAND_150[15:0];
  _RAND_151 = {1{`RANDOM}};
  V2_31 = _RAND_151[15:0];
  _RAND_152 = {1{`RANDOM}};
  V2_32 = _RAND_152[15:0];
  _RAND_153 = {1{`RANDOM}};
  V2_33 = _RAND_153[15:0];
  _RAND_154 = {1{`RANDOM}};
  V2_34 = _RAND_154[15:0];
  _RAND_155 = {1{`RANDOM}};
  V2_35 = _RAND_155[15:0];
  _RAND_156 = {1{`RANDOM}};
  V2_36 = _RAND_156[15:0];
  _RAND_157 = {1{`RANDOM}};
  V2_37 = _RAND_157[15:0];
  _RAND_158 = {1{`RANDOM}};
  V2_38 = _RAND_158[15:0];
  _RAND_159 = {1{`RANDOM}};
  V2_39 = _RAND_159[15:0];
  _RAND_160 = {1{`RANDOM}};
  start_reg_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  start_reg_1 = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  start_reg_2 = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  start_reg_3 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  start_reg_4 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  start_reg_5 = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  start_reg_6 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  start_reg_7 = _RAND_167[0:0];
  _RAND_168 = {1{`RANDOM}};
  start_reg_8 = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  start_reg_9 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  start_reg_10 = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  start_reg_11 = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  start_reg_12 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  start_reg_13 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  start_reg_14 = _RAND_174[0:0];
  _RAND_175 = {1{`RANDOM}};
  start_reg_15 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  start_reg_16 = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  start_reg_17 = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  start_reg_18 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  start_reg_19 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  start_reg_20 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  start_reg_21 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  start_reg_22 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  start_reg_23 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  start_reg_24 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  start_reg_25 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  start_reg_26 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  start_reg_27 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  start_reg_28 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  start_reg_29 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  start_reg_30 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  start_reg_31 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  start_reg_32 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  start_reg_33 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  start_reg_34 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  start_reg_35 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  start_reg_36 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  start_reg_37 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  start_reg_38 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  start_reg_39 = _RAND_199[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
