module SWCell(
  input  [1:0]  io_q,
  input  [1:0]  io_r,
  input  [15:0] io_e_i,
  input  [15:0] io_f_i,
  input  [15:0] io_ve_i,
  input  [15:0] io_vf_i,
  input  [15:0] io_vv_i,
  output [15:0] io_e_o,
  output [15:0] io_f_o,
  output [15:0] io_v_o
);
  wire [15:0] _T_2 = $signed(io_ve_i) - 16'sh2; // @[SWChisel.scala 78:17]
  wire [15:0] _T_5 = $signed(io_e_i) - 16'sh1; // @[SWChisel.scala 78:39]
  wire [15:0] e_max = $signed(_T_2) >= $signed(_T_5) ? $signed(_T_2) : $signed(_T_5); // @[SWChisel.scala 78:51 79:11 81:11]
  wire [15:0] _T_9 = $signed(io_vf_i) - 16'sh2; // @[SWChisel.scala 85:17]
  wire [15:0] _T_12 = $signed(io_f_i) - 16'sh1; // @[SWChisel.scala 85:38]
  wire [15:0] f_max = $signed(_T_9) > $signed(_T_12) ? $signed(_T_9) : $signed(_T_12); // @[SWChisel.scala 85:50 86:11 88:11]
  wire [15:0] ef_temp = $signed(e_max) > $signed(f_max) ? $signed(e_max) : $signed(f_max); // @[SWChisel.scala 92:24 93:13 95:13]
  wire [15:0] _v_temp_T_2 = $signed(io_vv_i) + 16'sh2; // @[SWChisel.scala 100:23]
  wire [15:0] _v_temp_T_5 = $signed(io_vv_i) - 16'sh2; // @[SWChisel.scala 102:23]
  wire [15:0] v_temp = io_q == io_r ? $signed(_v_temp_T_2) : $signed(_v_temp_T_5); // @[SWChisel.scala 100:12 102:12 99:24]
  assign io_e_o = $signed(_T_2) >= $signed(_T_5) ? $signed(_T_2) : $signed(_T_5); // @[SWChisel.scala 78:51 79:11 81:11]
  assign io_f_o = $signed(_T_9) > $signed(_T_12) ? $signed(_T_9) : $signed(_T_12); // @[SWChisel.scala 85:50 86:11 88:11]
  assign io_v_o = $signed(v_temp) > $signed(ef_temp) ? $signed(v_temp) : $signed(ef_temp); // @[SWChisel.scala 106:27 107:11 109:11]
endmodule
module MyCounter(
  input        clock,
  input        reset,
  input        io_en,
  output [6:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [6:0] _io_out_T_2 = io_out + 7'h1; // @[SWChisel.scala 155:55]
  reg [6:0] io_out_r; // @[Reg.scala 35:20]
  assign io_out = io_out_r; // @[SWChisel.scala 155:12]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 35:20]
      io_out_r <= 7'h0; // @[Reg.scala 35:20]
    end else if (io_en) begin // @[Reg.scala 36:18]
      if (io_out < 7'h64) begin // @[SWChisel.scala 155:28]
        io_out_r <= _io_out_T_2;
      end else begin
        io_out_r <= 7'h0;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_out_r = _RAND_0[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MAX(
  input         clock,
  input         reset,
  input         io_start,
  input  [15:0] io_in,
  output        io_done,
  output [15:0] io_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] max; // @[SWChisel.scala 122:20]
  reg [6:0] counter; // @[SWChisel.scala 133:24]
  wire [6:0] _counter_T_1 = counter - 7'h1; // @[SWChisel.scala 135:24]
  assign io_done = counter == 7'h0; // @[SWChisel.scala 141:17]
  assign io_out = max; // @[SWChisel.scala 123:10]
  always @(posedge clock) begin
    if (reset) begin // @[SWChisel.scala 122:20]
      max <= 16'sh8000; // @[SWChisel.scala 122:20]
    end else if ($signed(io_in) > $signed(max)) begin // @[SWChisel.scala 126:22]
      max <= io_in; // @[SWChisel.scala 127:9]
    end
    if (reset) begin // @[SWChisel.scala 133:24]
      counter <= 7'h65; // @[SWChisel.scala 133:24]
    end else if (counter == 7'h0) begin // @[SWChisel.scala 141:26]
      counter <= 7'h0; // @[SWChisel.scala 143:13]
    end else if (io_start) begin // @[SWChisel.scala 134:19]
      counter <= _counter_T_1; // @[SWChisel.scala 135:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  max = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  counter = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SW(
  input         clock,
  input         reset,
  input  [1:0]  io_q_0_b,
  input  [1:0]  io_q_1_b,
  input  [1:0]  io_q_2_b,
  input  [1:0]  io_q_3_b,
  input  [1:0]  io_q_4_b,
  input  [1:0]  io_q_5_b,
  input  [1:0]  io_q_6_b,
  input  [1:0]  io_q_7_b,
  input  [1:0]  io_q_8_b,
  input  [1:0]  io_q_9_b,
  input  [1:0]  io_q_10_b,
  input  [1:0]  io_q_11_b,
  input  [1:0]  io_q_12_b,
  input  [1:0]  io_q_13_b,
  input  [1:0]  io_q_14_b,
  input  [1:0]  io_q_15_b,
  input  [1:0]  io_q_16_b,
  input  [1:0]  io_q_17_b,
  input  [1:0]  io_q_18_b,
  input  [1:0]  io_q_19_b,
  input  [1:0]  io_q_20_b,
  input  [1:0]  io_q_21_b,
  input  [1:0]  io_q_22_b,
  input  [1:0]  io_q_23_b,
  input  [1:0]  io_q_24_b,
  input  [1:0]  io_q_25_b,
  input  [1:0]  io_q_26_b,
  input  [1:0]  io_q_27_b,
  input  [1:0]  io_q_28_b,
  input  [1:0]  io_q_29_b,
  input  [1:0]  io_q_30_b,
  input  [1:0]  io_q_31_b,
  input  [1:0]  io_q_32_b,
  input  [1:0]  io_q_33_b,
  input  [1:0]  io_q_34_b,
  input  [1:0]  io_q_35_b,
  input  [1:0]  io_q_36_b,
  input  [1:0]  io_q_37_b,
  input  [1:0]  io_q_38_b,
  input  [1:0]  io_q_39_b,
  input  [1:0]  io_q_40_b,
  input  [1:0]  io_q_41_b,
  input  [1:0]  io_q_42_b,
  input  [1:0]  io_q_43_b,
  input  [1:0]  io_q_44_b,
  input  [1:0]  io_q_45_b,
  input  [1:0]  io_q_46_b,
  input  [1:0]  io_q_47_b,
  input  [1:0]  io_q_48_b,
  input  [1:0]  io_q_49_b,
  input  [1:0]  io_r_0_b,
  input  [1:0]  io_r_1_b,
  input  [1:0]  io_r_2_b,
  input  [1:0]  io_r_3_b,
  input  [1:0]  io_r_4_b,
  input  [1:0]  io_r_5_b,
  input  [1:0]  io_r_6_b,
  input  [1:0]  io_r_7_b,
  input  [1:0]  io_r_8_b,
  input  [1:0]  io_r_9_b,
  input  [1:0]  io_r_10_b,
  input  [1:0]  io_r_11_b,
  input  [1:0]  io_r_12_b,
  input  [1:0]  io_r_13_b,
  input  [1:0]  io_r_14_b,
  input  [1:0]  io_r_15_b,
  input  [1:0]  io_r_16_b,
  input  [1:0]  io_r_17_b,
  input  [1:0]  io_r_18_b,
  input  [1:0]  io_r_19_b,
  input  [1:0]  io_r_20_b,
  input  [1:0]  io_r_21_b,
  input  [1:0]  io_r_22_b,
  input  [1:0]  io_r_23_b,
  input  [1:0]  io_r_24_b,
  input  [1:0]  io_r_25_b,
  input  [1:0]  io_r_26_b,
  input  [1:0]  io_r_27_b,
  input  [1:0]  io_r_28_b,
  input  [1:0]  io_r_29_b,
  input  [1:0]  io_r_30_b,
  input  [1:0]  io_r_31_b,
  input  [1:0]  io_r_32_b,
  input  [1:0]  io_r_33_b,
  input  [1:0]  io_r_34_b,
  input  [1:0]  io_r_35_b,
  input  [1:0]  io_r_36_b,
  input  [1:0]  io_r_37_b,
  input  [1:0]  io_r_38_b,
  input  [1:0]  io_r_39_b,
  input  [1:0]  io_r_40_b,
  input  [1:0]  io_r_41_b,
  input  [1:0]  io_r_42_b,
  input  [1:0]  io_r_43_b,
  input  [1:0]  io_r_44_b,
  input  [1:0]  io_r_45_b,
  input  [1:0]  io_r_46_b,
  input  [1:0]  io_r_47_b,
  input  [1:0]  io_r_48_b,
  input  [1:0]  io_r_49_b,
  input  [1:0]  io_r_50_b,
  input  [1:0]  io_r_51_b,
  input  [1:0]  io_r_52_b,
  input  [1:0]  io_r_53_b,
  input  [1:0]  io_r_54_b,
  input  [1:0]  io_r_55_b,
  input  [1:0]  io_r_56_b,
  input  [1:0]  io_r_57_b,
  input  [1:0]  io_r_58_b,
  input  [1:0]  io_r_59_b,
  input  [1:0]  io_r_60_b,
  input  [1:0]  io_r_61_b,
  input  [1:0]  io_r_62_b,
  input  [1:0]  io_r_63_b,
  input  [1:0]  io_r_64_b,
  input  [1:0]  io_r_65_b,
  input  [1:0]  io_r_66_b,
  input  [1:0]  io_r_67_b,
  input  [1:0]  io_r_68_b,
  input  [1:0]  io_r_69_b,
  input  [1:0]  io_r_70_b,
  input  [1:0]  io_r_71_b,
  input  [1:0]  io_r_72_b,
  input  [1:0]  io_r_73_b,
  input  [1:0]  io_r_74_b,
  input  [1:0]  io_r_75_b,
  input  [1:0]  io_r_76_b,
  input  [1:0]  io_r_77_b,
  input  [1:0]  io_r_78_b,
  input  [1:0]  io_r_79_b,
  input  [1:0]  io_r_80_b,
  input  [1:0]  io_r_81_b,
  input  [1:0]  io_r_82_b,
  input  [1:0]  io_r_83_b,
  input  [1:0]  io_r_84_b,
  input  [1:0]  io_r_85_b,
  input  [1:0]  io_r_86_b,
  input  [1:0]  io_r_87_b,
  input  [1:0]  io_r_88_b,
  input  [1:0]  io_r_89_b,
  input  [1:0]  io_r_90_b,
  input  [1:0]  io_r_91_b,
  input  [1:0]  io_r_92_b,
  input  [1:0]  io_r_93_b,
  input  [1:0]  io_r_94_b,
  input  [1:0]  io_r_95_b,
  input  [1:0]  io_r_96_b,
  input  [1:0]  io_r_97_b,
  input  [1:0]  io_r_98_b,
  input  [1:0]  io_r_99_b,
  input         io_start,
  output [15:0] io_result,
  output        io_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
`endif // RANDOMIZE_REG_INIT
  wire [1:0] array_0_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_0_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_0_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_1_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_1_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_1_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_2_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_2_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_2_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_3_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_3_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_3_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_4_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_4_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_4_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_5_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_5_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_5_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_6_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_6_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_6_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_7_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_7_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_7_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_8_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_8_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_8_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_9_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_9_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_9_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_10_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_10_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_10_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_11_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_11_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_11_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_12_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_12_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_12_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_13_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_13_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_13_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_14_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_14_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_14_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_15_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_15_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_15_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_16_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_16_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_16_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_17_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_17_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_17_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_18_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_18_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_18_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_19_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_19_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_19_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_20_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_20_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_20_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_21_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_21_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_21_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_22_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_22_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_22_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_23_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_23_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_23_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_24_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_24_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_24_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_25_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_25_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_25_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_26_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_26_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_26_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_27_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_27_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_27_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_28_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_28_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_28_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_29_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_29_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_29_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_30_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_30_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_30_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_31_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_31_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_31_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_32_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_32_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_32_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_33_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_33_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_33_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_34_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_34_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_34_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_35_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_35_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_35_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_36_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_36_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_36_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_37_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_37_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_37_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_38_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_38_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_38_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_39_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_39_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_39_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_40_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_40_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_40_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_41_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_41_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_41_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_42_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_42_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_42_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_43_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_43_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_43_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_44_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_44_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_44_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_45_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_45_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_45_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_46_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_46_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_46_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_47_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_47_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_47_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_48_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_48_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_48_io_v_o; // @[SWChisel.scala 170:39]
  wire [1:0] array_49_io_q; // @[SWChisel.scala 170:39]
  wire [1:0] array_49_io_r; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_e_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_f_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_ve_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_vf_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_vv_i; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_e_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_f_o; // @[SWChisel.scala 170:39]
  wire [15:0] array_49_io_v_o; // @[SWChisel.scala 170:39]
  wire  r_count_0_clock; // @[SWChisel.scala 171:41]
  wire  r_count_0_reset; // @[SWChisel.scala 171:41]
  wire  r_count_0_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_0_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_1_clock; // @[SWChisel.scala 171:41]
  wire  r_count_1_reset; // @[SWChisel.scala 171:41]
  wire  r_count_1_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_1_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_2_clock; // @[SWChisel.scala 171:41]
  wire  r_count_2_reset; // @[SWChisel.scala 171:41]
  wire  r_count_2_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_2_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_3_clock; // @[SWChisel.scala 171:41]
  wire  r_count_3_reset; // @[SWChisel.scala 171:41]
  wire  r_count_3_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_3_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_4_clock; // @[SWChisel.scala 171:41]
  wire  r_count_4_reset; // @[SWChisel.scala 171:41]
  wire  r_count_4_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_4_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_5_clock; // @[SWChisel.scala 171:41]
  wire  r_count_5_reset; // @[SWChisel.scala 171:41]
  wire  r_count_5_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_5_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_6_clock; // @[SWChisel.scala 171:41]
  wire  r_count_6_reset; // @[SWChisel.scala 171:41]
  wire  r_count_6_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_6_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_7_clock; // @[SWChisel.scala 171:41]
  wire  r_count_7_reset; // @[SWChisel.scala 171:41]
  wire  r_count_7_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_7_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_8_clock; // @[SWChisel.scala 171:41]
  wire  r_count_8_reset; // @[SWChisel.scala 171:41]
  wire  r_count_8_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_8_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_9_clock; // @[SWChisel.scala 171:41]
  wire  r_count_9_reset; // @[SWChisel.scala 171:41]
  wire  r_count_9_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_9_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_10_clock; // @[SWChisel.scala 171:41]
  wire  r_count_10_reset; // @[SWChisel.scala 171:41]
  wire  r_count_10_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_10_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_11_clock; // @[SWChisel.scala 171:41]
  wire  r_count_11_reset; // @[SWChisel.scala 171:41]
  wire  r_count_11_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_11_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_12_clock; // @[SWChisel.scala 171:41]
  wire  r_count_12_reset; // @[SWChisel.scala 171:41]
  wire  r_count_12_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_12_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_13_clock; // @[SWChisel.scala 171:41]
  wire  r_count_13_reset; // @[SWChisel.scala 171:41]
  wire  r_count_13_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_13_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_14_clock; // @[SWChisel.scala 171:41]
  wire  r_count_14_reset; // @[SWChisel.scala 171:41]
  wire  r_count_14_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_14_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_15_clock; // @[SWChisel.scala 171:41]
  wire  r_count_15_reset; // @[SWChisel.scala 171:41]
  wire  r_count_15_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_15_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_16_clock; // @[SWChisel.scala 171:41]
  wire  r_count_16_reset; // @[SWChisel.scala 171:41]
  wire  r_count_16_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_16_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_17_clock; // @[SWChisel.scala 171:41]
  wire  r_count_17_reset; // @[SWChisel.scala 171:41]
  wire  r_count_17_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_17_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_18_clock; // @[SWChisel.scala 171:41]
  wire  r_count_18_reset; // @[SWChisel.scala 171:41]
  wire  r_count_18_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_18_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_19_clock; // @[SWChisel.scala 171:41]
  wire  r_count_19_reset; // @[SWChisel.scala 171:41]
  wire  r_count_19_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_19_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_20_clock; // @[SWChisel.scala 171:41]
  wire  r_count_20_reset; // @[SWChisel.scala 171:41]
  wire  r_count_20_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_20_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_21_clock; // @[SWChisel.scala 171:41]
  wire  r_count_21_reset; // @[SWChisel.scala 171:41]
  wire  r_count_21_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_21_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_22_clock; // @[SWChisel.scala 171:41]
  wire  r_count_22_reset; // @[SWChisel.scala 171:41]
  wire  r_count_22_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_22_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_23_clock; // @[SWChisel.scala 171:41]
  wire  r_count_23_reset; // @[SWChisel.scala 171:41]
  wire  r_count_23_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_23_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_24_clock; // @[SWChisel.scala 171:41]
  wire  r_count_24_reset; // @[SWChisel.scala 171:41]
  wire  r_count_24_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_24_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_25_clock; // @[SWChisel.scala 171:41]
  wire  r_count_25_reset; // @[SWChisel.scala 171:41]
  wire  r_count_25_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_25_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_26_clock; // @[SWChisel.scala 171:41]
  wire  r_count_26_reset; // @[SWChisel.scala 171:41]
  wire  r_count_26_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_26_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_27_clock; // @[SWChisel.scala 171:41]
  wire  r_count_27_reset; // @[SWChisel.scala 171:41]
  wire  r_count_27_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_27_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_28_clock; // @[SWChisel.scala 171:41]
  wire  r_count_28_reset; // @[SWChisel.scala 171:41]
  wire  r_count_28_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_28_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_29_clock; // @[SWChisel.scala 171:41]
  wire  r_count_29_reset; // @[SWChisel.scala 171:41]
  wire  r_count_29_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_29_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_30_clock; // @[SWChisel.scala 171:41]
  wire  r_count_30_reset; // @[SWChisel.scala 171:41]
  wire  r_count_30_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_30_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_31_clock; // @[SWChisel.scala 171:41]
  wire  r_count_31_reset; // @[SWChisel.scala 171:41]
  wire  r_count_31_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_31_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_32_clock; // @[SWChisel.scala 171:41]
  wire  r_count_32_reset; // @[SWChisel.scala 171:41]
  wire  r_count_32_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_32_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_33_clock; // @[SWChisel.scala 171:41]
  wire  r_count_33_reset; // @[SWChisel.scala 171:41]
  wire  r_count_33_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_33_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_34_clock; // @[SWChisel.scala 171:41]
  wire  r_count_34_reset; // @[SWChisel.scala 171:41]
  wire  r_count_34_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_34_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_35_clock; // @[SWChisel.scala 171:41]
  wire  r_count_35_reset; // @[SWChisel.scala 171:41]
  wire  r_count_35_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_35_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_36_clock; // @[SWChisel.scala 171:41]
  wire  r_count_36_reset; // @[SWChisel.scala 171:41]
  wire  r_count_36_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_36_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_37_clock; // @[SWChisel.scala 171:41]
  wire  r_count_37_reset; // @[SWChisel.scala 171:41]
  wire  r_count_37_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_37_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_38_clock; // @[SWChisel.scala 171:41]
  wire  r_count_38_reset; // @[SWChisel.scala 171:41]
  wire  r_count_38_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_38_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_39_clock; // @[SWChisel.scala 171:41]
  wire  r_count_39_reset; // @[SWChisel.scala 171:41]
  wire  r_count_39_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_39_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_40_clock; // @[SWChisel.scala 171:41]
  wire  r_count_40_reset; // @[SWChisel.scala 171:41]
  wire  r_count_40_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_40_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_41_clock; // @[SWChisel.scala 171:41]
  wire  r_count_41_reset; // @[SWChisel.scala 171:41]
  wire  r_count_41_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_41_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_42_clock; // @[SWChisel.scala 171:41]
  wire  r_count_42_reset; // @[SWChisel.scala 171:41]
  wire  r_count_42_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_42_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_43_clock; // @[SWChisel.scala 171:41]
  wire  r_count_43_reset; // @[SWChisel.scala 171:41]
  wire  r_count_43_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_43_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_44_clock; // @[SWChisel.scala 171:41]
  wire  r_count_44_reset; // @[SWChisel.scala 171:41]
  wire  r_count_44_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_44_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_45_clock; // @[SWChisel.scala 171:41]
  wire  r_count_45_reset; // @[SWChisel.scala 171:41]
  wire  r_count_45_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_45_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_46_clock; // @[SWChisel.scala 171:41]
  wire  r_count_46_reset; // @[SWChisel.scala 171:41]
  wire  r_count_46_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_46_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_47_clock; // @[SWChisel.scala 171:41]
  wire  r_count_47_reset; // @[SWChisel.scala 171:41]
  wire  r_count_47_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_47_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_48_clock; // @[SWChisel.scala 171:41]
  wire  r_count_48_reset; // @[SWChisel.scala 171:41]
  wire  r_count_48_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_48_io_out; // @[SWChisel.scala 171:41]
  wire  r_count_49_clock; // @[SWChisel.scala 171:41]
  wire  r_count_49_reset; // @[SWChisel.scala 171:41]
  wire  r_count_49_io_en; // @[SWChisel.scala 171:41]
  wire [6:0] r_count_49_io_out; // @[SWChisel.scala 171:41]
  wire  max_clock; // @[SWChisel.scala 174:19]
  wire  max_reset; // @[SWChisel.scala 174:19]
  wire  max_io_start; // @[SWChisel.scala 174:19]
  wire [15:0] max_io_in; // @[SWChisel.scala 174:19]
  wire  max_io_done; // @[SWChisel.scala 174:19]
  wire [15:0] max_io_out; // @[SWChisel.scala 174:19]
  reg [15:0] E_0; // @[SWChisel.scala 162:18]
  reg [15:0] E_1; // @[SWChisel.scala 162:18]
  reg [15:0] E_2; // @[SWChisel.scala 162:18]
  reg [15:0] E_3; // @[SWChisel.scala 162:18]
  reg [15:0] E_4; // @[SWChisel.scala 162:18]
  reg [15:0] E_5; // @[SWChisel.scala 162:18]
  reg [15:0] E_6; // @[SWChisel.scala 162:18]
  reg [15:0] E_7; // @[SWChisel.scala 162:18]
  reg [15:0] E_8; // @[SWChisel.scala 162:18]
  reg [15:0] E_9; // @[SWChisel.scala 162:18]
  reg [15:0] E_10; // @[SWChisel.scala 162:18]
  reg [15:0] E_11; // @[SWChisel.scala 162:18]
  reg [15:0] E_12; // @[SWChisel.scala 162:18]
  reg [15:0] E_13; // @[SWChisel.scala 162:18]
  reg [15:0] E_14; // @[SWChisel.scala 162:18]
  reg [15:0] E_15; // @[SWChisel.scala 162:18]
  reg [15:0] E_16; // @[SWChisel.scala 162:18]
  reg [15:0] E_17; // @[SWChisel.scala 162:18]
  reg [15:0] E_18; // @[SWChisel.scala 162:18]
  reg [15:0] E_19; // @[SWChisel.scala 162:18]
  reg [15:0] E_20; // @[SWChisel.scala 162:18]
  reg [15:0] E_21; // @[SWChisel.scala 162:18]
  reg [15:0] E_22; // @[SWChisel.scala 162:18]
  reg [15:0] E_23; // @[SWChisel.scala 162:18]
  reg [15:0] E_24; // @[SWChisel.scala 162:18]
  reg [15:0] E_25; // @[SWChisel.scala 162:18]
  reg [15:0] E_26; // @[SWChisel.scala 162:18]
  reg [15:0] E_27; // @[SWChisel.scala 162:18]
  reg [15:0] E_28; // @[SWChisel.scala 162:18]
  reg [15:0] E_29; // @[SWChisel.scala 162:18]
  reg [15:0] E_30; // @[SWChisel.scala 162:18]
  reg [15:0] E_31; // @[SWChisel.scala 162:18]
  reg [15:0] E_32; // @[SWChisel.scala 162:18]
  reg [15:0] E_33; // @[SWChisel.scala 162:18]
  reg [15:0] E_34; // @[SWChisel.scala 162:18]
  reg [15:0] E_35; // @[SWChisel.scala 162:18]
  reg [15:0] E_36; // @[SWChisel.scala 162:18]
  reg [15:0] E_37; // @[SWChisel.scala 162:18]
  reg [15:0] E_38; // @[SWChisel.scala 162:18]
  reg [15:0] E_39; // @[SWChisel.scala 162:18]
  reg [15:0] E_40; // @[SWChisel.scala 162:18]
  reg [15:0] E_41; // @[SWChisel.scala 162:18]
  reg [15:0] E_42; // @[SWChisel.scala 162:18]
  reg [15:0] E_43; // @[SWChisel.scala 162:18]
  reg [15:0] E_44; // @[SWChisel.scala 162:18]
  reg [15:0] E_45; // @[SWChisel.scala 162:18]
  reg [15:0] E_46; // @[SWChisel.scala 162:18]
  reg [15:0] E_47; // @[SWChisel.scala 162:18]
  reg [15:0] E_48; // @[SWChisel.scala 162:18]
  reg [15:0] E_49; // @[SWChisel.scala 162:18]
  reg [15:0] F_1; // @[SWChisel.scala 163:18]
  reg [15:0] F_2; // @[SWChisel.scala 163:18]
  reg [15:0] F_3; // @[SWChisel.scala 163:18]
  reg [15:0] F_4; // @[SWChisel.scala 163:18]
  reg [15:0] F_5; // @[SWChisel.scala 163:18]
  reg [15:0] F_6; // @[SWChisel.scala 163:18]
  reg [15:0] F_7; // @[SWChisel.scala 163:18]
  reg [15:0] F_8; // @[SWChisel.scala 163:18]
  reg [15:0] F_9; // @[SWChisel.scala 163:18]
  reg [15:0] F_10; // @[SWChisel.scala 163:18]
  reg [15:0] F_11; // @[SWChisel.scala 163:18]
  reg [15:0] F_12; // @[SWChisel.scala 163:18]
  reg [15:0] F_13; // @[SWChisel.scala 163:18]
  reg [15:0] F_14; // @[SWChisel.scala 163:18]
  reg [15:0] F_15; // @[SWChisel.scala 163:18]
  reg [15:0] F_16; // @[SWChisel.scala 163:18]
  reg [15:0] F_17; // @[SWChisel.scala 163:18]
  reg [15:0] F_18; // @[SWChisel.scala 163:18]
  reg [15:0] F_19; // @[SWChisel.scala 163:18]
  reg [15:0] F_20; // @[SWChisel.scala 163:18]
  reg [15:0] F_21; // @[SWChisel.scala 163:18]
  reg [15:0] F_22; // @[SWChisel.scala 163:18]
  reg [15:0] F_23; // @[SWChisel.scala 163:18]
  reg [15:0] F_24; // @[SWChisel.scala 163:18]
  reg [15:0] F_25; // @[SWChisel.scala 163:18]
  reg [15:0] F_26; // @[SWChisel.scala 163:18]
  reg [15:0] F_27; // @[SWChisel.scala 163:18]
  reg [15:0] F_28; // @[SWChisel.scala 163:18]
  reg [15:0] F_29; // @[SWChisel.scala 163:18]
  reg [15:0] F_30; // @[SWChisel.scala 163:18]
  reg [15:0] F_31; // @[SWChisel.scala 163:18]
  reg [15:0] F_32; // @[SWChisel.scala 163:18]
  reg [15:0] F_33; // @[SWChisel.scala 163:18]
  reg [15:0] F_34; // @[SWChisel.scala 163:18]
  reg [15:0] F_35; // @[SWChisel.scala 163:18]
  reg [15:0] F_36; // @[SWChisel.scala 163:18]
  reg [15:0] F_37; // @[SWChisel.scala 163:18]
  reg [15:0] F_38; // @[SWChisel.scala 163:18]
  reg [15:0] F_39; // @[SWChisel.scala 163:18]
  reg [15:0] F_40; // @[SWChisel.scala 163:18]
  reg [15:0] F_41; // @[SWChisel.scala 163:18]
  reg [15:0] F_42; // @[SWChisel.scala 163:18]
  reg [15:0] F_43; // @[SWChisel.scala 163:18]
  reg [15:0] F_44; // @[SWChisel.scala 163:18]
  reg [15:0] F_45; // @[SWChisel.scala 163:18]
  reg [15:0] F_46; // @[SWChisel.scala 163:18]
  reg [15:0] F_47; // @[SWChisel.scala 163:18]
  reg [15:0] F_48; // @[SWChisel.scala 163:18]
  reg [15:0] F_49; // @[SWChisel.scala 163:18]
  reg [15:0] V1_0; // @[SWChisel.scala 164:19]
  reg [15:0] V1_1; // @[SWChisel.scala 164:19]
  reg [15:0] V1_2; // @[SWChisel.scala 164:19]
  reg [15:0] V1_3; // @[SWChisel.scala 164:19]
  reg [15:0] V1_4; // @[SWChisel.scala 164:19]
  reg [15:0] V1_5; // @[SWChisel.scala 164:19]
  reg [15:0] V1_6; // @[SWChisel.scala 164:19]
  reg [15:0] V1_7; // @[SWChisel.scala 164:19]
  reg [15:0] V1_8; // @[SWChisel.scala 164:19]
  reg [15:0] V1_9; // @[SWChisel.scala 164:19]
  reg [15:0] V1_10; // @[SWChisel.scala 164:19]
  reg [15:0] V1_11; // @[SWChisel.scala 164:19]
  reg [15:0] V1_12; // @[SWChisel.scala 164:19]
  reg [15:0] V1_13; // @[SWChisel.scala 164:19]
  reg [15:0] V1_14; // @[SWChisel.scala 164:19]
  reg [15:0] V1_15; // @[SWChisel.scala 164:19]
  reg [15:0] V1_16; // @[SWChisel.scala 164:19]
  reg [15:0] V1_17; // @[SWChisel.scala 164:19]
  reg [15:0] V1_18; // @[SWChisel.scala 164:19]
  reg [15:0] V1_19; // @[SWChisel.scala 164:19]
  reg [15:0] V1_20; // @[SWChisel.scala 164:19]
  reg [15:0] V1_21; // @[SWChisel.scala 164:19]
  reg [15:0] V1_22; // @[SWChisel.scala 164:19]
  reg [15:0] V1_23; // @[SWChisel.scala 164:19]
  reg [15:0] V1_24; // @[SWChisel.scala 164:19]
  reg [15:0] V1_25; // @[SWChisel.scala 164:19]
  reg [15:0] V1_26; // @[SWChisel.scala 164:19]
  reg [15:0] V1_27; // @[SWChisel.scala 164:19]
  reg [15:0] V1_28; // @[SWChisel.scala 164:19]
  reg [15:0] V1_29; // @[SWChisel.scala 164:19]
  reg [15:0] V1_30; // @[SWChisel.scala 164:19]
  reg [15:0] V1_31; // @[SWChisel.scala 164:19]
  reg [15:0] V1_32; // @[SWChisel.scala 164:19]
  reg [15:0] V1_33; // @[SWChisel.scala 164:19]
  reg [15:0] V1_34; // @[SWChisel.scala 164:19]
  reg [15:0] V1_35; // @[SWChisel.scala 164:19]
  reg [15:0] V1_36; // @[SWChisel.scala 164:19]
  reg [15:0] V1_37; // @[SWChisel.scala 164:19]
  reg [15:0] V1_38; // @[SWChisel.scala 164:19]
  reg [15:0] V1_39; // @[SWChisel.scala 164:19]
  reg [15:0] V1_40; // @[SWChisel.scala 164:19]
  reg [15:0] V1_41; // @[SWChisel.scala 164:19]
  reg [15:0] V1_42; // @[SWChisel.scala 164:19]
  reg [15:0] V1_43; // @[SWChisel.scala 164:19]
  reg [15:0] V1_44; // @[SWChisel.scala 164:19]
  reg [15:0] V1_45; // @[SWChisel.scala 164:19]
  reg [15:0] V1_46; // @[SWChisel.scala 164:19]
  reg [15:0] V1_47; // @[SWChisel.scala 164:19]
  reg [15:0] V1_48; // @[SWChisel.scala 164:19]
  reg [15:0] V1_49; // @[SWChisel.scala 164:19]
  reg [15:0] V1_50; // @[SWChisel.scala 164:19]
  reg [15:0] V2_0; // @[SWChisel.scala 166:19]
  reg [15:0] V2_1; // @[SWChisel.scala 166:19]
  reg [15:0] V2_2; // @[SWChisel.scala 166:19]
  reg [15:0] V2_3; // @[SWChisel.scala 166:19]
  reg [15:0] V2_4; // @[SWChisel.scala 166:19]
  reg [15:0] V2_5; // @[SWChisel.scala 166:19]
  reg [15:0] V2_6; // @[SWChisel.scala 166:19]
  reg [15:0] V2_7; // @[SWChisel.scala 166:19]
  reg [15:0] V2_8; // @[SWChisel.scala 166:19]
  reg [15:0] V2_9; // @[SWChisel.scala 166:19]
  reg [15:0] V2_10; // @[SWChisel.scala 166:19]
  reg [15:0] V2_11; // @[SWChisel.scala 166:19]
  reg [15:0] V2_12; // @[SWChisel.scala 166:19]
  reg [15:0] V2_13; // @[SWChisel.scala 166:19]
  reg [15:0] V2_14; // @[SWChisel.scala 166:19]
  reg [15:0] V2_15; // @[SWChisel.scala 166:19]
  reg [15:0] V2_16; // @[SWChisel.scala 166:19]
  reg [15:0] V2_17; // @[SWChisel.scala 166:19]
  reg [15:0] V2_18; // @[SWChisel.scala 166:19]
  reg [15:0] V2_19; // @[SWChisel.scala 166:19]
  reg [15:0] V2_20; // @[SWChisel.scala 166:19]
  reg [15:0] V2_21; // @[SWChisel.scala 166:19]
  reg [15:0] V2_22; // @[SWChisel.scala 166:19]
  reg [15:0] V2_23; // @[SWChisel.scala 166:19]
  reg [15:0] V2_24; // @[SWChisel.scala 166:19]
  reg [15:0] V2_25; // @[SWChisel.scala 166:19]
  reg [15:0] V2_26; // @[SWChisel.scala 166:19]
  reg [15:0] V2_27; // @[SWChisel.scala 166:19]
  reg [15:0] V2_28; // @[SWChisel.scala 166:19]
  reg [15:0] V2_29; // @[SWChisel.scala 166:19]
  reg [15:0] V2_30; // @[SWChisel.scala 166:19]
  reg [15:0] V2_31; // @[SWChisel.scala 166:19]
  reg [15:0] V2_32; // @[SWChisel.scala 166:19]
  reg [15:0] V2_33; // @[SWChisel.scala 166:19]
  reg [15:0] V2_34; // @[SWChisel.scala 166:19]
  reg [15:0] V2_35; // @[SWChisel.scala 166:19]
  reg [15:0] V2_36; // @[SWChisel.scala 166:19]
  reg [15:0] V2_37; // @[SWChisel.scala 166:19]
  reg [15:0] V2_38; // @[SWChisel.scala 166:19]
  reg [15:0] V2_39; // @[SWChisel.scala 166:19]
  reg [15:0] V2_40; // @[SWChisel.scala 166:19]
  reg [15:0] V2_41; // @[SWChisel.scala 166:19]
  reg [15:0] V2_42; // @[SWChisel.scala 166:19]
  reg [15:0] V2_43; // @[SWChisel.scala 166:19]
  reg [15:0] V2_44; // @[SWChisel.scala 166:19]
  reg [15:0] V2_45; // @[SWChisel.scala 166:19]
  reg [15:0] V2_46; // @[SWChisel.scala 166:19]
  reg [15:0] V2_47; // @[SWChisel.scala 166:19]
  reg [15:0] V2_48; // @[SWChisel.scala 166:19]
  reg [15:0] V2_49; // @[SWChisel.scala 166:19]
  reg  start_reg_0; // @[SWChisel.scala 167:26]
  reg  start_reg_1; // @[SWChisel.scala 167:26]
  reg  start_reg_2; // @[SWChisel.scala 167:26]
  reg  start_reg_3; // @[SWChisel.scala 167:26]
  reg  start_reg_4; // @[SWChisel.scala 167:26]
  reg  start_reg_5; // @[SWChisel.scala 167:26]
  reg  start_reg_6; // @[SWChisel.scala 167:26]
  reg  start_reg_7; // @[SWChisel.scala 167:26]
  reg  start_reg_8; // @[SWChisel.scala 167:26]
  reg  start_reg_9; // @[SWChisel.scala 167:26]
  reg  start_reg_10; // @[SWChisel.scala 167:26]
  reg  start_reg_11; // @[SWChisel.scala 167:26]
  reg  start_reg_12; // @[SWChisel.scala 167:26]
  reg  start_reg_13; // @[SWChisel.scala 167:26]
  reg  start_reg_14; // @[SWChisel.scala 167:26]
  reg  start_reg_15; // @[SWChisel.scala 167:26]
  reg  start_reg_16; // @[SWChisel.scala 167:26]
  reg  start_reg_17; // @[SWChisel.scala 167:26]
  reg  start_reg_18; // @[SWChisel.scala 167:26]
  reg  start_reg_19; // @[SWChisel.scala 167:26]
  reg  start_reg_20; // @[SWChisel.scala 167:26]
  reg  start_reg_21; // @[SWChisel.scala 167:26]
  reg  start_reg_22; // @[SWChisel.scala 167:26]
  reg  start_reg_23; // @[SWChisel.scala 167:26]
  reg  start_reg_24; // @[SWChisel.scala 167:26]
  reg  start_reg_25; // @[SWChisel.scala 167:26]
  reg  start_reg_26; // @[SWChisel.scala 167:26]
  reg  start_reg_27; // @[SWChisel.scala 167:26]
  reg  start_reg_28; // @[SWChisel.scala 167:26]
  reg  start_reg_29; // @[SWChisel.scala 167:26]
  reg  start_reg_30; // @[SWChisel.scala 167:26]
  reg  start_reg_31; // @[SWChisel.scala 167:26]
  reg  start_reg_32; // @[SWChisel.scala 167:26]
  reg  start_reg_33; // @[SWChisel.scala 167:26]
  reg  start_reg_34; // @[SWChisel.scala 167:26]
  reg  start_reg_35; // @[SWChisel.scala 167:26]
  reg  start_reg_36; // @[SWChisel.scala 167:26]
  reg  start_reg_37; // @[SWChisel.scala 167:26]
  reg  start_reg_38; // @[SWChisel.scala 167:26]
  reg  start_reg_39; // @[SWChisel.scala 167:26]
  reg  start_reg_40; // @[SWChisel.scala 167:26]
  reg  start_reg_41; // @[SWChisel.scala 167:26]
  reg  start_reg_42; // @[SWChisel.scala 167:26]
  reg  start_reg_43; // @[SWChisel.scala 167:26]
  reg  start_reg_44; // @[SWChisel.scala 167:26]
  reg  start_reg_45; // @[SWChisel.scala 167:26]
  reg  start_reg_46; // @[SWChisel.scala 167:26]
  reg  start_reg_47; // @[SWChisel.scala 167:26]
  reg  start_reg_48; // @[SWChisel.scala 167:26]
  reg  start_reg_49; // @[SWChisel.scala 167:26]
  wire [1:0] _GEN_151 = 7'h1 == r_count_0_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_152 = 7'h2 == r_count_0_io_out ? io_r_2_b : _GEN_151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_153 = 7'h3 == r_count_0_io_out ? io_r_3_b : _GEN_152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_154 = 7'h4 == r_count_0_io_out ? io_r_4_b : _GEN_153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_155 = 7'h5 == r_count_0_io_out ? io_r_5_b : _GEN_154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_156 = 7'h6 == r_count_0_io_out ? io_r_6_b : _GEN_155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_157 = 7'h7 == r_count_0_io_out ? io_r_7_b : _GEN_156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_158 = 7'h8 == r_count_0_io_out ? io_r_8_b : _GEN_157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_159 = 7'h9 == r_count_0_io_out ? io_r_9_b : _GEN_158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_160 = 7'ha == r_count_0_io_out ? io_r_10_b : _GEN_159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_161 = 7'hb == r_count_0_io_out ? io_r_11_b : _GEN_160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_162 = 7'hc == r_count_0_io_out ? io_r_12_b : _GEN_161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_163 = 7'hd == r_count_0_io_out ? io_r_13_b : _GEN_162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_164 = 7'he == r_count_0_io_out ? io_r_14_b : _GEN_163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_165 = 7'hf == r_count_0_io_out ? io_r_15_b : _GEN_164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_166 = 7'h10 == r_count_0_io_out ? io_r_16_b : _GEN_165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_167 = 7'h11 == r_count_0_io_out ? io_r_17_b : _GEN_166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_168 = 7'h12 == r_count_0_io_out ? io_r_18_b : _GEN_167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_169 = 7'h13 == r_count_0_io_out ? io_r_19_b : _GEN_168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_170 = 7'h14 == r_count_0_io_out ? io_r_20_b : _GEN_169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_171 = 7'h15 == r_count_0_io_out ? io_r_21_b : _GEN_170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_172 = 7'h16 == r_count_0_io_out ? io_r_22_b : _GEN_171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_173 = 7'h17 == r_count_0_io_out ? io_r_23_b : _GEN_172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_174 = 7'h18 == r_count_0_io_out ? io_r_24_b : _GEN_173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_175 = 7'h19 == r_count_0_io_out ? io_r_25_b : _GEN_174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_176 = 7'h1a == r_count_0_io_out ? io_r_26_b : _GEN_175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_177 = 7'h1b == r_count_0_io_out ? io_r_27_b : _GEN_176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_178 = 7'h1c == r_count_0_io_out ? io_r_28_b : _GEN_177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_179 = 7'h1d == r_count_0_io_out ? io_r_29_b : _GEN_178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_180 = 7'h1e == r_count_0_io_out ? io_r_30_b : _GEN_179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_181 = 7'h1f == r_count_0_io_out ? io_r_31_b : _GEN_180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_182 = 7'h20 == r_count_0_io_out ? io_r_32_b : _GEN_181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_183 = 7'h21 == r_count_0_io_out ? io_r_33_b : _GEN_182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_184 = 7'h22 == r_count_0_io_out ? io_r_34_b : _GEN_183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_185 = 7'h23 == r_count_0_io_out ? io_r_35_b : _GEN_184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_186 = 7'h24 == r_count_0_io_out ? io_r_36_b : _GEN_185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_187 = 7'h25 == r_count_0_io_out ? io_r_37_b : _GEN_186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_188 = 7'h26 == r_count_0_io_out ? io_r_38_b : _GEN_187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_189 = 7'h27 == r_count_0_io_out ? io_r_39_b : _GEN_188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_190 = 7'h28 == r_count_0_io_out ? io_r_40_b : _GEN_189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_191 = 7'h29 == r_count_0_io_out ? io_r_41_b : _GEN_190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_192 = 7'h2a == r_count_0_io_out ? io_r_42_b : _GEN_191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_193 = 7'h2b == r_count_0_io_out ? io_r_43_b : _GEN_192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_194 = 7'h2c == r_count_0_io_out ? io_r_44_b : _GEN_193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_195 = 7'h2d == r_count_0_io_out ? io_r_45_b : _GEN_194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_196 = 7'h2e == r_count_0_io_out ? io_r_46_b : _GEN_195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_197 = 7'h2f == r_count_0_io_out ? io_r_47_b : _GEN_196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_198 = 7'h30 == r_count_0_io_out ? io_r_48_b : _GEN_197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_199 = 7'h31 == r_count_0_io_out ? io_r_49_b : _GEN_198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_200 = 7'h32 == r_count_0_io_out ? io_r_50_b : _GEN_199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_201 = 7'h33 == r_count_0_io_out ? io_r_51_b : _GEN_200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_202 = 7'h34 == r_count_0_io_out ? io_r_52_b : _GEN_201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_203 = 7'h35 == r_count_0_io_out ? io_r_53_b : _GEN_202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_204 = 7'h36 == r_count_0_io_out ? io_r_54_b : _GEN_203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_205 = 7'h37 == r_count_0_io_out ? io_r_55_b : _GEN_204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_206 = 7'h38 == r_count_0_io_out ? io_r_56_b : _GEN_205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_207 = 7'h39 == r_count_0_io_out ? io_r_57_b : _GEN_206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_208 = 7'h3a == r_count_0_io_out ? io_r_58_b : _GEN_207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_209 = 7'h3b == r_count_0_io_out ? io_r_59_b : _GEN_208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_210 = 7'h3c == r_count_0_io_out ? io_r_60_b : _GEN_209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_211 = 7'h3d == r_count_0_io_out ? io_r_61_b : _GEN_210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_212 = 7'h3e == r_count_0_io_out ? io_r_62_b : _GEN_211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_213 = 7'h3f == r_count_0_io_out ? io_r_63_b : _GEN_212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_214 = 7'h40 == r_count_0_io_out ? io_r_64_b : _GEN_213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_215 = 7'h41 == r_count_0_io_out ? io_r_65_b : _GEN_214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_216 = 7'h42 == r_count_0_io_out ? io_r_66_b : _GEN_215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_217 = 7'h43 == r_count_0_io_out ? io_r_67_b : _GEN_216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_218 = 7'h44 == r_count_0_io_out ? io_r_68_b : _GEN_217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_219 = 7'h45 == r_count_0_io_out ? io_r_69_b : _GEN_218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_220 = 7'h46 == r_count_0_io_out ? io_r_70_b : _GEN_219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_221 = 7'h47 == r_count_0_io_out ? io_r_71_b : _GEN_220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_222 = 7'h48 == r_count_0_io_out ? io_r_72_b : _GEN_221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_223 = 7'h49 == r_count_0_io_out ? io_r_73_b : _GEN_222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_224 = 7'h4a == r_count_0_io_out ? io_r_74_b : _GEN_223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_225 = 7'h4b == r_count_0_io_out ? io_r_75_b : _GEN_224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_226 = 7'h4c == r_count_0_io_out ? io_r_76_b : _GEN_225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_227 = 7'h4d == r_count_0_io_out ? io_r_77_b : _GEN_226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_228 = 7'h4e == r_count_0_io_out ? io_r_78_b : _GEN_227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_229 = 7'h4f == r_count_0_io_out ? io_r_79_b : _GEN_228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_230 = 7'h50 == r_count_0_io_out ? io_r_80_b : _GEN_229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_231 = 7'h51 == r_count_0_io_out ? io_r_81_b : _GEN_230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_232 = 7'h52 == r_count_0_io_out ? io_r_82_b : _GEN_231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_233 = 7'h53 == r_count_0_io_out ? io_r_83_b : _GEN_232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_234 = 7'h54 == r_count_0_io_out ? io_r_84_b : _GEN_233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_235 = 7'h55 == r_count_0_io_out ? io_r_85_b : _GEN_234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_236 = 7'h56 == r_count_0_io_out ? io_r_86_b : _GEN_235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_237 = 7'h57 == r_count_0_io_out ? io_r_87_b : _GEN_236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_238 = 7'h58 == r_count_0_io_out ? io_r_88_b : _GEN_237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_239 = 7'h59 == r_count_0_io_out ? io_r_89_b : _GEN_238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_240 = 7'h5a == r_count_0_io_out ? io_r_90_b : _GEN_239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_241 = 7'h5b == r_count_0_io_out ? io_r_91_b : _GEN_240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_242 = 7'h5c == r_count_0_io_out ? io_r_92_b : _GEN_241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_243 = 7'h5d == r_count_0_io_out ? io_r_93_b : _GEN_242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_244 = 7'h5e == r_count_0_io_out ? io_r_94_b : _GEN_243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_245 = 7'h5f == r_count_0_io_out ? io_r_95_b : _GEN_244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_246 = 7'h60 == r_count_0_io_out ? io_r_96_b : _GEN_245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_247 = 7'h61 == r_count_0_io_out ? io_r_97_b : _GEN_246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_248 = 7'h62 == r_count_0_io_out ? io_r_98_b : _GEN_247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_251 = 7'h1 == r_count_1_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_252 = 7'h2 == r_count_1_io_out ? io_r_2_b : _GEN_251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_253 = 7'h3 == r_count_1_io_out ? io_r_3_b : _GEN_252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_254 = 7'h4 == r_count_1_io_out ? io_r_4_b : _GEN_253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_255 = 7'h5 == r_count_1_io_out ? io_r_5_b : _GEN_254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_256 = 7'h6 == r_count_1_io_out ? io_r_6_b : _GEN_255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_257 = 7'h7 == r_count_1_io_out ? io_r_7_b : _GEN_256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_258 = 7'h8 == r_count_1_io_out ? io_r_8_b : _GEN_257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_259 = 7'h9 == r_count_1_io_out ? io_r_9_b : _GEN_258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_260 = 7'ha == r_count_1_io_out ? io_r_10_b : _GEN_259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_261 = 7'hb == r_count_1_io_out ? io_r_11_b : _GEN_260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_262 = 7'hc == r_count_1_io_out ? io_r_12_b : _GEN_261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_263 = 7'hd == r_count_1_io_out ? io_r_13_b : _GEN_262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_264 = 7'he == r_count_1_io_out ? io_r_14_b : _GEN_263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_265 = 7'hf == r_count_1_io_out ? io_r_15_b : _GEN_264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_266 = 7'h10 == r_count_1_io_out ? io_r_16_b : _GEN_265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_267 = 7'h11 == r_count_1_io_out ? io_r_17_b : _GEN_266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_268 = 7'h12 == r_count_1_io_out ? io_r_18_b : _GEN_267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_269 = 7'h13 == r_count_1_io_out ? io_r_19_b : _GEN_268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_270 = 7'h14 == r_count_1_io_out ? io_r_20_b : _GEN_269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_271 = 7'h15 == r_count_1_io_out ? io_r_21_b : _GEN_270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_272 = 7'h16 == r_count_1_io_out ? io_r_22_b : _GEN_271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_273 = 7'h17 == r_count_1_io_out ? io_r_23_b : _GEN_272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_274 = 7'h18 == r_count_1_io_out ? io_r_24_b : _GEN_273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_275 = 7'h19 == r_count_1_io_out ? io_r_25_b : _GEN_274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_276 = 7'h1a == r_count_1_io_out ? io_r_26_b : _GEN_275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_277 = 7'h1b == r_count_1_io_out ? io_r_27_b : _GEN_276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_278 = 7'h1c == r_count_1_io_out ? io_r_28_b : _GEN_277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_279 = 7'h1d == r_count_1_io_out ? io_r_29_b : _GEN_278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_280 = 7'h1e == r_count_1_io_out ? io_r_30_b : _GEN_279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_281 = 7'h1f == r_count_1_io_out ? io_r_31_b : _GEN_280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_282 = 7'h20 == r_count_1_io_out ? io_r_32_b : _GEN_281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_283 = 7'h21 == r_count_1_io_out ? io_r_33_b : _GEN_282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_284 = 7'h22 == r_count_1_io_out ? io_r_34_b : _GEN_283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_285 = 7'h23 == r_count_1_io_out ? io_r_35_b : _GEN_284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_286 = 7'h24 == r_count_1_io_out ? io_r_36_b : _GEN_285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_287 = 7'h25 == r_count_1_io_out ? io_r_37_b : _GEN_286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_288 = 7'h26 == r_count_1_io_out ? io_r_38_b : _GEN_287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_289 = 7'h27 == r_count_1_io_out ? io_r_39_b : _GEN_288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_290 = 7'h28 == r_count_1_io_out ? io_r_40_b : _GEN_289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_291 = 7'h29 == r_count_1_io_out ? io_r_41_b : _GEN_290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_292 = 7'h2a == r_count_1_io_out ? io_r_42_b : _GEN_291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_293 = 7'h2b == r_count_1_io_out ? io_r_43_b : _GEN_292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_294 = 7'h2c == r_count_1_io_out ? io_r_44_b : _GEN_293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_295 = 7'h2d == r_count_1_io_out ? io_r_45_b : _GEN_294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_296 = 7'h2e == r_count_1_io_out ? io_r_46_b : _GEN_295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_297 = 7'h2f == r_count_1_io_out ? io_r_47_b : _GEN_296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_298 = 7'h30 == r_count_1_io_out ? io_r_48_b : _GEN_297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_299 = 7'h31 == r_count_1_io_out ? io_r_49_b : _GEN_298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_300 = 7'h32 == r_count_1_io_out ? io_r_50_b : _GEN_299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_301 = 7'h33 == r_count_1_io_out ? io_r_51_b : _GEN_300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_302 = 7'h34 == r_count_1_io_out ? io_r_52_b : _GEN_301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_303 = 7'h35 == r_count_1_io_out ? io_r_53_b : _GEN_302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_304 = 7'h36 == r_count_1_io_out ? io_r_54_b : _GEN_303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_305 = 7'h37 == r_count_1_io_out ? io_r_55_b : _GEN_304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_306 = 7'h38 == r_count_1_io_out ? io_r_56_b : _GEN_305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_307 = 7'h39 == r_count_1_io_out ? io_r_57_b : _GEN_306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_308 = 7'h3a == r_count_1_io_out ? io_r_58_b : _GEN_307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_309 = 7'h3b == r_count_1_io_out ? io_r_59_b : _GEN_308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_310 = 7'h3c == r_count_1_io_out ? io_r_60_b : _GEN_309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_311 = 7'h3d == r_count_1_io_out ? io_r_61_b : _GEN_310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_312 = 7'h3e == r_count_1_io_out ? io_r_62_b : _GEN_311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_313 = 7'h3f == r_count_1_io_out ? io_r_63_b : _GEN_312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_314 = 7'h40 == r_count_1_io_out ? io_r_64_b : _GEN_313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_315 = 7'h41 == r_count_1_io_out ? io_r_65_b : _GEN_314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_316 = 7'h42 == r_count_1_io_out ? io_r_66_b : _GEN_315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_317 = 7'h43 == r_count_1_io_out ? io_r_67_b : _GEN_316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_318 = 7'h44 == r_count_1_io_out ? io_r_68_b : _GEN_317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_319 = 7'h45 == r_count_1_io_out ? io_r_69_b : _GEN_318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_320 = 7'h46 == r_count_1_io_out ? io_r_70_b : _GEN_319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_321 = 7'h47 == r_count_1_io_out ? io_r_71_b : _GEN_320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_322 = 7'h48 == r_count_1_io_out ? io_r_72_b : _GEN_321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_323 = 7'h49 == r_count_1_io_out ? io_r_73_b : _GEN_322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_324 = 7'h4a == r_count_1_io_out ? io_r_74_b : _GEN_323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_325 = 7'h4b == r_count_1_io_out ? io_r_75_b : _GEN_324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_326 = 7'h4c == r_count_1_io_out ? io_r_76_b : _GEN_325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_327 = 7'h4d == r_count_1_io_out ? io_r_77_b : _GEN_326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_328 = 7'h4e == r_count_1_io_out ? io_r_78_b : _GEN_327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_329 = 7'h4f == r_count_1_io_out ? io_r_79_b : _GEN_328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_330 = 7'h50 == r_count_1_io_out ? io_r_80_b : _GEN_329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_331 = 7'h51 == r_count_1_io_out ? io_r_81_b : _GEN_330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_332 = 7'h52 == r_count_1_io_out ? io_r_82_b : _GEN_331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_333 = 7'h53 == r_count_1_io_out ? io_r_83_b : _GEN_332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_334 = 7'h54 == r_count_1_io_out ? io_r_84_b : _GEN_333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_335 = 7'h55 == r_count_1_io_out ? io_r_85_b : _GEN_334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_336 = 7'h56 == r_count_1_io_out ? io_r_86_b : _GEN_335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_337 = 7'h57 == r_count_1_io_out ? io_r_87_b : _GEN_336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_338 = 7'h58 == r_count_1_io_out ? io_r_88_b : _GEN_337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_339 = 7'h59 == r_count_1_io_out ? io_r_89_b : _GEN_338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_340 = 7'h5a == r_count_1_io_out ? io_r_90_b : _GEN_339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_341 = 7'h5b == r_count_1_io_out ? io_r_91_b : _GEN_340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_342 = 7'h5c == r_count_1_io_out ? io_r_92_b : _GEN_341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_343 = 7'h5d == r_count_1_io_out ? io_r_93_b : _GEN_342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_344 = 7'h5e == r_count_1_io_out ? io_r_94_b : _GEN_343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_345 = 7'h5f == r_count_1_io_out ? io_r_95_b : _GEN_344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_346 = 7'h60 == r_count_1_io_out ? io_r_96_b : _GEN_345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_347 = 7'h61 == r_count_1_io_out ? io_r_97_b : _GEN_346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_348 = 7'h62 == r_count_1_io_out ? io_r_98_b : _GEN_347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_351 = 7'h1 == r_count_2_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_352 = 7'h2 == r_count_2_io_out ? io_r_2_b : _GEN_351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_353 = 7'h3 == r_count_2_io_out ? io_r_3_b : _GEN_352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_354 = 7'h4 == r_count_2_io_out ? io_r_4_b : _GEN_353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_355 = 7'h5 == r_count_2_io_out ? io_r_5_b : _GEN_354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_356 = 7'h6 == r_count_2_io_out ? io_r_6_b : _GEN_355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_357 = 7'h7 == r_count_2_io_out ? io_r_7_b : _GEN_356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_358 = 7'h8 == r_count_2_io_out ? io_r_8_b : _GEN_357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_359 = 7'h9 == r_count_2_io_out ? io_r_9_b : _GEN_358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_360 = 7'ha == r_count_2_io_out ? io_r_10_b : _GEN_359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_361 = 7'hb == r_count_2_io_out ? io_r_11_b : _GEN_360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_362 = 7'hc == r_count_2_io_out ? io_r_12_b : _GEN_361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_363 = 7'hd == r_count_2_io_out ? io_r_13_b : _GEN_362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_364 = 7'he == r_count_2_io_out ? io_r_14_b : _GEN_363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_365 = 7'hf == r_count_2_io_out ? io_r_15_b : _GEN_364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_366 = 7'h10 == r_count_2_io_out ? io_r_16_b : _GEN_365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_367 = 7'h11 == r_count_2_io_out ? io_r_17_b : _GEN_366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_368 = 7'h12 == r_count_2_io_out ? io_r_18_b : _GEN_367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_369 = 7'h13 == r_count_2_io_out ? io_r_19_b : _GEN_368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_370 = 7'h14 == r_count_2_io_out ? io_r_20_b : _GEN_369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_371 = 7'h15 == r_count_2_io_out ? io_r_21_b : _GEN_370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_372 = 7'h16 == r_count_2_io_out ? io_r_22_b : _GEN_371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_373 = 7'h17 == r_count_2_io_out ? io_r_23_b : _GEN_372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_374 = 7'h18 == r_count_2_io_out ? io_r_24_b : _GEN_373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_375 = 7'h19 == r_count_2_io_out ? io_r_25_b : _GEN_374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_376 = 7'h1a == r_count_2_io_out ? io_r_26_b : _GEN_375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_377 = 7'h1b == r_count_2_io_out ? io_r_27_b : _GEN_376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_378 = 7'h1c == r_count_2_io_out ? io_r_28_b : _GEN_377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_379 = 7'h1d == r_count_2_io_out ? io_r_29_b : _GEN_378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_380 = 7'h1e == r_count_2_io_out ? io_r_30_b : _GEN_379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_381 = 7'h1f == r_count_2_io_out ? io_r_31_b : _GEN_380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_382 = 7'h20 == r_count_2_io_out ? io_r_32_b : _GEN_381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_383 = 7'h21 == r_count_2_io_out ? io_r_33_b : _GEN_382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_384 = 7'h22 == r_count_2_io_out ? io_r_34_b : _GEN_383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_385 = 7'h23 == r_count_2_io_out ? io_r_35_b : _GEN_384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_386 = 7'h24 == r_count_2_io_out ? io_r_36_b : _GEN_385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_387 = 7'h25 == r_count_2_io_out ? io_r_37_b : _GEN_386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_388 = 7'h26 == r_count_2_io_out ? io_r_38_b : _GEN_387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_389 = 7'h27 == r_count_2_io_out ? io_r_39_b : _GEN_388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_390 = 7'h28 == r_count_2_io_out ? io_r_40_b : _GEN_389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_391 = 7'h29 == r_count_2_io_out ? io_r_41_b : _GEN_390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_392 = 7'h2a == r_count_2_io_out ? io_r_42_b : _GEN_391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_393 = 7'h2b == r_count_2_io_out ? io_r_43_b : _GEN_392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_394 = 7'h2c == r_count_2_io_out ? io_r_44_b : _GEN_393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_395 = 7'h2d == r_count_2_io_out ? io_r_45_b : _GEN_394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_396 = 7'h2e == r_count_2_io_out ? io_r_46_b : _GEN_395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_397 = 7'h2f == r_count_2_io_out ? io_r_47_b : _GEN_396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_398 = 7'h30 == r_count_2_io_out ? io_r_48_b : _GEN_397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_399 = 7'h31 == r_count_2_io_out ? io_r_49_b : _GEN_398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_400 = 7'h32 == r_count_2_io_out ? io_r_50_b : _GEN_399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_401 = 7'h33 == r_count_2_io_out ? io_r_51_b : _GEN_400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_402 = 7'h34 == r_count_2_io_out ? io_r_52_b : _GEN_401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_403 = 7'h35 == r_count_2_io_out ? io_r_53_b : _GEN_402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_404 = 7'h36 == r_count_2_io_out ? io_r_54_b : _GEN_403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_405 = 7'h37 == r_count_2_io_out ? io_r_55_b : _GEN_404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_406 = 7'h38 == r_count_2_io_out ? io_r_56_b : _GEN_405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_407 = 7'h39 == r_count_2_io_out ? io_r_57_b : _GEN_406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_408 = 7'h3a == r_count_2_io_out ? io_r_58_b : _GEN_407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_409 = 7'h3b == r_count_2_io_out ? io_r_59_b : _GEN_408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_410 = 7'h3c == r_count_2_io_out ? io_r_60_b : _GEN_409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_411 = 7'h3d == r_count_2_io_out ? io_r_61_b : _GEN_410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_412 = 7'h3e == r_count_2_io_out ? io_r_62_b : _GEN_411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_413 = 7'h3f == r_count_2_io_out ? io_r_63_b : _GEN_412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_414 = 7'h40 == r_count_2_io_out ? io_r_64_b : _GEN_413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_415 = 7'h41 == r_count_2_io_out ? io_r_65_b : _GEN_414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_416 = 7'h42 == r_count_2_io_out ? io_r_66_b : _GEN_415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_417 = 7'h43 == r_count_2_io_out ? io_r_67_b : _GEN_416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_418 = 7'h44 == r_count_2_io_out ? io_r_68_b : _GEN_417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_419 = 7'h45 == r_count_2_io_out ? io_r_69_b : _GEN_418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_420 = 7'h46 == r_count_2_io_out ? io_r_70_b : _GEN_419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_421 = 7'h47 == r_count_2_io_out ? io_r_71_b : _GEN_420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_422 = 7'h48 == r_count_2_io_out ? io_r_72_b : _GEN_421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_423 = 7'h49 == r_count_2_io_out ? io_r_73_b : _GEN_422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_424 = 7'h4a == r_count_2_io_out ? io_r_74_b : _GEN_423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_425 = 7'h4b == r_count_2_io_out ? io_r_75_b : _GEN_424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_426 = 7'h4c == r_count_2_io_out ? io_r_76_b : _GEN_425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_427 = 7'h4d == r_count_2_io_out ? io_r_77_b : _GEN_426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_428 = 7'h4e == r_count_2_io_out ? io_r_78_b : _GEN_427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_429 = 7'h4f == r_count_2_io_out ? io_r_79_b : _GEN_428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_430 = 7'h50 == r_count_2_io_out ? io_r_80_b : _GEN_429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_431 = 7'h51 == r_count_2_io_out ? io_r_81_b : _GEN_430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_432 = 7'h52 == r_count_2_io_out ? io_r_82_b : _GEN_431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_433 = 7'h53 == r_count_2_io_out ? io_r_83_b : _GEN_432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_434 = 7'h54 == r_count_2_io_out ? io_r_84_b : _GEN_433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_435 = 7'h55 == r_count_2_io_out ? io_r_85_b : _GEN_434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_436 = 7'h56 == r_count_2_io_out ? io_r_86_b : _GEN_435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_437 = 7'h57 == r_count_2_io_out ? io_r_87_b : _GEN_436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_438 = 7'h58 == r_count_2_io_out ? io_r_88_b : _GEN_437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_439 = 7'h59 == r_count_2_io_out ? io_r_89_b : _GEN_438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_440 = 7'h5a == r_count_2_io_out ? io_r_90_b : _GEN_439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_441 = 7'h5b == r_count_2_io_out ? io_r_91_b : _GEN_440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_442 = 7'h5c == r_count_2_io_out ? io_r_92_b : _GEN_441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_443 = 7'h5d == r_count_2_io_out ? io_r_93_b : _GEN_442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_444 = 7'h5e == r_count_2_io_out ? io_r_94_b : _GEN_443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_445 = 7'h5f == r_count_2_io_out ? io_r_95_b : _GEN_444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_446 = 7'h60 == r_count_2_io_out ? io_r_96_b : _GEN_445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_447 = 7'h61 == r_count_2_io_out ? io_r_97_b : _GEN_446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_448 = 7'h62 == r_count_2_io_out ? io_r_98_b : _GEN_447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_451 = 7'h1 == r_count_3_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_452 = 7'h2 == r_count_3_io_out ? io_r_2_b : _GEN_451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_453 = 7'h3 == r_count_3_io_out ? io_r_3_b : _GEN_452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_454 = 7'h4 == r_count_3_io_out ? io_r_4_b : _GEN_453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_455 = 7'h5 == r_count_3_io_out ? io_r_5_b : _GEN_454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_456 = 7'h6 == r_count_3_io_out ? io_r_6_b : _GEN_455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_457 = 7'h7 == r_count_3_io_out ? io_r_7_b : _GEN_456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_458 = 7'h8 == r_count_3_io_out ? io_r_8_b : _GEN_457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_459 = 7'h9 == r_count_3_io_out ? io_r_9_b : _GEN_458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_460 = 7'ha == r_count_3_io_out ? io_r_10_b : _GEN_459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_461 = 7'hb == r_count_3_io_out ? io_r_11_b : _GEN_460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_462 = 7'hc == r_count_3_io_out ? io_r_12_b : _GEN_461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_463 = 7'hd == r_count_3_io_out ? io_r_13_b : _GEN_462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_464 = 7'he == r_count_3_io_out ? io_r_14_b : _GEN_463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_465 = 7'hf == r_count_3_io_out ? io_r_15_b : _GEN_464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_466 = 7'h10 == r_count_3_io_out ? io_r_16_b : _GEN_465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_467 = 7'h11 == r_count_3_io_out ? io_r_17_b : _GEN_466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_468 = 7'h12 == r_count_3_io_out ? io_r_18_b : _GEN_467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_469 = 7'h13 == r_count_3_io_out ? io_r_19_b : _GEN_468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_470 = 7'h14 == r_count_3_io_out ? io_r_20_b : _GEN_469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_471 = 7'h15 == r_count_3_io_out ? io_r_21_b : _GEN_470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_472 = 7'h16 == r_count_3_io_out ? io_r_22_b : _GEN_471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_473 = 7'h17 == r_count_3_io_out ? io_r_23_b : _GEN_472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_474 = 7'h18 == r_count_3_io_out ? io_r_24_b : _GEN_473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_475 = 7'h19 == r_count_3_io_out ? io_r_25_b : _GEN_474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_476 = 7'h1a == r_count_3_io_out ? io_r_26_b : _GEN_475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_477 = 7'h1b == r_count_3_io_out ? io_r_27_b : _GEN_476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_478 = 7'h1c == r_count_3_io_out ? io_r_28_b : _GEN_477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_479 = 7'h1d == r_count_3_io_out ? io_r_29_b : _GEN_478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_480 = 7'h1e == r_count_3_io_out ? io_r_30_b : _GEN_479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_481 = 7'h1f == r_count_3_io_out ? io_r_31_b : _GEN_480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_482 = 7'h20 == r_count_3_io_out ? io_r_32_b : _GEN_481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_483 = 7'h21 == r_count_3_io_out ? io_r_33_b : _GEN_482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_484 = 7'h22 == r_count_3_io_out ? io_r_34_b : _GEN_483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_485 = 7'h23 == r_count_3_io_out ? io_r_35_b : _GEN_484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_486 = 7'h24 == r_count_3_io_out ? io_r_36_b : _GEN_485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_487 = 7'h25 == r_count_3_io_out ? io_r_37_b : _GEN_486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_488 = 7'h26 == r_count_3_io_out ? io_r_38_b : _GEN_487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_489 = 7'h27 == r_count_3_io_out ? io_r_39_b : _GEN_488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_490 = 7'h28 == r_count_3_io_out ? io_r_40_b : _GEN_489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_491 = 7'h29 == r_count_3_io_out ? io_r_41_b : _GEN_490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_492 = 7'h2a == r_count_3_io_out ? io_r_42_b : _GEN_491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_493 = 7'h2b == r_count_3_io_out ? io_r_43_b : _GEN_492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_494 = 7'h2c == r_count_3_io_out ? io_r_44_b : _GEN_493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_495 = 7'h2d == r_count_3_io_out ? io_r_45_b : _GEN_494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_496 = 7'h2e == r_count_3_io_out ? io_r_46_b : _GEN_495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_497 = 7'h2f == r_count_3_io_out ? io_r_47_b : _GEN_496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_498 = 7'h30 == r_count_3_io_out ? io_r_48_b : _GEN_497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_499 = 7'h31 == r_count_3_io_out ? io_r_49_b : _GEN_498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_500 = 7'h32 == r_count_3_io_out ? io_r_50_b : _GEN_499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_501 = 7'h33 == r_count_3_io_out ? io_r_51_b : _GEN_500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_502 = 7'h34 == r_count_3_io_out ? io_r_52_b : _GEN_501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_503 = 7'h35 == r_count_3_io_out ? io_r_53_b : _GEN_502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_504 = 7'h36 == r_count_3_io_out ? io_r_54_b : _GEN_503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_505 = 7'h37 == r_count_3_io_out ? io_r_55_b : _GEN_504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_506 = 7'h38 == r_count_3_io_out ? io_r_56_b : _GEN_505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_507 = 7'h39 == r_count_3_io_out ? io_r_57_b : _GEN_506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_508 = 7'h3a == r_count_3_io_out ? io_r_58_b : _GEN_507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_509 = 7'h3b == r_count_3_io_out ? io_r_59_b : _GEN_508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_510 = 7'h3c == r_count_3_io_out ? io_r_60_b : _GEN_509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_511 = 7'h3d == r_count_3_io_out ? io_r_61_b : _GEN_510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_512 = 7'h3e == r_count_3_io_out ? io_r_62_b : _GEN_511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_513 = 7'h3f == r_count_3_io_out ? io_r_63_b : _GEN_512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_514 = 7'h40 == r_count_3_io_out ? io_r_64_b : _GEN_513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_515 = 7'h41 == r_count_3_io_out ? io_r_65_b : _GEN_514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_516 = 7'h42 == r_count_3_io_out ? io_r_66_b : _GEN_515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_517 = 7'h43 == r_count_3_io_out ? io_r_67_b : _GEN_516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_518 = 7'h44 == r_count_3_io_out ? io_r_68_b : _GEN_517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_519 = 7'h45 == r_count_3_io_out ? io_r_69_b : _GEN_518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_520 = 7'h46 == r_count_3_io_out ? io_r_70_b : _GEN_519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_521 = 7'h47 == r_count_3_io_out ? io_r_71_b : _GEN_520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_522 = 7'h48 == r_count_3_io_out ? io_r_72_b : _GEN_521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_523 = 7'h49 == r_count_3_io_out ? io_r_73_b : _GEN_522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_524 = 7'h4a == r_count_3_io_out ? io_r_74_b : _GEN_523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_525 = 7'h4b == r_count_3_io_out ? io_r_75_b : _GEN_524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_526 = 7'h4c == r_count_3_io_out ? io_r_76_b : _GEN_525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_527 = 7'h4d == r_count_3_io_out ? io_r_77_b : _GEN_526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_528 = 7'h4e == r_count_3_io_out ? io_r_78_b : _GEN_527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_529 = 7'h4f == r_count_3_io_out ? io_r_79_b : _GEN_528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_530 = 7'h50 == r_count_3_io_out ? io_r_80_b : _GEN_529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_531 = 7'h51 == r_count_3_io_out ? io_r_81_b : _GEN_530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_532 = 7'h52 == r_count_3_io_out ? io_r_82_b : _GEN_531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_533 = 7'h53 == r_count_3_io_out ? io_r_83_b : _GEN_532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_534 = 7'h54 == r_count_3_io_out ? io_r_84_b : _GEN_533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_535 = 7'h55 == r_count_3_io_out ? io_r_85_b : _GEN_534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_536 = 7'h56 == r_count_3_io_out ? io_r_86_b : _GEN_535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_537 = 7'h57 == r_count_3_io_out ? io_r_87_b : _GEN_536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_538 = 7'h58 == r_count_3_io_out ? io_r_88_b : _GEN_537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_539 = 7'h59 == r_count_3_io_out ? io_r_89_b : _GEN_538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_540 = 7'h5a == r_count_3_io_out ? io_r_90_b : _GEN_539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_541 = 7'h5b == r_count_3_io_out ? io_r_91_b : _GEN_540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_542 = 7'h5c == r_count_3_io_out ? io_r_92_b : _GEN_541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_543 = 7'h5d == r_count_3_io_out ? io_r_93_b : _GEN_542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_544 = 7'h5e == r_count_3_io_out ? io_r_94_b : _GEN_543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_545 = 7'h5f == r_count_3_io_out ? io_r_95_b : _GEN_544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_546 = 7'h60 == r_count_3_io_out ? io_r_96_b : _GEN_545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_547 = 7'h61 == r_count_3_io_out ? io_r_97_b : _GEN_546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_548 = 7'h62 == r_count_3_io_out ? io_r_98_b : _GEN_547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_551 = 7'h1 == r_count_4_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_552 = 7'h2 == r_count_4_io_out ? io_r_2_b : _GEN_551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_553 = 7'h3 == r_count_4_io_out ? io_r_3_b : _GEN_552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_554 = 7'h4 == r_count_4_io_out ? io_r_4_b : _GEN_553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_555 = 7'h5 == r_count_4_io_out ? io_r_5_b : _GEN_554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_556 = 7'h6 == r_count_4_io_out ? io_r_6_b : _GEN_555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_557 = 7'h7 == r_count_4_io_out ? io_r_7_b : _GEN_556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_558 = 7'h8 == r_count_4_io_out ? io_r_8_b : _GEN_557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_559 = 7'h9 == r_count_4_io_out ? io_r_9_b : _GEN_558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_560 = 7'ha == r_count_4_io_out ? io_r_10_b : _GEN_559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_561 = 7'hb == r_count_4_io_out ? io_r_11_b : _GEN_560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_562 = 7'hc == r_count_4_io_out ? io_r_12_b : _GEN_561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_563 = 7'hd == r_count_4_io_out ? io_r_13_b : _GEN_562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_564 = 7'he == r_count_4_io_out ? io_r_14_b : _GEN_563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_565 = 7'hf == r_count_4_io_out ? io_r_15_b : _GEN_564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_566 = 7'h10 == r_count_4_io_out ? io_r_16_b : _GEN_565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_567 = 7'h11 == r_count_4_io_out ? io_r_17_b : _GEN_566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_568 = 7'h12 == r_count_4_io_out ? io_r_18_b : _GEN_567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_569 = 7'h13 == r_count_4_io_out ? io_r_19_b : _GEN_568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_570 = 7'h14 == r_count_4_io_out ? io_r_20_b : _GEN_569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_571 = 7'h15 == r_count_4_io_out ? io_r_21_b : _GEN_570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_572 = 7'h16 == r_count_4_io_out ? io_r_22_b : _GEN_571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_573 = 7'h17 == r_count_4_io_out ? io_r_23_b : _GEN_572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_574 = 7'h18 == r_count_4_io_out ? io_r_24_b : _GEN_573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_575 = 7'h19 == r_count_4_io_out ? io_r_25_b : _GEN_574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_576 = 7'h1a == r_count_4_io_out ? io_r_26_b : _GEN_575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_577 = 7'h1b == r_count_4_io_out ? io_r_27_b : _GEN_576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_578 = 7'h1c == r_count_4_io_out ? io_r_28_b : _GEN_577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_579 = 7'h1d == r_count_4_io_out ? io_r_29_b : _GEN_578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_580 = 7'h1e == r_count_4_io_out ? io_r_30_b : _GEN_579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_581 = 7'h1f == r_count_4_io_out ? io_r_31_b : _GEN_580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_582 = 7'h20 == r_count_4_io_out ? io_r_32_b : _GEN_581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_583 = 7'h21 == r_count_4_io_out ? io_r_33_b : _GEN_582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_584 = 7'h22 == r_count_4_io_out ? io_r_34_b : _GEN_583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_585 = 7'h23 == r_count_4_io_out ? io_r_35_b : _GEN_584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_586 = 7'h24 == r_count_4_io_out ? io_r_36_b : _GEN_585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_587 = 7'h25 == r_count_4_io_out ? io_r_37_b : _GEN_586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_588 = 7'h26 == r_count_4_io_out ? io_r_38_b : _GEN_587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_589 = 7'h27 == r_count_4_io_out ? io_r_39_b : _GEN_588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_590 = 7'h28 == r_count_4_io_out ? io_r_40_b : _GEN_589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_591 = 7'h29 == r_count_4_io_out ? io_r_41_b : _GEN_590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_592 = 7'h2a == r_count_4_io_out ? io_r_42_b : _GEN_591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_593 = 7'h2b == r_count_4_io_out ? io_r_43_b : _GEN_592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_594 = 7'h2c == r_count_4_io_out ? io_r_44_b : _GEN_593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_595 = 7'h2d == r_count_4_io_out ? io_r_45_b : _GEN_594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_596 = 7'h2e == r_count_4_io_out ? io_r_46_b : _GEN_595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_597 = 7'h2f == r_count_4_io_out ? io_r_47_b : _GEN_596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_598 = 7'h30 == r_count_4_io_out ? io_r_48_b : _GEN_597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_599 = 7'h31 == r_count_4_io_out ? io_r_49_b : _GEN_598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_600 = 7'h32 == r_count_4_io_out ? io_r_50_b : _GEN_599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_601 = 7'h33 == r_count_4_io_out ? io_r_51_b : _GEN_600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_602 = 7'h34 == r_count_4_io_out ? io_r_52_b : _GEN_601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_603 = 7'h35 == r_count_4_io_out ? io_r_53_b : _GEN_602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_604 = 7'h36 == r_count_4_io_out ? io_r_54_b : _GEN_603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_605 = 7'h37 == r_count_4_io_out ? io_r_55_b : _GEN_604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_606 = 7'h38 == r_count_4_io_out ? io_r_56_b : _GEN_605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_607 = 7'h39 == r_count_4_io_out ? io_r_57_b : _GEN_606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_608 = 7'h3a == r_count_4_io_out ? io_r_58_b : _GEN_607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_609 = 7'h3b == r_count_4_io_out ? io_r_59_b : _GEN_608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_610 = 7'h3c == r_count_4_io_out ? io_r_60_b : _GEN_609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_611 = 7'h3d == r_count_4_io_out ? io_r_61_b : _GEN_610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_612 = 7'h3e == r_count_4_io_out ? io_r_62_b : _GEN_611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_613 = 7'h3f == r_count_4_io_out ? io_r_63_b : _GEN_612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_614 = 7'h40 == r_count_4_io_out ? io_r_64_b : _GEN_613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_615 = 7'h41 == r_count_4_io_out ? io_r_65_b : _GEN_614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_616 = 7'h42 == r_count_4_io_out ? io_r_66_b : _GEN_615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_617 = 7'h43 == r_count_4_io_out ? io_r_67_b : _GEN_616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_618 = 7'h44 == r_count_4_io_out ? io_r_68_b : _GEN_617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_619 = 7'h45 == r_count_4_io_out ? io_r_69_b : _GEN_618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_620 = 7'h46 == r_count_4_io_out ? io_r_70_b : _GEN_619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_621 = 7'h47 == r_count_4_io_out ? io_r_71_b : _GEN_620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_622 = 7'h48 == r_count_4_io_out ? io_r_72_b : _GEN_621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_623 = 7'h49 == r_count_4_io_out ? io_r_73_b : _GEN_622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_624 = 7'h4a == r_count_4_io_out ? io_r_74_b : _GEN_623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_625 = 7'h4b == r_count_4_io_out ? io_r_75_b : _GEN_624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_626 = 7'h4c == r_count_4_io_out ? io_r_76_b : _GEN_625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_627 = 7'h4d == r_count_4_io_out ? io_r_77_b : _GEN_626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_628 = 7'h4e == r_count_4_io_out ? io_r_78_b : _GEN_627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_629 = 7'h4f == r_count_4_io_out ? io_r_79_b : _GEN_628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_630 = 7'h50 == r_count_4_io_out ? io_r_80_b : _GEN_629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_631 = 7'h51 == r_count_4_io_out ? io_r_81_b : _GEN_630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_632 = 7'h52 == r_count_4_io_out ? io_r_82_b : _GEN_631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_633 = 7'h53 == r_count_4_io_out ? io_r_83_b : _GEN_632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_634 = 7'h54 == r_count_4_io_out ? io_r_84_b : _GEN_633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_635 = 7'h55 == r_count_4_io_out ? io_r_85_b : _GEN_634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_636 = 7'h56 == r_count_4_io_out ? io_r_86_b : _GEN_635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_637 = 7'h57 == r_count_4_io_out ? io_r_87_b : _GEN_636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_638 = 7'h58 == r_count_4_io_out ? io_r_88_b : _GEN_637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_639 = 7'h59 == r_count_4_io_out ? io_r_89_b : _GEN_638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_640 = 7'h5a == r_count_4_io_out ? io_r_90_b : _GEN_639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_641 = 7'h5b == r_count_4_io_out ? io_r_91_b : _GEN_640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_642 = 7'h5c == r_count_4_io_out ? io_r_92_b : _GEN_641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_643 = 7'h5d == r_count_4_io_out ? io_r_93_b : _GEN_642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_644 = 7'h5e == r_count_4_io_out ? io_r_94_b : _GEN_643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_645 = 7'h5f == r_count_4_io_out ? io_r_95_b : _GEN_644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_646 = 7'h60 == r_count_4_io_out ? io_r_96_b : _GEN_645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_647 = 7'h61 == r_count_4_io_out ? io_r_97_b : _GEN_646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_648 = 7'h62 == r_count_4_io_out ? io_r_98_b : _GEN_647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_651 = 7'h1 == r_count_5_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_652 = 7'h2 == r_count_5_io_out ? io_r_2_b : _GEN_651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_653 = 7'h3 == r_count_5_io_out ? io_r_3_b : _GEN_652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_654 = 7'h4 == r_count_5_io_out ? io_r_4_b : _GEN_653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_655 = 7'h5 == r_count_5_io_out ? io_r_5_b : _GEN_654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_656 = 7'h6 == r_count_5_io_out ? io_r_6_b : _GEN_655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_657 = 7'h7 == r_count_5_io_out ? io_r_7_b : _GEN_656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_658 = 7'h8 == r_count_5_io_out ? io_r_8_b : _GEN_657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_659 = 7'h9 == r_count_5_io_out ? io_r_9_b : _GEN_658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_660 = 7'ha == r_count_5_io_out ? io_r_10_b : _GEN_659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_661 = 7'hb == r_count_5_io_out ? io_r_11_b : _GEN_660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_662 = 7'hc == r_count_5_io_out ? io_r_12_b : _GEN_661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_663 = 7'hd == r_count_5_io_out ? io_r_13_b : _GEN_662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_664 = 7'he == r_count_5_io_out ? io_r_14_b : _GEN_663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_665 = 7'hf == r_count_5_io_out ? io_r_15_b : _GEN_664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_666 = 7'h10 == r_count_5_io_out ? io_r_16_b : _GEN_665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_667 = 7'h11 == r_count_5_io_out ? io_r_17_b : _GEN_666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_668 = 7'h12 == r_count_5_io_out ? io_r_18_b : _GEN_667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_669 = 7'h13 == r_count_5_io_out ? io_r_19_b : _GEN_668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_670 = 7'h14 == r_count_5_io_out ? io_r_20_b : _GEN_669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_671 = 7'h15 == r_count_5_io_out ? io_r_21_b : _GEN_670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_672 = 7'h16 == r_count_5_io_out ? io_r_22_b : _GEN_671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_673 = 7'h17 == r_count_5_io_out ? io_r_23_b : _GEN_672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_674 = 7'h18 == r_count_5_io_out ? io_r_24_b : _GEN_673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_675 = 7'h19 == r_count_5_io_out ? io_r_25_b : _GEN_674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_676 = 7'h1a == r_count_5_io_out ? io_r_26_b : _GEN_675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_677 = 7'h1b == r_count_5_io_out ? io_r_27_b : _GEN_676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_678 = 7'h1c == r_count_5_io_out ? io_r_28_b : _GEN_677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_679 = 7'h1d == r_count_5_io_out ? io_r_29_b : _GEN_678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_680 = 7'h1e == r_count_5_io_out ? io_r_30_b : _GEN_679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_681 = 7'h1f == r_count_5_io_out ? io_r_31_b : _GEN_680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_682 = 7'h20 == r_count_5_io_out ? io_r_32_b : _GEN_681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_683 = 7'h21 == r_count_5_io_out ? io_r_33_b : _GEN_682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_684 = 7'h22 == r_count_5_io_out ? io_r_34_b : _GEN_683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_685 = 7'h23 == r_count_5_io_out ? io_r_35_b : _GEN_684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_686 = 7'h24 == r_count_5_io_out ? io_r_36_b : _GEN_685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_687 = 7'h25 == r_count_5_io_out ? io_r_37_b : _GEN_686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_688 = 7'h26 == r_count_5_io_out ? io_r_38_b : _GEN_687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_689 = 7'h27 == r_count_5_io_out ? io_r_39_b : _GEN_688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_690 = 7'h28 == r_count_5_io_out ? io_r_40_b : _GEN_689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_691 = 7'h29 == r_count_5_io_out ? io_r_41_b : _GEN_690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_692 = 7'h2a == r_count_5_io_out ? io_r_42_b : _GEN_691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_693 = 7'h2b == r_count_5_io_out ? io_r_43_b : _GEN_692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_694 = 7'h2c == r_count_5_io_out ? io_r_44_b : _GEN_693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_695 = 7'h2d == r_count_5_io_out ? io_r_45_b : _GEN_694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_696 = 7'h2e == r_count_5_io_out ? io_r_46_b : _GEN_695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_697 = 7'h2f == r_count_5_io_out ? io_r_47_b : _GEN_696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_698 = 7'h30 == r_count_5_io_out ? io_r_48_b : _GEN_697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_699 = 7'h31 == r_count_5_io_out ? io_r_49_b : _GEN_698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_700 = 7'h32 == r_count_5_io_out ? io_r_50_b : _GEN_699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_701 = 7'h33 == r_count_5_io_out ? io_r_51_b : _GEN_700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_702 = 7'h34 == r_count_5_io_out ? io_r_52_b : _GEN_701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_703 = 7'h35 == r_count_5_io_out ? io_r_53_b : _GEN_702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_704 = 7'h36 == r_count_5_io_out ? io_r_54_b : _GEN_703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_705 = 7'h37 == r_count_5_io_out ? io_r_55_b : _GEN_704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_706 = 7'h38 == r_count_5_io_out ? io_r_56_b : _GEN_705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_707 = 7'h39 == r_count_5_io_out ? io_r_57_b : _GEN_706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_708 = 7'h3a == r_count_5_io_out ? io_r_58_b : _GEN_707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_709 = 7'h3b == r_count_5_io_out ? io_r_59_b : _GEN_708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_710 = 7'h3c == r_count_5_io_out ? io_r_60_b : _GEN_709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_711 = 7'h3d == r_count_5_io_out ? io_r_61_b : _GEN_710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_712 = 7'h3e == r_count_5_io_out ? io_r_62_b : _GEN_711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_713 = 7'h3f == r_count_5_io_out ? io_r_63_b : _GEN_712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_714 = 7'h40 == r_count_5_io_out ? io_r_64_b : _GEN_713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_715 = 7'h41 == r_count_5_io_out ? io_r_65_b : _GEN_714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_716 = 7'h42 == r_count_5_io_out ? io_r_66_b : _GEN_715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_717 = 7'h43 == r_count_5_io_out ? io_r_67_b : _GEN_716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_718 = 7'h44 == r_count_5_io_out ? io_r_68_b : _GEN_717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_719 = 7'h45 == r_count_5_io_out ? io_r_69_b : _GEN_718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_720 = 7'h46 == r_count_5_io_out ? io_r_70_b : _GEN_719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_721 = 7'h47 == r_count_5_io_out ? io_r_71_b : _GEN_720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_722 = 7'h48 == r_count_5_io_out ? io_r_72_b : _GEN_721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_723 = 7'h49 == r_count_5_io_out ? io_r_73_b : _GEN_722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_724 = 7'h4a == r_count_5_io_out ? io_r_74_b : _GEN_723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_725 = 7'h4b == r_count_5_io_out ? io_r_75_b : _GEN_724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_726 = 7'h4c == r_count_5_io_out ? io_r_76_b : _GEN_725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_727 = 7'h4d == r_count_5_io_out ? io_r_77_b : _GEN_726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_728 = 7'h4e == r_count_5_io_out ? io_r_78_b : _GEN_727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_729 = 7'h4f == r_count_5_io_out ? io_r_79_b : _GEN_728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_730 = 7'h50 == r_count_5_io_out ? io_r_80_b : _GEN_729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_731 = 7'h51 == r_count_5_io_out ? io_r_81_b : _GEN_730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_732 = 7'h52 == r_count_5_io_out ? io_r_82_b : _GEN_731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_733 = 7'h53 == r_count_5_io_out ? io_r_83_b : _GEN_732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_734 = 7'h54 == r_count_5_io_out ? io_r_84_b : _GEN_733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_735 = 7'h55 == r_count_5_io_out ? io_r_85_b : _GEN_734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_736 = 7'h56 == r_count_5_io_out ? io_r_86_b : _GEN_735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_737 = 7'h57 == r_count_5_io_out ? io_r_87_b : _GEN_736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_738 = 7'h58 == r_count_5_io_out ? io_r_88_b : _GEN_737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_739 = 7'h59 == r_count_5_io_out ? io_r_89_b : _GEN_738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_740 = 7'h5a == r_count_5_io_out ? io_r_90_b : _GEN_739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_741 = 7'h5b == r_count_5_io_out ? io_r_91_b : _GEN_740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_742 = 7'h5c == r_count_5_io_out ? io_r_92_b : _GEN_741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_743 = 7'h5d == r_count_5_io_out ? io_r_93_b : _GEN_742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_744 = 7'h5e == r_count_5_io_out ? io_r_94_b : _GEN_743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_745 = 7'h5f == r_count_5_io_out ? io_r_95_b : _GEN_744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_746 = 7'h60 == r_count_5_io_out ? io_r_96_b : _GEN_745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_747 = 7'h61 == r_count_5_io_out ? io_r_97_b : _GEN_746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_748 = 7'h62 == r_count_5_io_out ? io_r_98_b : _GEN_747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_751 = 7'h1 == r_count_6_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_752 = 7'h2 == r_count_6_io_out ? io_r_2_b : _GEN_751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_753 = 7'h3 == r_count_6_io_out ? io_r_3_b : _GEN_752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_754 = 7'h4 == r_count_6_io_out ? io_r_4_b : _GEN_753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_755 = 7'h5 == r_count_6_io_out ? io_r_5_b : _GEN_754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_756 = 7'h6 == r_count_6_io_out ? io_r_6_b : _GEN_755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_757 = 7'h7 == r_count_6_io_out ? io_r_7_b : _GEN_756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_758 = 7'h8 == r_count_6_io_out ? io_r_8_b : _GEN_757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_759 = 7'h9 == r_count_6_io_out ? io_r_9_b : _GEN_758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_760 = 7'ha == r_count_6_io_out ? io_r_10_b : _GEN_759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_761 = 7'hb == r_count_6_io_out ? io_r_11_b : _GEN_760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_762 = 7'hc == r_count_6_io_out ? io_r_12_b : _GEN_761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_763 = 7'hd == r_count_6_io_out ? io_r_13_b : _GEN_762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_764 = 7'he == r_count_6_io_out ? io_r_14_b : _GEN_763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_765 = 7'hf == r_count_6_io_out ? io_r_15_b : _GEN_764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_766 = 7'h10 == r_count_6_io_out ? io_r_16_b : _GEN_765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_767 = 7'h11 == r_count_6_io_out ? io_r_17_b : _GEN_766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_768 = 7'h12 == r_count_6_io_out ? io_r_18_b : _GEN_767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_769 = 7'h13 == r_count_6_io_out ? io_r_19_b : _GEN_768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_770 = 7'h14 == r_count_6_io_out ? io_r_20_b : _GEN_769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_771 = 7'h15 == r_count_6_io_out ? io_r_21_b : _GEN_770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_772 = 7'h16 == r_count_6_io_out ? io_r_22_b : _GEN_771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_773 = 7'h17 == r_count_6_io_out ? io_r_23_b : _GEN_772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_774 = 7'h18 == r_count_6_io_out ? io_r_24_b : _GEN_773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_775 = 7'h19 == r_count_6_io_out ? io_r_25_b : _GEN_774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_776 = 7'h1a == r_count_6_io_out ? io_r_26_b : _GEN_775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_777 = 7'h1b == r_count_6_io_out ? io_r_27_b : _GEN_776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_778 = 7'h1c == r_count_6_io_out ? io_r_28_b : _GEN_777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_779 = 7'h1d == r_count_6_io_out ? io_r_29_b : _GEN_778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_780 = 7'h1e == r_count_6_io_out ? io_r_30_b : _GEN_779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_781 = 7'h1f == r_count_6_io_out ? io_r_31_b : _GEN_780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_782 = 7'h20 == r_count_6_io_out ? io_r_32_b : _GEN_781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_783 = 7'h21 == r_count_6_io_out ? io_r_33_b : _GEN_782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_784 = 7'h22 == r_count_6_io_out ? io_r_34_b : _GEN_783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_785 = 7'h23 == r_count_6_io_out ? io_r_35_b : _GEN_784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_786 = 7'h24 == r_count_6_io_out ? io_r_36_b : _GEN_785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_787 = 7'h25 == r_count_6_io_out ? io_r_37_b : _GEN_786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_788 = 7'h26 == r_count_6_io_out ? io_r_38_b : _GEN_787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_789 = 7'h27 == r_count_6_io_out ? io_r_39_b : _GEN_788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_790 = 7'h28 == r_count_6_io_out ? io_r_40_b : _GEN_789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_791 = 7'h29 == r_count_6_io_out ? io_r_41_b : _GEN_790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_792 = 7'h2a == r_count_6_io_out ? io_r_42_b : _GEN_791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_793 = 7'h2b == r_count_6_io_out ? io_r_43_b : _GEN_792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_794 = 7'h2c == r_count_6_io_out ? io_r_44_b : _GEN_793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_795 = 7'h2d == r_count_6_io_out ? io_r_45_b : _GEN_794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_796 = 7'h2e == r_count_6_io_out ? io_r_46_b : _GEN_795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_797 = 7'h2f == r_count_6_io_out ? io_r_47_b : _GEN_796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_798 = 7'h30 == r_count_6_io_out ? io_r_48_b : _GEN_797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_799 = 7'h31 == r_count_6_io_out ? io_r_49_b : _GEN_798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_800 = 7'h32 == r_count_6_io_out ? io_r_50_b : _GEN_799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_801 = 7'h33 == r_count_6_io_out ? io_r_51_b : _GEN_800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_802 = 7'h34 == r_count_6_io_out ? io_r_52_b : _GEN_801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_803 = 7'h35 == r_count_6_io_out ? io_r_53_b : _GEN_802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_804 = 7'h36 == r_count_6_io_out ? io_r_54_b : _GEN_803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_805 = 7'h37 == r_count_6_io_out ? io_r_55_b : _GEN_804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_806 = 7'h38 == r_count_6_io_out ? io_r_56_b : _GEN_805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_807 = 7'h39 == r_count_6_io_out ? io_r_57_b : _GEN_806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_808 = 7'h3a == r_count_6_io_out ? io_r_58_b : _GEN_807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_809 = 7'h3b == r_count_6_io_out ? io_r_59_b : _GEN_808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_810 = 7'h3c == r_count_6_io_out ? io_r_60_b : _GEN_809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_811 = 7'h3d == r_count_6_io_out ? io_r_61_b : _GEN_810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_812 = 7'h3e == r_count_6_io_out ? io_r_62_b : _GEN_811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_813 = 7'h3f == r_count_6_io_out ? io_r_63_b : _GEN_812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_814 = 7'h40 == r_count_6_io_out ? io_r_64_b : _GEN_813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_815 = 7'h41 == r_count_6_io_out ? io_r_65_b : _GEN_814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_816 = 7'h42 == r_count_6_io_out ? io_r_66_b : _GEN_815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_817 = 7'h43 == r_count_6_io_out ? io_r_67_b : _GEN_816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_818 = 7'h44 == r_count_6_io_out ? io_r_68_b : _GEN_817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_819 = 7'h45 == r_count_6_io_out ? io_r_69_b : _GEN_818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_820 = 7'h46 == r_count_6_io_out ? io_r_70_b : _GEN_819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_821 = 7'h47 == r_count_6_io_out ? io_r_71_b : _GEN_820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_822 = 7'h48 == r_count_6_io_out ? io_r_72_b : _GEN_821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_823 = 7'h49 == r_count_6_io_out ? io_r_73_b : _GEN_822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_824 = 7'h4a == r_count_6_io_out ? io_r_74_b : _GEN_823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_825 = 7'h4b == r_count_6_io_out ? io_r_75_b : _GEN_824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_826 = 7'h4c == r_count_6_io_out ? io_r_76_b : _GEN_825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_827 = 7'h4d == r_count_6_io_out ? io_r_77_b : _GEN_826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_828 = 7'h4e == r_count_6_io_out ? io_r_78_b : _GEN_827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_829 = 7'h4f == r_count_6_io_out ? io_r_79_b : _GEN_828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_830 = 7'h50 == r_count_6_io_out ? io_r_80_b : _GEN_829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_831 = 7'h51 == r_count_6_io_out ? io_r_81_b : _GEN_830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_832 = 7'h52 == r_count_6_io_out ? io_r_82_b : _GEN_831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_833 = 7'h53 == r_count_6_io_out ? io_r_83_b : _GEN_832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_834 = 7'h54 == r_count_6_io_out ? io_r_84_b : _GEN_833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_835 = 7'h55 == r_count_6_io_out ? io_r_85_b : _GEN_834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_836 = 7'h56 == r_count_6_io_out ? io_r_86_b : _GEN_835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_837 = 7'h57 == r_count_6_io_out ? io_r_87_b : _GEN_836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_838 = 7'h58 == r_count_6_io_out ? io_r_88_b : _GEN_837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_839 = 7'h59 == r_count_6_io_out ? io_r_89_b : _GEN_838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_840 = 7'h5a == r_count_6_io_out ? io_r_90_b : _GEN_839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_841 = 7'h5b == r_count_6_io_out ? io_r_91_b : _GEN_840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_842 = 7'h5c == r_count_6_io_out ? io_r_92_b : _GEN_841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_843 = 7'h5d == r_count_6_io_out ? io_r_93_b : _GEN_842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_844 = 7'h5e == r_count_6_io_out ? io_r_94_b : _GEN_843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_845 = 7'h5f == r_count_6_io_out ? io_r_95_b : _GEN_844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_846 = 7'h60 == r_count_6_io_out ? io_r_96_b : _GEN_845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_847 = 7'h61 == r_count_6_io_out ? io_r_97_b : _GEN_846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_848 = 7'h62 == r_count_6_io_out ? io_r_98_b : _GEN_847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_851 = 7'h1 == r_count_7_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_852 = 7'h2 == r_count_7_io_out ? io_r_2_b : _GEN_851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_853 = 7'h3 == r_count_7_io_out ? io_r_3_b : _GEN_852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_854 = 7'h4 == r_count_7_io_out ? io_r_4_b : _GEN_853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_855 = 7'h5 == r_count_7_io_out ? io_r_5_b : _GEN_854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_856 = 7'h6 == r_count_7_io_out ? io_r_6_b : _GEN_855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_857 = 7'h7 == r_count_7_io_out ? io_r_7_b : _GEN_856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_858 = 7'h8 == r_count_7_io_out ? io_r_8_b : _GEN_857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_859 = 7'h9 == r_count_7_io_out ? io_r_9_b : _GEN_858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_860 = 7'ha == r_count_7_io_out ? io_r_10_b : _GEN_859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_861 = 7'hb == r_count_7_io_out ? io_r_11_b : _GEN_860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_862 = 7'hc == r_count_7_io_out ? io_r_12_b : _GEN_861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_863 = 7'hd == r_count_7_io_out ? io_r_13_b : _GEN_862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_864 = 7'he == r_count_7_io_out ? io_r_14_b : _GEN_863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_865 = 7'hf == r_count_7_io_out ? io_r_15_b : _GEN_864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_866 = 7'h10 == r_count_7_io_out ? io_r_16_b : _GEN_865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_867 = 7'h11 == r_count_7_io_out ? io_r_17_b : _GEN_866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_868 = 7'h12 == r_count_7_io_out ? io_r_18_b : _GEN_867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_869 = 7'h13 == r_count_7_io_out ? io_r_19_b : _GEN_868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_870 = 7'h14 == r_count_7_io_out ? io_r_20_b : _GEN_869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_871 = 7'h15 == r_count_7_io_out ? io_r_21_b : _GEN_870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_872 = 7'h16 == r_count_7_io_out ? io_r_22_b : _GEN_871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_873 = 7'h17 == r_count_7_io_out ? io_r_23_b : _GEN_872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_874 = 7'h18 == r_count_7_io_out ? io_r_24_b : _GEN_873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_875 = 7'h19 == r_count_7_io_out ? io_r_25_b : _GEN_874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_876 = 7'h1a == r_count_7_io_out ? io_r_26_b : _GEN_875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_877 = 7'h1b == r_count_7_io_out ? io_r_27_b : _GEN_876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_878 = 7'h1c == r_count_7_io_out ? io_r_28_b : _GEN_877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_879 = 7'h1d == r_count_7_io_out ? io_r_29_b : _GEN_878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_880 = 7'h1e == r_count_7_io_out ? io_r_30_b : _GEN_879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_881 = 7'h1f == r_count_7_io_out ? io_r_31_b : _GEN_880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_882 = 7'h20 == r_count_7_io_out ? io_r_32_b : _GEN_881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_883 = 7'h21 == r_count_7_io_out ? io_r_33_b : _GEN_882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_884 = 7'h22 == r_count_7_io_out ? io_r_34_b : _GEN_883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_885 = 7'h23 == r_count_7_io_out ? io_r_35_b : _GEN_884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_886 = 7'h24 == r_count_7_io_out ? io_r_36_b : _GEN_885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_887 = 7'h25 == r_count_7_io_out ? io_r_37_b : _GEN_886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_888 = 7'h26 == r_count_7_io_out ? io_r_38_b : _GEN_887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_889 = 7'h27 == r_count_7_io_out ? io_r_39_b : _GEN_888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_890 = 7'h28 == r_count_7_io_out ? io_r_40_b : _GEN_889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_891 = 7'h29 == r_count_7_io_out ? io_r_41_b : _GEN_890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_892 = 7'h2a == r_count_7_io_out ? io_r_42_b : _GEN_891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_893 = 7'h2b == r_count_7_io_out ? io_r_43_b : _GEN_892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_894 = 7'h2c == r_count_7_io_out ? io_r_44_b : _GEN_893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_895 = 7'h2d == r_count_7_io_out ? io_r_45_b : _GEN_894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_896 = 7'h2e == r_count_7_io_out ? io_r_46_b : _GEN_895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_897 = 7'h2f == r_count_7_io_out ? io_r_47_b : _GEN_896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_898 = 7'h30 == r_count_7_io_out ? io_r_48_b : _GEN_897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_899 = 7'h31 == r_count_7_io_out ? io_r_49_b : _GEN_898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_900 = 7'h32 == r_count_7_io_out ? io_r_50_b : _GEN_899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_901 = 7'h33 == r_count_7_io_out ? io_r_51_b : _GEN_900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_902 = 7'h34 == r_count_7_io_out ? io_r_52_b : _GEN_901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_903 = 7'h35 == r_count_7_io_out ? io_r_53_b : _GEN_902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_904 = 7'h36 == r_count_7_io_out ? io_r_54_b : _GEN_903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_905 = 7'h37 == r_count_7_io_out ? io_r_55_b : _GEN_904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_906 = 7'h38 == r_count_7_io_out ? io_r_56_b : _GEN_905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_907 = 7'h39 == r_count_7_io_out ? io_r_57_b : _GEN_906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_908 = 7'h3a == r_count_7_io_out ? io_r_58_b : _GEN_907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_909 = 7'h3b == r_count_7_io_out ? io_r_59_b : _GEN_908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_910 = 7'h3c == r_count_7_io_out ? io_r_60_b : _GEN_909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_911 = 7'h3d == r_count_7_io_out ? io_r_61_b : _GEN_910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_912 = 7'h3e == r_count_7_io_out ? io_r_62_b : _GEN_911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_913 = 7'h3f == r_count_7_io_out ? io_r_63_b : _GEN_912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_914 = 7'h40 == r_count_7_io_out ? io_r_64_b : _GEN_913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_915 = 7'h41 == r_count_7_io_out ? io_r_65_b : _GEN_914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_916 = 7'h42 == r_count_7_io_out ? io_r_66_b : _GEN_915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_917 = 7'h43 == r_count_7_io_out ? io_r_67_b : _GEN_916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_918 = 7'h44 == r_count_7_io_out ? io_r_68_b : _GEN_917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_919 = 7'h45 == r_count_7_io_out ? io_r_69_b : _GEN_918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_920 = 7'h46 == r_count_7_io_out ? io_r_70_b : _GEN_919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_921 = 7'h47 == r_count_7_io_out ? io_r_71_b : _GEN_920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_922 = 7'h48 == r_count_7_io_out ? io_r_72_b : _GEN_921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_923 = 7'h49 == r_count_7_io_out ? io_r_73_b : _GEN_922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_924 = 7'h4a == r_count_7_io_out ? io_r_74_b : _GEN_923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_925 = 7'h4b == r_count_7_io_out ? io_r_75_b : _GEN_924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_926 = 7'h4c == r_count_7_io_out ? io_r_76_b : _GEN_925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_927 = 7'h4d == r_count_7_io_out ? io_r_77_b : _GEN_926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_928 = 7'h4e == r_count_7_io_out ? io_r_78_b : _GEN_927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_929 = 7'h4f == r_count_7_io_out ? io_r_79_b : _GEN_928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_930 = 7'h50 == r_count_7_io_out ? io_r_80_b : _GEN_929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_931 = 7'h51 == r_count_7_io_out ? io_r_81_b : _GEN_930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_932 = 7'h52 == r_count_7_io_out ? io_r_82_b : _GEN_931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_933 = 7'h53 == r_count_7_io_out ? io_r_83_b : _GEN_932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_934 = 7'h54 == r_count_7_io_out ? io_r_84_b : _GEN_933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_935 = 7'h55 == r_count_7_io_out ? io_r_85_b : _GEN_934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_936 = 7'h56 == r_count_7_io_out ? io_r_86_b : _GEN_935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_937 = 7'h57 == r_count_7_io_out ? io_r_87_b : _GEN_936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_938 = 7'h58 == r_count_7_io_out ? io_r_88_b : _GEN_937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_939 = 7'h59 == r_count_7_io_out ? io_r_89_b : _GEN_938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_940 = 7'h5a == r_count_7_io_out ? io_r_90_b : _GEN_939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_941 = 7'h5b == r_count_7_io_out ? io_r_91_b : _GEN_940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_942 = 7'h5c == r_count_7_io_out ? io_r_92_b : _GEN_941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_943 = 7'h5d == r_count_7_io_out ? io_r_93_b : _GEN_942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_944 = 7'h5e == r_count_7_io_out ? io_r_94_b : _GEN_943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_945 = 7'h5f == r_count_7_io_out ? io_r_95_b : _GEN_944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_946 = 7'h60 == r_count_7_io_out ? io_r_96_b : _GEN_945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_947 = 7'h61 == r_count_7_io_out ? io_r_97_b : _GEN_946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_948 = 7'h62 == r_count_7_io_out ? io_r_98_b : _GEN_947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_951 = 7'h1 == r_count_8_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_952 = 7'h2 == r_count_8_io_out ? io_r_2_b : _GEN_951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_953 = 7'h3 == r_count_8_io_out ? io_r_3_b : _GEN_952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_954 = 7'h4 == r_count_8_io_out ? io_r_4_b : _GEN_953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_955 = 7'h5 == r_count_8_io_out ? io_r_5_b : _GEN_954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_956 = 7'h6 == r_count_8_io_out ? io_r_6_b : _GEN_955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_957 = 7'h7 == r_count_8_io_out ? io_r_7_b : _GEN_956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_958 = 7'h8 == r_count_8_io_out ? io_r_8_b : _GEN_957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_959 = 7'h9 == r_count_8_io_out ? io_r_9_b : _GEN_958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_960 = 7'ha == r_count_8_io_out ? io_r_10_b : _GEN_959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_961 = 7'hb == r_count_8_io_out ? io_r_11_b : _GEN_960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_962 = 7'hc == r_count_8_io_out ? io_r_12_b : _GEN_961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_963 = 7'hd == r_count_8_io_out ? io_r_13_b : _GEN_962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_964 = 7'he == r_count_8_io_out ? io_r_14_b : _GEN_963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_965 = 7'hf == r_count_8_io_out ? io_r_15_b : _GEN_964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_966 = 7'h10 == r_count_8_io_out ? io_r_16_b : _GEN_965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_967 = 7'h11 == r_count_8_io_out ? io_r_17_b : _GEN_966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_968 = 7'h12 == r_count_8_io_out ? io_r_18_b : _GEN_967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_969 = 7'h13 == r_count_8_io_out ? io_r_19_b : _GEN_968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_970 = 7'h14 == r_count_8_io_out ? io_r_20_b : _GEN_969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_971 = 7'h15 == r_count_8_io_out ? io_r_21_b : _GEN_970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_972 = 7'h16 == r_count_8_io_out ? io_r_22_b : _GEN_971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_973 = 7'h17 == r_count_8_io_out ? io_r_23_b : _GEN_972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_974 = 7'h18 == r_count_8_io_out ? io_r_24_b : _GEN_973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_975 = 7'h19 == r_count_8_io_out ? io_r_25_b : _GEN_974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_976 = 7'h1a == r_count_8_io_out ? io_r_26_b : _GEN_975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_977 = 7'h1b == r_count_8_io_out ? io_r_27_b : _GEN_976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_978 = 7'h1c == r_count_8_io_out ? io_r_28_b : _GEN_977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_979 = 7'h1d == r_count_8_io_out ? io_r_29_b : _GEN_978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_980 = 7'h1e == r_count_8_io_out ? io_r_30_b : _GEN_979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_981 = 7'h1f == r_count_8_io_out ? io_r_31_b : _GEN_980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_982 = 7'h20 == r_count_8_io_out ? io_r_32_b : _GEN_981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_983 = 7'h21 == r_count_8_io_out ? io_r_33_b : _GEN_982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_984 = 7'h22 == r_count_8_io_out ? io_r_34_b : _GEN_983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_985 = 7'h23 == r_count_8_io_out ? io_r_35_b : _GEN_984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_986 = 7'h24 == r_count_8_io_out ? io_r_36_b : _GEN_985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_987 = 7'h25 == r_count_8_io_out ? io_r_37_b : _GEN_986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_988 = 7'h26 == r_count_8_io_out ? io_r_38_b : _GEN_987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_989 = 7'h27 == r_count_8_io_out ? io_r_39_b : _GEN_988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_990 = 7'h28 == r_count_8_io_out ? io_r_40_b : _GEN_989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_991 = 7'h29 == r_count_8_io_out ? io_r_41_b : _GEN_990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_992 = 7'h2a == r_count_8_io_out ? io_r_42_b : _GEN_991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_993 = 7'h2b == r_count_8_io_out ? io_r_43_b : _GEN_992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_994 = 7'h2c == r_count_8_io_out ? io_r_44_b : _GEN_993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_995 = 7'h2d == r_count_8_io_out ? io_r_45_b : _GEN_994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_996 = 7'h2e == r_count_8_io_out ? io_r_46_b : _GEN_995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_997 = 7'h2f == r_count_8_io_out ? io_r_47_b : _GEN_996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_998 = 7'h30 == r_count_8_io_out ? io_r_48_b : _GEN_997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_999 = 7'h31 == r_count_8_io_out ? io_r_49_b : _GEN_998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1000 = 7'h32 == r_count_8_io_out ? io_r_50_b : _GEN_999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1001 = 7'h33 == r_count_8_io_out ? io_r_51_b : _GEN_1000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1002 = 7'h34 == r_count_8_io_out ? io_r_52_b : _GEN_1001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1003 = 7'h35 == r_count_8_io_out ? io_r_53_b : _GEN_1002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1004 = 7'h36 == r_count_8_io_out ? io_r_54_b : _GEN_1003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1005 = 7'h37 == r_count_8_io_out ? io_r_55_b : _GEN_1004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1006 = 7'h38 == r_count_8_io_out ? io_r_56_b : _GEN_1005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1007 = 7'h39 == r_count_8_io_out ? io_r_57_b : _GEN_1006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1008 = 7'h3a == r_count_8_io_out ? io_r_58_b : _GEN_1007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1009 = 7'h3b == r_count_8_io_out ? io_r_59_b : _GEN_1008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1010 = 7'h3c == r_count_8_io_out ? io_r_60_b : _GEN_1009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1011 = 7'h3d == r_count_8_io_out ? io_r_61_b : _GEN_1010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1012 = 7'h3e == r_count_8_io_out ? io_r_62_b : _GEN_1011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1013 = 7'h3f == r_count_8_io_out ? io_r_63_b : _GEN_1012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1014 = 7'h40 == r_count_8_io_out ? io_r_64_b : _GEN_1013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1015 = 7'h41 == r_count_8_io_out ? io_r_65_b : _GEN_1014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1016 = 7'h42 == r_count_8_io_out ? io_r_66_b : _GEN_1015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1017 = 7'h43 == r_count_8_io_out ? io_r_67_b : _GEN_1016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1018 = 7'h44 == r_count_8_io_out ? io_r_68_b : _GEN_1017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1019 = 7'h45 == r_count_8_io_out ? io_r_69_b : _GEN_1018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1020 = 7'h46 == r_count_8_io_out ? io_r_70_b : _GEN_1019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1021 = 7'h47 == r_count_8_io_out ? io_r_71_b : _GEN_1020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1022 = 7'h48 == r_count_8_io_out ? io_r_72_b : _GEN_1021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1023 = 7'h49 == r_count_8_io_out ? io_r_73_b : _GEN_1022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1024 = 7'h4a == r_count_8_io_out ? io_r_74_b : _GEN_1023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1025 = 7'h4b == r_count_8_io_out ? io_r_75_b : _GEN_1024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1026 = 7'h4c == r_count_8_io_out ? io_r_76_b : _GEN_1025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1027 = 7'h4d == r_count_8_io_out ? io_r_77_b : _GEN_1026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1028 = 7'h4e == r_count_8_io_out ? io_r_78_b : _GEN_1027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1029 = 7'h4f == r_count_8_io_out ? io_r_79_b : _GEN_1028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1030 = 7'h50 == r_count_8_io_out ? io_r_80_b : _GEN_1029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1031 = 7'h51 == r_count_8_io_out ? io_r_81_b : _GEN_1030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1032 = 7'h52 == r_count_8_io_out ? io_r_82_b : _GEN_1031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1033 = 7'h53 == r_count_8_io_out ? io_r_83_b : _GEN_1032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1034 = 7'h54 == r_count_8_io_out ? io_r_84_b : _GEN_1033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1035 = 7'h55 == r_count_8_io_out ? io_r_85_b : _GEN_1034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1036 = 7'h56 == r_count_8_io_out ? io_r_86_b : _GEN_1035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1037 = 7'h57 == r_count_8_io_out ? io_r_87_b : _GEN_1036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1038 = 7'h58 == r_count_8_io_out ? io_r_88_b : _GEN_1037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1039 = 7'h59 == r_count_8_io_out ? io_r_89_b : _GEN_1038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1040 = 7'h5a == r_count_8_io_out ? io_r_90_b : _GEN_1039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1041 = 7'h5b == r_count_8_io_out ? io_r_91_b : _GEN_1040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1042 = 7'h5c == r_count_8_io_out ? io_r_92_b : _GEN_1041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1043 = 7'h5d == r_count_8_io_out ? io_r_93_b : _GEN_1042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1044 = 7'h5e == r_count_8_io_out ? io_r_94_b : _GEN_1043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1045 = 7'h5f == r_count_8_io_out ? io_r_95_b : _GEN_1044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1046 = 7'h60 == r_count_8_io_out ? io_r_96_b : _GEN_1045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1047 = 7'h61 == r_count_8_io_out ? io_r_97_b : _GEN_1046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1048 = 7'h62 == r_count_8_io_out ? io_r_98_b : _GEN_1047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1051 = 7'h1 == r_count_9_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1052 = 7'h2 == r_count_9_io_out ? io_r_2_b : _GEN_1051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1053 = 7'h3 == r_count_9_io_out ? io_r_3_b : _GEN_1052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1054 = 7'h4 == r_count_9_io_out ? io_r_4_b : _GEN_1053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1055 = 7'h5 == r_count_9_io_out ? io_r_5_b : _GEN_1054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1056 = 7'h6 == r_count_9_io_out ? io_r_6_b : _GEN_1055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1057 = 7'h7 == r_count_9_io_out ? io_r_7_b : _GEN_1056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1058 = 7'h8 == r_count_9_io_out ? io_r_8_b : _GEN_1057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1059 = 7'h9 == r_count_9_io_out ? io_r_9_b : _GEN_1058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1060 = 7'ha == r_count_9_io_out ? io_r_10_b : _GEN_1059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1061 = 7'hb == r_count_9_io_out ? io_r_11_b : _GEN_1060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1062 = 7'hc == r_count_9_io_out ? io_r_12_b : _GEN_1061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1063 = 7'hd == r_count_9_io_out ? io_r_13_b : _GEN_1062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1064 = 7'he == r_count_9_io_out ? io_r_14_b : _GEN_1063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1065 = 7'hf == r_count_9_io_out ? io_r_15_b : _GEN_1064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1066 = 7'h10 == r_count_9_io_out ? io_r_16_b : _GEN_1065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1067 = 7'h11 == r_count_9_io_out ? io_r_17_b : _GEN_1066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1068 = 7'h12 == r_count_9_io_out ? io_r_18_b : _GEN_1067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1069 = 7'h13 == r_count_9_io_out ? io_r_19_b : _GEN_1068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1070 = 7'h14 == r_count_9_io_out ? io_r_20_b : _GEN_1069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1071 = 7'h15 == r_count_9_io_out ? io_r_21_b : _GEN_1070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1072 = 7'h16 == r_count_9_io_out ? io_r_22_b : _GEN_1071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1073 = 7'h17 == r_count_9_io_out ? io_r_23_b : _GEN_1072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1074 = 7'h18 == r_count_9_io_out ? io_r_24_b : _GEN_1073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1075 = 7'h19 == r_count_9_io_out ? io_r_25_b : _GEN_1074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1076 = 7'h1a == r_count_9_io_out ? io_r_26_b : _GEN_1075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1077 = 7'h1b == r_count_9_io_out ? io_r_27_b : _GEN_1076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1078 = 7'h1c == r_count_9_io_out ? io_r_28_b : _GEN_1077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1079 = 7'h1d == r_count_9_io_out ? io_r_29_b : _GEN_1078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1080 = 7'h1e == r_count_9_io_out ? io_r_30_b : _GEN_1079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1081 = 7'h1f == r_count_9_io_out ? io_r_31_b : _GEN_1080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1082 = 7'h20 == r_count_9_io_out ? io_r_32_b : _GEN_1081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1083 = 7'h21 == r_count_9_io_out ? io_r_33_b : _GEN_1082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1084 = 7'h22 == r_count_9_io_out ? io_r_34_b : _GEN_1083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1085 = 7'h23 == r_count_9_io_out ? io_r_35_b : _GEN_1084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1086 = 7'h24 == r_count_9_io_out ? io_r_36_b : _GEN_1085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1087 = 7'h25 == r_count_9_io_out ? io_r_37_b : _GEN_1086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1088 = 7'h26 == r_count_9_io_out ? io_r_38_b : _GEN_1087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1089 = 7'h27 == r_count_9_io_out ? io_r_39_b : _GEN_1088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1090 = 7'h28 == r_count_9_io_out ? io_r_40_b : _GEN_1089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1091 = 7'h29 == r_count_9_io_out ? io_r_41_b : _GEN_1090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1092 = 7'h2a == r_count_9_io_out ? io_r_42_b : _GEN_1091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1093 = 7'h2b == r_count_9_io_out ? io_r_43_b : _GEN_1092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1094 = 7'h2c == r_count_9_io_out ? io_r_44_b : _GEN_1093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1095 = 7'h2d == r_count_9_io_out ? io_r_45_b : _GEN_1094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1096 = 7'h2e == r_count_9_io_out ? io_r_46_b : _GEN_1095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1097 = 7'h2f == r_count_9_io_out ? io_r_47_b : _GEN_1096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1098 = 7'h30 == r_count_9_io_out ? io_r_48_b : _GEN_1097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1099 = 7'h31 == r_count_9_io_out ? io_r_49_b : _GEN_1098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1100 = 7'h32 == r_count_9_io_out ? io_r_50_b : _GEN_1099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1101 = 7'h33 == r_count_9_io_out ? io_r_51_b : _GEN_1100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1102 = 7'h34 == r_count_9_io_out ? io_r_52_b : _GEN_1101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1103 = 7'h35 == r_count_9_io_out ? io_r_53_b : _GEN_1102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1104 = 7'h36 == r_count_9_io_out ? io_r_54_b : _GEN_1103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1105 = 7'h37 == r_count_9_io_out ? io_r_55_b : _GEN_1104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1106 = 7'h38 == r_count_9_io_out ? io_r_56_b : _GEN_1105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1107 = 7'h39 == r_count_9_io_out ? io_r_57_b : _GEN_1106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1108 = 7'h3a == r_count_9_io_out ? io_r_58_b : _GEN_1107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1109 = 7'h3b == r_count_9_io_out ? io_r_59_b : _GEN_1108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1110 = 7'h3c == r_count_9_io_out ? io_r_60_b : _GEN_1109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1111 = 7'h3d == r_count_9_io_out ? io_r_61_b : _GEN_1110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1112 = 7'h3e == r_count_9_io_out ? io_r_62_b : _GEN_1111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1113 = 7'h3f == r_count_9_io_out ? io_r_63_b : _GEN_1112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1114 = 7'h40 == r_count_9_io_out ? io_r_64_b : _GEN_1113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1115 = 7'h41 == r_count_9_io_out ? io_r_65_b : _GEN_1114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1116 = 7'h42 == r_count_9_io_out ? io_r_66_b : _GEN_1115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1117 = 7'h43 == r_count_9_io_out ? io_r_67_b : _GEN_1116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1118 = 7'h44 == r_count_9_io_out ? io_r_68_b : _GEN_1117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1119 = 7'h45 == r_count_9_io_out ? io_r_69_b : _GEN_1118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1120 = 7'h46 == r_count_9_io_out ? io_r_70_b : _GEN_1119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1121 = 7'h47 == r_count_9_io_out ? io_r_71_b : _GEN_1120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1122 = 7'h48 == r_count_9_io_out ? io_r_72_b : _GEN_1121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1123 = 7'h49 == r_count_9_io_out ? io_r_73_b : _GEN_1122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1124 = 7'h4a == r_count_9_io_out ? io_r_74_b : _GEN_1123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1125 = 7'h4b == r_count_9_io_out ? io_r_75_b : _GEN_1124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1126 = 7'h4c == r_count_9_io_out ? io_r_76_b : _GEN_1125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1127 = 7'h4d == r_count_9_io_out ? io_r_77_b : _GEN_1126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1128 = 7'h4e == r_count_9_io_out ? io_r_78_b : _GEN_1127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1129 = 7'h4f == r_count_9_io_out ? io_r_79_b : _GEN_1128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1130 = 7'h50 == r_count_9_io_out ? io_r_80_b : _GEN_1129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1131 = 7'h51 == r_count_9_io_out ? io_r_81_b : _GEN_1130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1132 = 7'h52 == r_count_9_io_out ? io_r_82_b : _GEN_1131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1133 = 7'h53 == r_count_9_io_out ? io_r_83_b : _GEN_1132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1134 = 7'h54 == r_count_9_io_out ? io_r_84_b : _GEN_1133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1135 = 7'h55 == r_count_9_io_out ? io_r_85_b : _GEN_1134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1136 = 7'h56 == r_count_9_io_out ? io_r_86_b : _GEN_1135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1137 = 7'h57 == r_count_9_io_out ? io_r_87_b : _GEN_1136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1138 = 7'h58 == r_count_9_io_out ? io_r_88_b : _GEN_1137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1139 = 7'h59 == r_count_9_io_out ? io_r_89_b : _GEN_1138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1140 = 7'h5a == r_count_9_io_out ? io_r_90_b : _GEN_1139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1141 = 7'h5b == r_count_9_io_out ? io_r_91_b : _GEN_1140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1142 = 7'h5c == r_count_9_io_out ? io_r_92_b : _GEN_1141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1143 = 7'h5d == r_count_9_io_out ? io_r_93_b : _GEN_1142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1144 = 7'h5e == r_count_9_io_out ? io_r_94_b : _GEN_1143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1145 = 7'h5f == r_count_9_io_out ? io_r_95_b : _GEN_1144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1146 = 7'h60 == r_count_9_io_out ? io_r_96_b : _GEN_1145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1147 = 7'h61 == r_count_9_io_out ? io_r_97_b : _GEN_1146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1148 = 7'h62 == r_count_9_io_out ? io_r_98_b : _GEN_1147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1151 = 7'h1 == r_count_10_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1152 = 7'h2 == r_count_10_io_out ? io_r_2_b : _GEN_1151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1153 = 7'h3 == r_count_10_io_out ? io_r_3_b : _GEN_1152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1154 = 7'h4 == r_count_10_io_out ? io_r_4_b : _GEN_1153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1155 = 7'h5 == r_count_10_io_out ? io_r_5_b : _GEN_1154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1156 = 7'h6 == r_count_10_io_out ? io_r_6_b : _GEN_1155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1157 = 7'h7 == r_count_10_io_out ? io_r_7_b : _GEN_1156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1158 = 7'h8 == r_count_10_io_out ? io_r_8_b : _GEN_1157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1159 = 7'h9 == r_count_10_io_out ? io_r_9_b : _GEN_1158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1160 = 7'ha == r_count_10_io_out ? io_r_10_b : _GEN_1159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1161 = 7'hb == r_count_10_io_out ? io_r_11_b : _GEN_1160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1162 = 7'hc == r_count_10_io_out ? io_r_12_b : _GEN_1161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1163 = 7'hd == r_count_10_io_out ? io_r_13_b : _GEN_1162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1164 = 7'he == r_count_10_io_out ? io_r_14_b : _GEN_1163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1165 = 7'hf == r_count_10_io_out ? io_r_15_b : _GEN_1164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1166 = 7'h10 == r_count_10_io_out ? io_r_16_b : _GEN_1165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1167 = 7'h11 == r_count_10_io_out ? io_r_17_b : _GEN_1166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1168 = 7'h12 == r_count_10_io_out ? io_r_18_b : _GEN_1167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1169 = 7'h13 == r_count_10_io_out ? io_r_19_b : _GEN_1168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1170 = 7'h14 == r_count_10_io_out ? io_r_20_b : _GEN_1169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1171 = 7'h15 == r_count_10_io_out ? io_r_21_b : _GEN_1170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1172 = 7'h16 == r_count_10_io_out ? io_r_22_b : _GEN_1171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1173 = 7'h17 == r_count_10_io_out ? io_r_23_b : _GEN_1172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1174 = 7'h18 == r_count_10_io_out ? io_r_24_b : _GEN_1173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1175 = 7'h19 == r_count_10_io_out ? io_r_25_b : _GEN_1174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1176 = 7'h1a == r_count_10_io_out ? io_r_26_b : _GEN_1175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1177 = 7'h1b == r_count_10_io_out ? io_r_27_b : _GEN_1176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1178 = 7'h1c == r_count_10_io_out ? io_r_28_b : _GEN_1177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1179 = 7'h1d == r_count_10_io_out ? io_r_29_b : _GEN_1178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1180 = 7'h1e == r_count_10_io_out ? io_r_30_b : _GEN_1179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1181 = 7'h1f == r_count_10_io_out ? io_r_31_b : _GEN_1180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1182 = 7'h20 == r_count_10_io_out ? io_r_32_b : _GEN_1181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1183 = 7'h21 == r_count_10_io_out ? io_r_33_b : _GEN_1182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1184 = 7'h22 == r_count_10_io_out ? io_r_34_b : _GEN_1183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1185 = 7'h23 == r_count_10_io_out ? io_r_35_b : _GEN_1184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1186 = 7'h24 == r_count_10_io_out ? io_r_36_b : _GEN_1185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1187 = 7'h25 == r_count_10_io_out ? io_r_37_b : _GEN_1186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1188 = 7'h26 == r_count_10_io_out ? io_r_38_b : _GEN_1187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1189 = 7'h27 == r_count_10_io_out ? io_r_39_b : _GEN_1188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1190 = 7'h28 == r_count_10_io_out ? io_r_40_b : _GEN_1189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1191 = 7'h29 == r_count_10_io_out ? io_r_41_b : _GEN_1190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1192 = 7'h2a == r_count_10_io_out ? io_r_42_b : _GEN_1191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1193 = 7'h2b == r_count_10_io_out ? io_r_43_b : _GEN_1192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1194 = 7'h2c == r_count_10_io_out ? io_r_44_b : _GEN_1193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1195 = 7'h2d == r_count_10_io_out ? io_r_45_b : _GEN_1194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1196 = 7'h2e == r_count_10_io_out ? io_r_46_b : _GEN_1195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1197 = 7'h2f == r_count_10_io_out ? io_r_47_b : _GEN_1196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1198 = 7'h30 == r_count_10_io_out ? io_r_48_b : _GEN_1197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1199 = 7'h31 == r_count_10_io_out ? io_r_49_b : _GEN_1198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1200 = 7'h32 == r_count_10_io_out ? io_r_50_b : _GEN_1199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1201 = 7'h33 == r_count_10_io_out ? io_r_51_b : _GEN_1200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1202 = 7'h34 == r_count_10_io_out ? io_r_52_b : _GEN_1201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1203 = 7'h35 == r_count_10_io_out ? io_r_53_b : _GEN_1202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1204 = 7'h36 == r_count_10_io_out ? io_r_54_b : _GEN_1203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1205 = 7'h37 == r_count_10_io_out ? io_r_55_b : _GEN_1204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1206 = 7'h38 == r_count_10_io_out ? io_r_56_b : _GEN_1205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1207 = 7'h39 == r_count_10_io_out ? io_r_57_b : _GEN_1206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1208 = 7'h3a == r_count_10_io_out ? io_r_58_b : _GEN_1207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1209 = 7'h3b == r_count_10_io_out ? io_r_59_b : _GEN_1208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1210 = 7'h3c == r_count_10_io_out ? io_r_60_b : _GEN_1209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1211 = 7'h3d == r_count_10_io_out ? io_r_61_b : _GEN_1210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1212 = 7'h3e == r_count_10_io_out ? io_r_62_b : _GEN_1211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1213 = 7'h3f == r_count_10_io_out ? io_r_63_b : _GEN_1212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1214 = 7'h40 == r_count_10_io_out ? io_r_64_b : _GEN_1213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1215 = 7'h41 == r_count_10_io_out ? io_r_65_b : _GEN_1214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1216 = 7'h42 == r_count_10_io_out ? io_r_66_b : _GEN_1215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1217 = 7'h43 == r_count_10_io_out ? io_r_67_b : _GEN_1216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1218 = 7'h44 == r_count_10_io_out ? io_r_68_b : _GEN_1217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1219 = 7'h45 == r_count_10_io_out ? io_r_69_b : _GEN_1218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1220 = 7'h46 == r_count_10_io_out ? io_r_70_b : _GEN_1219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1221 = 7'h47 == r_count_10_io_out ? io_r_71_b : _GEN_1220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1222 = 7'h48 == r_count_10_io_out ? io_r_72_b : _GEN_1221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1223 = 7'h49 == r_count_10_io_out ? io_r_73_b : _GEN_1222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1224 = 7'h4a == r_count_10_io_out ? io_r_74_b : _GEN_1223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1225 = 7'h4b == r_count_10_io_out ? io_r_75_b : _GEN_1224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1226 = 7'h4c == r_count_10_io_out ? io_r_76_b : _GEN_1225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1227 = 7'h4d == r_count_10_io_out ? io_r_77_b : _GEN_1226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1228 = 7'h4e == r_count_10_io_out ? io_r_78_b : _GEN_1227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1229 = 7'h4f == r_count_10_io_out ? io_r_79_b : _GEN_1228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1230 = 7'h50 == r_count_10_io_out ? io_r_80_b : _GEN_1229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1231 = 7'h51 == r_count_10_io_out ? io_r_81_b : _GEN_1230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1232 = 7'h52 == r_count_10_io_out ? io_r_82_b : _GEN_1231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1233 = 7'h53 == r_count_10_io_out ? io_r_83_b : _GEN_1232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1234 = 7'h54 == r_count_10_io_out ? io_r_84_b : _GEN_1233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1235 = 7'h55 == r_count_10_io_out ? io_r_85_b : _GEN_1234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1236 = 7'h56 == r_count_10_io_out ? io_r_86_b : _GEN_1235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1237 = 7'h57 == r_count_10_io_out ? io_r_87_b : _GEN_1236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1238 = 7'h58 == r_count_10_io_out ? io_r_88_b : _GEN_1237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1239 = 7'h59 == r_count_10_io_out ? io_r_89_b : _GEN_1238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1240 = 7'h5a == r_count_10_io_out ? io_r_90_b : _GEN_1239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1241 = 7'h5b == r_count_10_io_out ? io_r_91_b : _GEN_1240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1242 = 7'h5c == r_count_10_io_out ? io_r_92_b : _GEN_1241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1243 = 7'h5d == r_count_10_io_out ? io_r_93_b : _GEN_1242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1244 = 7'h5e == r_count_10_io_out ? io_r_94_b : _GEN_1243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1245 = 7'h5f == r_count_10_io_out ? io_r_95_b : _GEN_1244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1246 = 7'h60 == r_count_10_io_out ? io_r_96_b : _GEN_1245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1247 = 7'h61 == r_count_10_io_out ? io_r_97_b : _GEN_1246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1248 = 7'h62 == r_count_10_io_out ? io_r_98_b : _GEN_1247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1251 = 7'h1 == r_count_11_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1252 = 7'h2 == r_count_11_io_out ? io_r_2_b : _GEN_1251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1253 = 7'h3 == r_count_11_io_out ? io_r_3_b : _GEN_1252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1254 = 7'h4 == r_count_11_io_out ? io_r_4_b : _GEN_1253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1255 = 7'h5 == r_count_11_io_out ? io_r_5_b : _GEN_1254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1256 = 7'h6 == r_count_11_io_out ? io_r_6_b : _GEN_1255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1257 = 7'h7 == r_count_11_io_out ? io_r_7_b : _GEN_1256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1258 = 7'h8 == r_count_11_io_out ? io_r_8_b : _GEN_1257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1259 = 7'h9 == r_count_11_io_out ? io_r_9_b : _GEN_1258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1260 = 7'ha == r_count_11_io_out ? io_r_10_b : _GEN_1259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1261 = 7'hb == r_count_11_io_out ? io_r_11_b : _GEN_1260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1262 = 7'hc == r_count_11_io_out ? io_r_12_b : _GEN_1261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1263 = 7'hd == r_count_11_io_out ? io_r_13_b : _GEN_1262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1264 = 7'he == r_count_11_io_out ? io_r_14_b : _GEN_1263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1265 = 7'hf == r_count_11_io_out ? io_r_15_b : _GEN_1264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1266 = 7'h10 == r_count_11_io_out ? io_r_16_b : _GEN_1265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1267 = 7'h11 == r_count_11_io_out ? io_r_17_b : _GEN_1266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1268 = 7'h12 == r_count_11_io_out ? io_r_18_b : _GEN_1267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1269 = 7'h13 == r_count_11_io_out ? io_r_19_b : _GEN_1268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1270 = 7'h14 == r_count_11_io_out ? io_r_20_b : _GEN_1269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1271 = 7'h15 == r_count_11_io_out ? io_r_21_b : _GEN_1270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1272 = 7'h16 == r_count_11_io_out ? io_r_22_b : _GEN_1271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1273 = 7'h17 == r_count_11_io_out ? io_r_23_b : _GEN_1272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1274 = 7'h18 == r_count_11_io_out ? io_r_24_b : _GEN_1273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1275 = 7'h19 == r_count_11_io_out ? io_r_25_b : _GEN_1274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1276 = 7'h1a == r_count_11_io_out ? io_r_26_b : _GEN_1275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1277 = 7'h1b == r_count_11_io_out ? io_r_27_b : _GEN_1276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1278 = 7'h1c == r_count_11_io_out ? io_r_28_b : _GEN_1277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1279 = 7'h1d == r_count_11_io_out ? io_r_29_b : _GEN_1278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1280 = 7'h1e == r_count_11_io_out ? io_r_30_b : _GEN_1279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1281 = 7'h1f == r_count_11_io_out ? io_r_31_b : _GEN_1280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1282 = 7'h20 == r_count_11_io_out ? io_r_32_b : _GEN_1281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1283 = 7'h21 == r_count_11_io_out ? io_r_33_b : _GEN_1282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1284 = 7'h22 == r_count_11_io_out ? io_r_34_b : _GEN_1283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1285 = 7'h23 == r_count_11_io_out ? io_r_35_b : _GEN_1284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1286 = 7'h24 == r_count_11_io_out ? io_r_36_b : _GEN_1285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1287 = 7'h25 == r_count_11_io_out ? io_r_37_b : _GEN_1286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1288 = 7'h26 == r_count_11_io_out ? io_r_38_b : _GEN_1287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1289 = 7'h27 == r_count_11_io_out ? io_r_39_b : _GEN_1288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1290 = 7'h28 == r_count_11_io_out ? io_r_40_b : _GEN_1289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1291 = 7'h29 == r_count_11_io_out ? io_r_41_b : _GEN_1290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1292 = 7'h2a == r_count_11_io_out ? io_r_42_b : _GEN_1291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1293 = 7'h2b == r_count_11_io_out ? io_r_43_b : _GEN_1292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1294 = 7'h2c == r_count_11_io_out ? io_r_44_b : _GEN_1293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1295 = 7'h2d == r_count_11_io_out ? io_r_45_b : _GEN_1294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1296 = 7'h2e == r_count_11_io_out ? io_r_46_b : _GEN_1295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1297 = 7'h2f == r_count_11_io_out ? io_r_47_b : _GEN_1296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1298 = 7'h30 == r_count_11_io_out ? io_r_48_b : _GEN_1297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1299 = 7'h31 == r_count_11_io_out ? io_r_49_b : _GEN_1298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1300 = 7'h32 == r_count_11_io_out ? io_r_50_b : _GEN_1299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1301 = 7'h33 == r_count_11_io_out ? io_r_51_b : _GEN_1300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1302 = 7'h34 == r_count_11_io_out ? io_r_52_b : _GEN_1301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1303 = 7'h35 == r_count_11_io_out ? io_r_53_b : _GEN_1302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1304 = 7'h36 == r_count_11_io_out ? io_r_54_b : _GEN_1303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1305 = 7'h37 == r_count_11_io_out ? io_r_55_b : _GEN_1304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1306 = 7'h38 == r_count_11_io_out ? io_r_56_b : _GEN_1305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1307 = 7'h39 == r_count_11_io_out ? io_r_57_b : _GEN_1306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1308 = 7'h3a == r_count_11_io_out ? io_r_58_b : _GEN_1307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1309 = 7'h3b == r_count_11_io_out ? io_r_59_b : _GEN_1308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1310 = 7'h3c == r_count_11_io_out ? io_r_60_b : _GEN_1309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1311 = 7'h3d == r_count_11_io_out ? io_r_61_b : _GEN_1310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1312 = 7'h3e == r_count_11_io_out ? io_r_62_b : _GEN_1311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1313 = 7'h3f == r_count_11_io_out ? io_r_63_b : _GEN_1312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1314 = 7'h40 == r_count_11_io_out ? io_r_64_b : _GEN_1313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1315 = 7'h41 == r_count_11_io_out ? io_r_65_b : _GEN_1314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1316 = 7'h42 == r_count_11_io_out ? io_r_66_b : _GEN_1315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1317 = 7'h43 == r_count_11_io_out ? io_r_67_b : _GEN_1316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1318 = 7'h44 == r_count_11_io_out ? io_r_68_b : _GEN_1317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1319 = 7'h45 == r_count_11_io_out ? io_r_69_b : _GEN_1318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1320 = 7'h46 == r_count_11_io_out ? io_r_70_b : _GEN_1319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1321 = 7'h47 == r_count_11_io_out ? io_r_71_b : _GEN_1320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1322 = 7'h48 == r_count_11_io_out ? io_r_72_b : _GEN_1321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1323 = 7'h49 == r_count_11_io_out ? io_r_73_b : _GEN_1322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1324 = 7'h4a == r_count_11_io_out ? io_r_74_b : _GEN_1323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1325 = 7'h4b == r_count_11_io_out ? io_r_75_b : _GEN_1324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1326 = 7'h4c == r_count_11_io_out ? io_r_76_b : _GEN_1325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1327 = 7'h4d == r_count_11_io_out ? io_r_77_b : _GEN_1326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1328 = 7'h4e == r_count_11_io_out ? io_r_78_b : _GEN_1327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1329 = 7'h4f == r_count_11_io_out ? io_r_79_b : _GEN_1328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1330 = 7'h50 == r_count_11_io_out ? io_r_80_b : _GEN_1329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1331 = 7'h51 == r_count_11_io_out ? io_r_81_b : _GEN_1330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1332 = 7'h52 == r_count_11_io_out ? io_r_82_b : _GEN_1331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1333 = 7'h53 == r_count_11_io_out ? io_r_83_b : _GEN_1332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1334 = 7'h54 == r_count_11_io_out ? io_r_84_b : _GEN_1333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1335 = 7'h55 == r_count_11_io_out ? io_r_85_b : _GEN_1334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1336 = 7'h56 == r_count_11_io_out ? io_r_86_b : _GEN_1335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1337 = 7'h57 == r_count_11_io_out ? io_r_87_b : _GEN_1336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1338 = 7'h58 == r_count_11_io_out ? io_r_88_b : _GEN_1337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1339 = 7'h59 == r_count_11_io_out ? io_r_89_b : _GEN_1338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1340 = 7'h5a == r_count_11_io_out ? io_r_90_b : _GEN_1339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1341 = 7'h5b == r_count_11_io_out ? io_r_91_b : _GEN_1340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1342 = 7'h5c == r_count_11_io_out ? io_r_92_b : _GEN_1341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1343 = 7'h5d == r_count_11_io_out ? io_r_93_b : _GEN_1342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1344 = 7'h5e == r_count_11_io_out ? io_r_94_b : _GEN_1343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1345 = 7'h5f == r_count_11_io_out ? io_r_95_b : _GEN_1344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1346 = 7'h60 == r_count_11_io_out ? io_r_96_b : _GEN_1345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1347 = 7'h61 == r_count_11_io_out ? io_r_97_b : _GEN_1346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1348 = 7'h62 == r_count_11_io_out ? io_r_98_b : _GEN_1347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1351 = 7'h1 == r_count_12_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1352 = 7'h2 == r_count_12_io_out ? io_r_2_b : _GEN_1351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1353 = 7'h3 == r_count_12_io_out ? io_r_3_b : _GEN_1352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1354 = 7'h4 == r_count_12_io_out ? io_r_4_b : _GEN_1353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1355 = 7'h5 == r_count_12_io_out ? io_r_5_b : _GEN_1354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1356 = 7'h6 == r_count_12_io_out ? io_r_6_b : _GEN_1355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1357 = 7'h7 == r_count_12_io_out ? io_r_7_b : _GEN_1356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1358 = 7'h8 == r_count_12_io_out ? io_r_8_b : _GEN_1357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1359 = 7'h9 == r_count_12_io_out ? io_r_9_b : _GEN_1358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1360 = 7'ha == r_count_12_io_out ? io_r_10_b : _GEN_1359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1361 = 7'hb == r_count_12_io_out ? io_r_11_b : _GEN_1360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1362 = 7'hc == r_count_12_io_out ? io_r_12_b : _GEN_1361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1363 = 7'hd == r_count_12_io_out ? io_r_13_b : _GEN_1362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1364 = 7'he == r_count_12_io_out ? io_r_14_b : _GEN_1363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1365 = 7'hf == r_count_12_io_out ? io_r_15_b : _GEN_1364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1366 = 7'h10 == r_count_12_io_out ? io_r_16_b : _GEN_1365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1367 = 7'h11 == r_count_12_io_out ? io_r_17_b : _GEN_1366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1368 = 7'h12 == r_count_12_io_out ? io_r_18_b : _GEN_1367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1369 = 7'h13 == r_count_12_io_out ? io_r_19_b : _GEN_1368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1370 = 7'h14 == r_count_12_io_out ? io_r_20_b : _GEN_1369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1371 = 7'h15 == r_count_12_io_out ? io_r_21_b : _GEN_1370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1372 = 7'h16 == r_count_12_io_out ? io_r_22_b : _GEN_1371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1373 = 7'h17 == r_count_12_io_out ? io_r_23_b : _GEN_1372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1374 = 7'h18 == r_count_12_io_out ? io_r_24_b : _GEN_1373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1375 = 7'h19 == r_count_12_io_out ? io_r_25_b : _GEN_1374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1376 = 7'h1a == r_count_12_io_out ? io_r_26_b : _GEN_1375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1377 = 7'h1b == r_count_12_io_out ? io_r_27_b : _GEN_1376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1378 = 7'h1c == r_count_12_io_out ? io_r_28_b : _GEN_1377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1379 = 7'h1d == r_count_12_io_out ? io_r_29_b : _GEN_1378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1380 = 7'h1e == r_count_12_io_out ? io_r_30_b : _GEN_1379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1381 = 7'h1f == r_count_12_io_out ? io_r_31_b : _GEN_1380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1382 = 7'h20 == r_count_12_io_out ? io_r_32_b : _GEN_1381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1383 = 7'h21 == r_count_12_io_out ? io_r_33_b : _GEN_1382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1384 = 7'h22 == r_count_12_io_out ? io_r_34_b : _GEN_1383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1385 = 7'h23 == r_count_12_io_out ? io_r_35_b : _GEN_1384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1386 = 7'h24 == r_count_12_io_out ? io_r_36_b : _GEN_1385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1387 = 7'h25 == r_count_12_io_out ? io_r_37_b : _GEN_1386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1388 = 7'h26 == r_count_12_io_out ? io_r_38_b : _GEN_1387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1389 = 7'h27 == r_count_12_io_out ? io_r_39_b : _GEN_1388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1390 = 7'h28 == r_count_12_io_out ? io_r_40_b : _GEN_1389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1391 = 7'h29 == r_count_12_io_out ? io_r_41_b : _GEN_1390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1392 = 7'h2a == r_count_12_io_out ? io_r_42_b : _GEN_1391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1393 = 7'h2b == r_count_12_io_out ? io_r_43_b : _GEN_1392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1394 = 7'h2c == r_count_12_io_out ? io_r_44_b : _GEN_1393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1395 = 7'h2d == r_count_12_io_out ? io_r_45_b : _GEN_1394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1396 = 7'h2e == r_count_12_io_out ? io_r_46_b : _GEN_1395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1397 = 7'h2f == r_count_12_io_out ? io_r_47_b : _GEN_1396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1398 = 7'h30 == r_count_12_io_out ? io_r_48_b : _GEN_1397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1399 = 7'h31 == r_count_12_io_out ? io_r_49_b : _GEN_1398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1400 = 7'h32 == r_count_12_io_out ? io_r_50_b : _GEN_1399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1401 = 7'h33 == r_count_12_io_out ? io_r_51_b : _GEN_1400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1402 = 7'h34 == r_count_12_io_out ? io_r_52_b : _GEN_1401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1403 = 7'h35 == r_count_12_io_out ? io_r_53_b : _GEN_1402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1404 = 7'h36 == r_count_12_io_out ? io_r_54_b : _GEN_1403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1405 = 7'h37 == r_count_12_io_out ? io_r_55_b : _GEN_1404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1406 = 7'h38 == r_count_12_io_out ? io_r_56_b : _GEN_1405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1407 = 7'h39 == r_count_12_io_out ? io_r_57_b : _GEN_1406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1408 = 7'h3a == r_count_12_io_out ? io_r_58_b : _GEN_1407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1409 = 7'h3b == r_count_12_io_out ? io_r_59_b : _GEN_1408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1410 = 7'h3c == r_count_12_io_out ? io_r_60_b : _GEN_1409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1411 = 7'h3d == r_count_12_io_out ? io_r_61_b : _GEN_1410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1412 = 7'h3e == r_count_12_io_out ? io_r_62_b : _GEN_1411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1413 = 7'h3f == r_count_12_io_out ? io_r_63_b : _GEN_1412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1414 = 7'h40 == r_count_12_io_out ? io_r_64_b : _GEN_1413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1415 = 7'h41 == r_count_12_io_out ? io_r_65_b : _GEN_1414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1416 = 7'h42 == r_count_12_io_out ? io_r_66_b : _GEN_1415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1417 = 7'h43 == r_count_12_io_out ? io_r_67_b : _GEN_1416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1418 = 7'h44 == r_count_12_io_out ? io_r_68_b : _GEN_1417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1419 = 7'h45 == r_count_12_io_out ? io_r_69_b : _GEN_1418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1420 = 7'h46 == r_count_12_io_out ? io_r_70_b : _GEN_1419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1421 = 7'h47 == r_count_12_io_out ? io_r_71_b : _GEN_1420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1422 = 7'h48 == r_count_12_io_out ? io_r_72_b : _GEN_1421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1423 = 7'h49 == r_count_12_io_out ? io_r_73_b : _GEN_1422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1424 = 7'h4a == r_count_12_io_out ? io_r_74_b : _GEN_1423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1425 = 7'h4b == r_count_12_io_out ? io_r_75_b : _GEN_1424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1426 = 7'h4c == r_count_12_io_out ? io_r_76_b : _GEN_1425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1427 = 7'h4d == r_count_12_io_out ? io_r_77_b : _GEN_1426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1428 = 7'h4e == r_count_12_io_out ? io_r_78_b : _GEN_1427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1429 = 7'h4f == r_count_12_io_out ? io_r_79_b : _GEN_1428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1430 = 7'h50 == r_count_12_io_out ? io_r_80_b : _GEN_1429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1431 = 7'h51 == r_count_12_io_out ? io_r_81_b : _GEN_1430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1432 = 7'h52 == r_count_12_io_out ? io_r_82_b : _GEN_1431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1433 = 7'h53 == r_count_12_io_out ? io_r_83_b : _GEN_1432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1434 = 7'h54 == r_count_12_io_out ? io_r_84_b : _GEN_1433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1435 = 7'h55 == r_count_12_io_out ? io_r_85_b : _GEN_1434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1436 = 7'h56 == r_count_12_io_out ? io_r_86_b : _GEN_1435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1437 = 7'h57 == r_count_12_io_out ? io_r_87_b : _GEN_1436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1438 = 7'h58 == r_count_12_io_out ? io_r_88_b : _GEN_1437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1439 = 7'h59 == r_count_12_io_out ? io_r_89_b : _GEN_1438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1440 = 7'h5a == r_count_12_io_out ? io_r_90_b : _GEN_1439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1441 = 7'h5b == r_count_12_io_out ? io_r_91_b : _GEN_1440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1442 = 7'h5c == r_count_12_io_out ? io_r_92_b : _GEN_1441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1443 = 7'h5d == r_count_12_io_out ? io_r_93_b : _GEN_1442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1444 = 7'h5e == r_count_12_io_out ? io_r_94_b : _GEN_1443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1445 = 7'h5f == r_count_12_io_out ? io_r_95_b : _GEN_1444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1446 = 7'h60 == r_count_12_io_out ? io_r_96_b : _GEN_1445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1447 = 7'h61 == r_count_12_io_out ? io_r_97_b : _GEN_1446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1448 = 7'h62 == r_count_12_io_out ? io_r_98_b : _GEN_1447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1451 = 7'h1 == r_count_13_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1452 = 7'h2 == r_count_13_io_out ? io_r_2_b : _GEN_1451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1453 = 7'h3 == r_count_13_io_out ? io_r_3_b : _GEN_1452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1454 = 7'h4 == r_count_13_io_out ? io_r_4_b : _GEN_1453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1455 = 7'h5 == r_count_13_io_out ? io_r_5_b : _GEN_1454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1456 = 7'h6 == r_count_13_io_out ? io_r_6_b : _GEN_1455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1457 = 7'h7 == r_count_13_io_out ? io_r_7_b : _GEN_1456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1458 = 7'h8 == r_count_13_io_out ? io_r_8_b : _GEN_1457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1459 = 7'h9 == r_count_13_io_out ? io_r_9_b : _GEN_1458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1460 = 7'ha == r_count_13_io_out ? io_r_10_b : _GEN_1459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1461 = 7'hb == r_count_13_io_out ? io_r_11_b : _GEN_1460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1462 = 7'hc == r_count_13_io_out ? io_r_12_b : _GEN_1461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1463 = 7'hd == r_count_13_io_out ? io_r_13_b : _GEN_1462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1464 = 7'he == r_count_13_io_out ? io_r_14_b : _GEN_1463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1465 = 7'hf == r_count_13_io_out ? io_r_15_b : _GEN_1464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1466 = 7'h10 == r_count_13_io_out ? io_r_16_b : _GEN_1465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1467 = 7'h11 == r_count_13_io_out ? io_r_17_b : _GEN_1466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1468 = 7'h12 == r_count_13_io_out ? io_r_18_b : _GEN_1467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1469 = 7'h13 == r_count_13_io_out ? io_r_19_b : _GEN_1468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1470 = 7'h14 == r_count_13_io_out ? io_r_20_b : _GEN_1469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1471 = 7'h15 == r_count_13_io_out ? io_r_21_b : _GEN_1470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1472 = 7'h16 == r_count_13_io_out ? io_r_22_b : _GEN_1471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1473 = 7'h17 == r_count_13_io_out ? io_r_23_b : _GEN_1472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1474 = 7'h18 == r_count_13_io_out ? io_r_24_b : _GEN_1473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1475 = 7'h19 == r_count_13_io_out ? io_r_25_b : _GEN_1474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1476 = 7'h1a == r_count_13_io_out ? io_r_26_b : _GEN_1475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1477 = 7'h1b == r_count_13_io_out ? io_r_27_b : _GEN_1476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1478 = 7'h1c == r_count_13_io_out ? io_r_28_b : _GEN_1477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1479 = 7'h1d == r_count_13_io_out ? io_r_29_b : _GEN_1478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1480 = 7'h1e == r_count_13_io_out ? io_r_30_b : _GEN_1479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1481 = 7'h1f == r_count_13_io_out ? io_r_31_b : _GEN_1480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1482 = 7'h20 == r_count_13_io_out ? io_r_32_b : _GEN_1481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1483 = 7'h21 == r_count_13_io_out ? io_r_33_b : _GEN_1482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1484 = 7'h22 == r_count_13_io_out ? io_r_34_b : _GEN_1483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1485 = 7'h23 == r_count_13_io_out ? io_r_35_b : _GEN_1484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1486 = 7'h24 == r_count_13_io_out ? io_r_36_b : _GEN_1485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1487 = 7'h25 == r_count_13_io_out ? io_r_37_b : _GEN_1486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1488 = 7'h26 == r_count_13_io_out ? io_r_38_b : _GEN_1487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1489 = 7'h27 == r_count_13_io_out ? io_r_39_b : _GEN_1488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1490 = 7'h28 == r_count_13_io_out ? io_r_40_b : _GEN_1489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1491 = 7'h29 == r_count_13_io_out ? io_r_41_b : _GEN_1490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1492 = 7'h2a == r_count_13_io_out ? io_r_42_b : _GEN_1491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1493 = 7'h2b == r_count_13_io_out ? io_r_43_b : _GEN_1492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1494 = 7'h2c == r_count_13_io_out ? io_r_44_b : _GEN_1493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1495 = 7'h2d == r_count_13_io_out ? io_r_45_b : _GEN_1494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1496 = 7'h2e == r_count_13_io_out ? io_r_46_b : _GEN_1495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1497 = 7'h2f == r_count_13_io_out ? io_r_47_b : _GEN_1496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1498 = 7'h30 == r_count_13_io_out ? io_r_48_b : _GEN_1497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1499 = 7'h31 == r_count_13_io_out ? io_r_49_b : _GEN_1498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1500 = 7'h32 == r_count_13_io_out ? io_r_50_b : _GEN_1499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1501 = 7'h33 == r_count_13_io_out ? io_r_51_b : _GEN_1500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1502 = 7'h34 == r_count_13_io_out ? io_r_52_b : _GEN_1501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1503 = 7'h35 == r_count_13_io_out ? io_r_53_b : _GEN_1502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1504 = 7'h36 == r_count_13_io_out ? io_r_54_b : _GEN_1503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1505 = 7'h37 == r_count_13_io_out ? io_r_55_b : _GEN_1504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1506 = 7'h38 == r_count_13_io_out ? io_r_56_b : _GEN_1505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1507 = 7'h39 == r_count_13_io_out ? io_r_57_b : _GEN_1506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1508 = 7'h3a == r_count_13_io_out ? io_r_58_b : _GEN_1507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1509 = 7'h3b == r_count_13_io_out ? io_r_59_b : _GEN_1508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1510 = 7'h3c == r_count_13_io_out ? io_r_60_b : _GEN_1509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1511 = 7'h3d == r_count_13_io_out ? io_r_61_b : _GEN_1510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1512 = 7'h3e == r_count_13_io_out ? io_r_62_b : _GEN_1511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1513 = 7'h3f == r_count_13_io_out ? io_r_63_b : _GEN_1512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1514 = 7'h40 == r_count_13_io_out ? io_r_64_b : _GEN_1513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1515 = 7'h41 == r_count_13_io_out ? io_r_65_b : _GEN_1514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1516 = 7'h42 == r_count_13_io_out ? io_r_66_b : _GEN_1515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1517 = 7'h43 == r_count_13_io_out ? io_r_67_b : _GEN_1516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1518 = 7'h44 == r_count_13_io_out ? io_r_68_b : _GEN_1517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1519 = 7'h45 == r_count_13_io_out ? io_r_69_b : _GEN_1518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1520 = 7'h46 == r_count_13_io_out ? io_r_70_b : _GEN_1519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1521 = 7'h47 == r_count_13_io_out ? io_r_71_b : _GEN_1520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1522 = 7'h48 == r_count_13_io_out ? io_r_72_b : _GEN_1521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1523 = 7'h49 == r_count_13_io_out ? io_r_73_b : _GEN_1522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1524 = 7'h4a == r_count_13_io_out ? io_r_74_b : _GEN_1523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1525 = 7'h4b == r_count_13_io_out ? io_r_75_b : _GEN_1524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1526 = 7'h4c == r_count_13_io_out ? io_r_76_b : _GEN_1525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1527 = 7'h4d == r_count_13_io_out ? io_r_77_b : _GEN_1526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1528 = 7'h4e == r_count_13_io_out ? io_r_78_b : _GEN_1527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1529 = 7'h4f == r_count_13_io_out ? io_r_79_b : _GEN_1528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1530 = 7'h50 == r_count_13_io_out ? io_r_80_b : _GEN_1529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1531 = 7'h51 == r_count_13_io_out ? io_r_81_b : _GEN_1530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1532 = 7'h52 == r_count_13_io_out ? io_r_82_b : _GEN_1531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1533 = 7'h53 == r_count_13_io_out ? io_r_83_b : _GEN_1532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1534 = 7'h54 == r_count_13_io_out ? io_r_84_b : _GEN_1533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1535 = 7'h55 == r_count_13_io_out ? io_r_85_b : _GEN_1534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1536 = 7'h56 == r_count_13_io_out ? io_r_86_b : _GEN_1535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1537 = 7'h57 == r_count_13_io_out ? io_r_87_b : _GEN_1536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1538 = 7'h58 == r_count_13_io_out ? io_r_88_b : _GEN_1537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1539 = 7'h59 == r_count_13_io_out ? io_r_89_b : _GEN_1538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1540 = 7'h5a == r_count_13_io_out ? io_r_90_b : _GEN_1539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1541 = 7'h5b == r_count_13_io_out ? io_r_91_b : _GEN_1540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1542 = 7'h5c == r_count_13_io_out ? io_r_92_b : _GEN_1541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1543 = 7'h5d == r_count_13_io_out ? io_r_93_b : _GEN_1542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1544 = 7'h5e == r_count_13_io_out ? io_r_94_b : _GEN_1543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1545 = 7'h5f == r_count_13_io_out ? io_r_95_b : _GEN_1544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1546 = 7'h60 == r_count_13_io_out ? io_r_96_b : _GEN_1545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1547 = 7'h61 == r_count_13_io_out ? io_r_97_b : _GEN_1546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1548 = 7'h62 == r_count_13_io_out ? io_r_98_b : _GEN_1547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1551 = 7'h1 == r_count_14_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1552 = 7'h2 == r_count_14_io_out ? io_r_2_b : _GEN_1551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1553 = 7'h3 == r_count_14_io_out ? io_r_3_b : _GEN_1552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1554 = 7'h4 == r_count_14_io_out ? io_r_4_b : _GEN_1553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1555 = 7'h5 == r_count_14_io_out ? io_r_5_b : _GEN_1554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1556 = 7'h6 == r_count_14_io_out ? io_r_6_b : _GEN_1555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1557 = 7'h7 == r_count_14_io_out ? io_r_7_b : _GEN_1556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1558 = 7'h8 == r_count_14_io_out ? io_r_8_b : _GEN_1557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1559 = 7'h9 == r_count_14_io_out ? io_r_9_b : _GEN_1558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1560 = 7'ha == r_count_14_io_out ? io_r_10_b : _GEN_1559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1561 = 7'hb == r_count_14_io_out ? io_r_11_b : _GEN_1560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1562 = 7'hc == r_count_14_io_out ? io_r_12_b : _GEN_1561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1563 = 7'hd == r_count_14_io_out ? io_r_13_b : _GEN_1562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1564 = 7'he == r_count_14_io_out ? io_r_14_b : _GEN_1563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1565 = 7'hf == r_count_14_io_out ? io_r_15_b : _GEN_1564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1566 = 7'h10 == r_count_14_io_out ? io_r_16_b : _GEN_1565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1567 = 7'h11 == r_count_14_io_out ? io_r_17_b : _GEN_1566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1568 = 7'h12 == r_count_14_io_out ? io_r_18_b : _GEN_1567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1569 = 7'h13 == r_count_14_io_out ? io_r_19_b : _GEN_1568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1570 = 7'h14 == r_count_14_io_out ? io_r_20_b : _GEN_1569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1571 = 7'h15 == r_count_14_io_out ? io_r_21_b : _GEN_1570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1572 = 7'h16 == r_count_14_io_out ? io_r_22_b : _GEN_1571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1573 = 7'h17 == r_count_14_io_out ? io_r_23_b : _GEN_1572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1574 = 7'h18 == r_count_14_io_out ? io_r_24_b : _GEN_1573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1575 = 7'h19 == r_count_14_io_out ? io_r_25_b : _GEN_1574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1576 = 7'h1a == r_count_14_io_out ? io_r_26_b : _GEN_1575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1577 = 7'h1b == r_count_14_io_out ? io_r_27_b : _GEN_1576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1578 = 7'h1c == r_count_14_io_out ? io_r_28_b : _GEN_1577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1579 = 7'h1d == r_count_14_io_out ? io_r_29_b : _GEN_1578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1580 = 7'h1e == r_count_14_io_out ? io_r_30_b : _GEN_1579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1581 = 7'h1f == r_count_14_io_out ? io_r_31_b : _GEN_1580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1582 = 7'h20 == r_count_14_io_out ? io_r_32_b : _GEN_1581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1583 = 7'h21 == r_count_14_io_out ? io_r_33_b : _GEN_1582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1584 = 7'h22 == r_count_14_io_out ? io_r_34_b : _GEN_1583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1585 = 7'h23 == r_count_14_io_out ? io_r_35_b : _GEN_1584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1586 = 7'h24 == r_count_14_io_out ? io_r_36_b : _GEN_1585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1587 = 7'h25 == r_count_14_io_out ? io_r_37_b : _GEN_1586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1588 = 7'h26 == r_count_14_io_out ? io_r_38_b : _GEN_1587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1589 = 7'h27 == r_count_14_io_out ? io_r_39_b : _GEN_1588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1590 = 7'h28 == r_count_14_io_out ? io_r_40_b : _GEN_1589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1591 = 7'h29 == r_count_14_io_out ? io_r_41_b : _GEN_1590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1592 = 7'h2a == r_count_14_io_out ? io_r_42_b : _GEN_1591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1593 = 7'h2b == r_count_14_io_out ? io_r_43_b : _GEN_1592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1594 = 7'h2c == r_count_14_io_out ? io_r_44_b : _GEN_1593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1595 = 7'h2d == r_count_14_io_out ? io_r_45_b : _GEN_1594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1596 = 7'h2e == r_count_14_io_out ? io_r_46_b : _GEN_1595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1597 = 7'h2f == r_count_14_io_out ? io_r_47_b : _GEN_1596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1598 = 7'h30 == r_count_14_io_out ? io_r_48_b : _GEN_1597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1599 = 7'h31 == r_count_14_io_out ? io_r_49_b : _GEN_1598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1600 = 7'h32 == r_count_14_io_out ? io_r_50_b : _GEN_1599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1601 = 7'h33 == r_count_14_io_out ? io_r_51_b : _GEN_1600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1602 = 7'h34 == r_count_14_io_out ? io_r_52_b : _GEN_1601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1603 = 7'h35 == r_count_14_io_out ? io_r_53_b : _GEN_1602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1604 = 7'h36 == r_count_14_io_out ? io_r_54_b : _GEN_1603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1605 = 7'h37 == r_count_14_io_out ? io_r_55_b : _GEN_1604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1606 = 7'h38 == r_count_14_io_out ? io_r_56_b : _GEN_1605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1607 = 7'h39 == r_count_14_io_out ? io_r_57_b : _GEN_1606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1608 = 7'h3a == r_count_14_io_out ? io_r_58_b : _GEN_1607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1609 = 7'h3b == r_count_14_io_out ? io_r_59_b : _GEN_1608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1610 = 7'h3c == r_count_14_io_out ? io_r_60_b : _GEN_1609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1611 = 7'h3d == r_count_14_io_out ? io_r_61_b : _GEN_1610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1612 = 7'h3e == r_count_14_io_out ? io_r_62_b : _GEN_1611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1613 = 7'h3f == r_count_14_io_out ? io_r_63_b : _GEN_1612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1614 = 7'h40 == r_count_14_io_out ? io_r_64_b : _GEN_1613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1615 = 7'h41 == r_count_14_io_out ? io_r_65_b : _GEN_1614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1616 = 7'h42 == r_count_14_io_out ? io_r_66_b : _GEN_1615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1617 = 7'h43 == r_count_14_io_out ? io_r_67_b : _GEN_1616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1618 = 7'h44 == r_count_14_io_out ? io_r_68_b : _GEN_1617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1619 = 7'h45 == r_count_14_io_out ? io_r_69_b : _GEN_1618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1620 = 7'h46 == r_count_14_io_out ? io_r_70_b : _GEN_1619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1621 = 7'h47 == r_count_14_io_out ? io_r_71_b : _GEN_1620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1622 = 7'h48 == r_count_14_io_out ? io_r_72_b : _GEN_1621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1623 = 7'h49 == r_count_14_io_out ? io_r_73_b : _GEN_1622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1624 = 7'h4a == r_count_14_io_out ? io_r_74_b : _GEN_1623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1625 = 7'h4b == r_count_14_io_out ? io_r_75_b : _GEN_1624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1626 = 7'h4c == r_count_14_io_out ? io_r_76_b : _GEN_1625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1627 = 7'h4d == r_count_14_io_out ? io_r_77_b : _GEN_1626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1628 = 7'h4e == r_count_14_io_out ? io_r_78_b : _GEN_1627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1629 = 7'h4f == r_count_14_io_out ? io_r_79_b : _GEN_1628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1630 = 7'h50 == r_count_14_io_out ? io_r_80_b : _GEN_1629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1631 = 7'h51 == r_count_14_io_out ? io_r_81_b : _GEN_1630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1632 = 7'h52 == r_count_14_io_out ? io_r_82_b : _GEN_1631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1633 = 7'h53 == r_count_14_io_out ? io_r_83_b : _GEN_1632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1634 = 7'h54 == r_count_14_io_out ? io_r_84_b : _GEN_1633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1635 = 7'h55 == r_count_14_io_out ? io_r_85_b : _GEN_1634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1636 = 7'h56 == r_count_14_io_out ? io_r_86_b : _GEN_1635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1637 = 7'h57 == r_count_14_io_out ? io_r_87_b : _GEN_1636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1638 = 7'h58 == r_count_14_io_out ? io_r_88_b : _GEN_1637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1639 = 7'h59 == r_count_14_io_out ? io_r_89_b : _GEN_1638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1640 = 7'h5a == r_count_14_io_out ? io_r_90_b : _GEN_1639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1641 = 7'h5b == r_count_14_io_out ? io_r_91_b : _GEN_1640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1642 = 7'h5c == r_count_14_io_out ? io_r_92_b : _GEN_1641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1643 = 7'h5d == r_count_14_io_out ? io_r_93_b : _GEN_1642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1644 = 7'h5e == r_count_14_io_out ? io_r_94_b : _GEN_1643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1645 = 7'h5f == r_count_14_io_out ? io_r_95_b : _GEN_1644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1646 = 7'h60 == r_count_14_io_out ? io_r_96_b : _GEN_1645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1647 = 7'h61 == r_count_14_io_out ? io_r_97_b : _GEN_1646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1648 = 7'h62 == r_count_14_io_out ? io_r_98_b : _GEN_1647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1651 = 7'h1 == r_count_15_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1652 = 7'h2 == r_count_15_io_out ? io_r_2_b : _GEN_1651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1653 = 7'h3 == r_count_15_io_out ? io_r_3_b : _GEN_1652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1654 = 7'h4 == r_count_15_io_out ? io_r_4_b : _GEN_1653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1655 = 7'h5 == r_count_15_io_out ? io_r_5_b : _GEN_1654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1656 = 7'h6 == r_count_15_io_out ? io_r_6_b : _GEN_1655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1657 = 7'h7 == r_count_15_io_out ? io_r_7_b : _GEN_1656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1658 = 7'h8 == r_count_15_io_out ? io_r_8_b : _GEN_1657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1659 = 7'h9 == r_count_15_io_out ? io_r_9_b : _GEN_1658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1660 = 7'ha == r_count_15_io_out ? io_r_10_b : _GEN_1659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1661 = 7'hb == r_count_15_io_out ? io_r_11_b : _GEN_1660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1662 = 7'hc == r_count_15_io_out ? io_r_12_b : _GEN_1661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1663 = 7'hd == r_count_15_io_out ? io_r_13_b : _GEN_1662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1664 = 7'he == r_count_15_io_out ? io_r_14_b : _GEN_1663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1665 = 7'hf == r_count_15_io_out ? io_r_15_b : _GEN_1664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1666 = 7'h10 == r_count_15_io_out ? io_r_16_b : _GEN_1665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1667 = 7'h11 == r_count_15_io_out ? io_r_17_b : _GEN_1666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1668 = 7'h12 == r_count_15_io_out ? io_r_18_b : _GEN_1667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1669 = 7'h13 == r_count_15_io_out ? io_r_19_b : _GEN_1668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1670 = 7'h14 == r_count_15_io_out ? io_r_20_b : _GEN_1669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1671 = 7'h15 == r_count_15_io_out ? io_r_21_b : _GEN_1670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1672 = 7'h16 == r_count_15_io_out ? io_r_22_b : _GEN_1671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1673 = 7'h17 == r_count_15_io_out ? io_r_23_b : _GEN_1672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1674 = 7'h18 == r_count_15_io_out ? io_r_24_b : _GEN_1673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1675 = 7'h19 == r_count_15_io_out ? io_r_25_b : _GEN_1674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1676 = 7'h1a == r_count_15_io_out ? io_r_26_b : _GEN_1675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1677 = 7'h1b == r_count_15_io_out ? io_r_27_b : _GEN_1676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1678 = 7'h1c == r_count_15_io_out ? io_r_28_b : _GEN_1677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1679 = 7'h1d == r_count_15_io_out ? io_r_29_b : _GEN_1678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1680 = 7'h1e == r_count_15_io_out ? io_r_30_b : _GEN_1679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1681 = 7'h1f == r_count_15_io_out ? io_r_31_b : _GEN_1680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1682 = 7'h20 == r_count_15_io_out ? io_r_32_b : _GEN_1681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1683 = 7'h21 == r_count_15_io_out ? io_r_33_b : _GEN_1682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1684 = 7'h22 == r_count_15_io_out ? io_r_34_b : _GEN_1683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1685 = 7'h23 == r_count_15_io_out ? io_r_35_b : _GEN_1684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1686 = 7'h24 == r_count_15_io_out ? io_r_36_b : _GEN_1685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1687 = 7'h25 == r_count_15_io_out ? io_r_37_b : _GEN_1686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1688 = 7'h26 == r_count_15_io_out ? io_r_38_b : _GEN_1687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1689 = 7'h27 == r_count_15_io_out ? io_r_39_b : _GEN_1688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1690 = 7'h28 == r_count_15_io_out ? io_r_40_b : _GEN_1689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1691 = 7'h29 == r_count_15_io_out ? io_r_41_b : _GEN_1690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1692 = 7'h2a == r_count_15_io_out ? io_r_42_b : _GEN_1691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1693 = 7'h2b == r_count_15_io_out ? io_r_43_b : _GEN_1692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1694 = 7'h2c == r_count_15_io_out ? io_r_44_b : _GEN_1693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1695 = 7'h2d == r_count_15_io_out ? io_r_45_b : _GEN_1694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1696 = 7'h2e == r_count_15_io_out ? io_r_46_b : _GEN_1695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1697 = 7'h2f == r_count_15_io_out ? io_r_47_b : _GEN_1696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1698 = 7'h30 == r_count_15_io_out ? io_r_48_b : _GEN_1697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1699 = 7'h31 == r_count_15_io_out ? io_r_49_b : _GEN_1698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1700 = 7'h32 == r_count_15_io_out ? io_r_50_b : _GEN_1699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1701 = 7'h33 == r_count_15_io_out ? io_r_51_b : _GEN_1700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1702 = 7'h34 == r_count_15_io_out ? io_r_52_b : _GEN_1701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1703 = 7'h35 == r_count_15_io_out ? io_r_53_b : _GEN_1702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1704 = 7'h36 == r_count_15_io_out ? io_r_54_b : _GEN_1703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1705 = 7'h37 == r_count_15_io_out ? io_r_55_b : _GEN_1704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1706 = 7'h38 == r_count_15_io_out ? io_r_56_b : _GEN_1705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1707 = 7'h39 == r_count_15_io_out ? io_r_57_b : _GEN_1706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1708 = 7'h3a == r_count_15_io_out ? io_r_58_b : _GEN_1707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1709 = 7'h3b == r_count_15_io_out ? io_r_59_b : _GEN_1708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1710 = 7'h3c == r_count_15_io_out ? io_r_60_b : _GEN_1709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1711 = 7'h3d == r_count_15_io_out ? io_r_61_b : _GEN_1710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1712 = 7'h3e == r_count_15_io_out ? io_r_62_b : _GEN_1711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1713 = 7'h3f == r_count_15_io_out ? io_r_63_b : _GEN_1712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1714 = 7'h40 == r_count_15_io_out ? io_r_64_b : _GEN_1713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1715 = 7'h41 == r_count_15_io_out ? io_r_65_b : _GEN_1714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1716 = 7'h42 == r_count_15_io_out ? io_r_66_b : _GEN_1715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1717 = 7'h43 == r_count_15_io_out ? io_r_67_b : _GEN_1716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1718 = 7'h44 == r_count_15_io_out ? io_r_68_b : _GEN_1717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1719 = 7'h45 == r_count_15_io_out ? io_r_69_b : _GEN_1718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1720 = 7'h46 == r_count_15_io_out ? io_r_70_b : _GEN_1719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1721 = 7'h47 == r_count_15_io_out ? io_r_71_b : _GEN_1720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1722 = 7'h48 == r_count_15_io_out ? io_r_72_b : _GEN_1721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1723 = 7'h49 == r_count_15_io_out ? io_r_73_b : _GEN_1722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1724 = 7'h4a == r_count_15_io_out ? io_r_74_b : _GEN_1723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1725 = 7'h4b == r_count_15_io_out ? io_r_75_b : _GEN_1724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1726 = 7'h4c == r_count_15_io_out ? io_r_76_b : _GEN_1725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1727 = 7'h4d == r_count_15_io_out ? io_r_77_b : _GEN_1726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1728 = 7'h4e == r_count_15_io_out ? io_r_78_b : _GEN_1727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1729 = 7'h4f == r_count_15_io_out ? io_r_79_b : _GEN_1728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1730 = 7'h50 == r_count_15_io_out ? io_r_80_b : _GEN_1729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1731 = 7'h51 == r_count_15_io_out ? io_r_81_b : _GEN_1730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1732 = 7'h52 == r_count_15_io_out ? io_r_82_b : _GEN_1731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1733 = 7'h53 == r_count_15_io_out ? io_r_83_b : _GEN_1732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1734 = 7'h54 == r_count_15_io_out ? io_r_84_b : _GEN_1733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1735 = 7'h55 == r_count_15_io_out ? io_r_85_b : _GEN_1734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1736 = 7'h56 == r_count_15_io_out ? io_r_86_b : _GEN_1735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1737 = 7'h57 == r_count_15_io_out ? io_r_87_b : _GEN_1736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1738 = 7'h58 == r_count_15_io_out ? io_r_88_b : _GEN_1737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1739 = 7'h59 == r_count_15_io_out ? io_r_89_b : _GEN_1738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1740 = 7'h5a == r_count_15_io_out ? io_r_90_b : _GEN_1739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1741 = 7'h5b == r_count_15_io_out ? io_r_91_b : _GEN_1740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1742 = 7'h5c == r_count_15_io_out ? io_r_92_b : _GEN_1741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1743 = 7'h5d == r_count_15_io_out ? io_r_93_b : _GEN_1742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1744 = 7'h5e == r_count_15_io_out ? io_r_94_b : _GEN_1743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1745 = 7'h5f == r_count_15_io_out ? io_r_95_b : _GEN_1744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1746 = 7'h60 == r_count_15_io_out ? io_r_96_b : _GEN_1745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1747 = 7'h61 == r_count_15_io_out ? io_r_97_b : _GEN_1746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1748 = 7'h62 == r_count_15_io_out ? io_r_98_b : _GEN_1747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1751 = 7'h1 == r_count_16_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1752 = 7'h2 == r_count_16_io_out ? io_r_2_b : _GEN_1751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1753 = 7'h3 == r_count_16_io_out ? io_r_3_b : _GEN_1752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1754 = 7'h4 == r_count_16_io_out ? io_r_4_b : _GEN_1753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1755 = 7'h5 == r_count_16_io_out ? io_r_5_b : _GEN_1754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1756 = 7'h6 == r_count_16_io_out ? io_r_6_b : _GEN_1755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1757 = 7'h7 == r_count_16_io_out ? io_r_7_b : _GEN_1756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1758 = 7'h8 == r_count_16_io_out ? io_r_8_b : _GEN_1757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1759 = 7'h9 == r_count_16_io_out ? io_r_9_b : _GEN_1758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1760 = 7'ha == r_count_16_io_out ? io_r_10_b : _GEN_1759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1761 = 7'hb == r_count_16_io_out ? io_r_11_b : _GEN_1760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1762 = 7'hc == r_count_16_io_out ? io_r_12_b : _GEN_1761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1763 = 7'hd == r_count_16_io_out ? io_r_13_b : _GEN_1762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1764 = 7'he == r_count_16_io_out ? io_r_14_b : _GEN_1763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1765 = 7'hf == r_count_16_io_out ? io_r_15_b : _GEN_1764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1766 = 7'h10 == r_count_16_io_out ? io_r_16_b : _GEN_1765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1767 = 7'h11 == r_count_16_io_out ? io_r_17_b : _GEN_1766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1768 = 7'h12 == r_count_16_io_out ? io_r_18_b : _GEN_1767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1769 = 7'h13 == r_count_16_io_out ? io_r_19_b : _GEN_1768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1770 = 7'h14 == r_count_16_io_out ? io_r_20_b : _GEN_1769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1771 = 7'h15 == r_count_16_io_out ? io_r_21_b : _GEN_1770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1772 = 7'h16 == r_count_16_io_out ? io_r_22_b : _GEN_1771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1773 = 7'h17 == r_count_16_io_out ? io_r_23_b : _GEN_1772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1774 = 7'h18 == r_count_16_io_out ? io_r_24_b : _GEN_1773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1775 = 7'h19 == r_count_16_io_out ? io_r_25_b : _GEN_1774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1776 = 7'h1a == r_count_16_io_out ? io_r_26_b : _GEN_1775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1777 = 7'h1b == r_count_16_io_out ? io_r_27_b : _GEN_1776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1778 = 7'h1c == r_count_16_io_out ? io_r_28_b : _GEN_1777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1779 = 7'h1d == r_count_16_io_out ? io_r_29_b : _GEN_1778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1780 = 7'h1e == r_count_16_io_out ? io_r_30_b : _GEN_1779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1781 = 7'h1f == r_count_16_io_out ? io_r_31_b : _GEN_1780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1782 = 7'h20 == r_count_16_io_out ? io_r_32_b : _GEN_1781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1783 = 7'h21 == r_count_16_io_out ? io_r_33_b : _GEN_1782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1784 = 7'h22 == r_count_16_io_out ? io_r_34_b : _GEN_1783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1785 = 7'h23 == r_count_16_io_out ? io_r_35_b : _GEN_1784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1786 = 7'h24 == r_count_16_io_out ? io_r_36_b : _GEN_1785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1787 = 7'h25 == r_count_16_io_out ? io_r_37_b : _GEN_1786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1788 = 7'h26 == r_count_16_io_out ? io_r_38_b : _GEN_1787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1789 = 7'h27 == r_count_16_io_out ? io_r_39_b : _GEN_1788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1790 = 7'h28 == r_count_16_io_out ? io_r_40_b : _GEN_1789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1791 = 7'h29 == r_count_16_io_out ? io_r_41_b : _GEN_1790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1792 = 7'h2a == r_count_16_io_out ? io_r_42_b : _GEN_1791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1793 = 7'h2b == r_count_16_io_out ? io_r_43_b : _GEN_1792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1794 = 7'h2c == r_count_16_io_out ? io_r_44_b : _GEN_1793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1795 = 7'h2d == r_count_16_io_out ? io_r_45_b : _GEN_1794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1796 = 7'h2e == r_count_16_io_out ? io_r_46_b : _GEN_1795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1797 = 7'h2f == r_count_16_io_out ? io_r_47_b : _GEN_1796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1798 = 7'h30 == r_count_16_io_out ? io_r_48_b : _GEN_1797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1799 = 7'h31 == r_count_16_io_out ? io_r_49_b : _GEN_1798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1800 = 7'h32 == r_count_16_io_out ? io_r_50_b : _GEN_1799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1801 = 7'h33 == r_count_16_io_out ? io_r_51_b : _GEN_1800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1802 = 7'h34 == r_count_16_io_out ? io_r_52_b : _GEN_1801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1803 = 7'h35 == r_count_16_io_out ? io_r_53_b : _GEN_1802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1804 = 7'h36 == r_count_16_io_out ? io_r_54_b : _GEN_1803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1805 = 7'h37 == r_count_16_io_out ? io_r_55_b : _GEN_1804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1806 = 7'h38 == r_count_16_io_out ? io_r_56_b : _GEN_1805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1807 = 7'h39 == r_count_16_io_out ? io_r_57_b : _GEN_1806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1808 = 7'h3a == r_count_16_io_out ? io_r_58_b : _GEN_1807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1809 = 7'h3b == r_count_16_io_out ? io_r_59_b : _GEN_1808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1810 = 7'h3c == r_count_16_io_out ? io_r_60_b : _GEN_1809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1811 = 7'h3d == r_count_16_io_out ? io_r_61_b : _GEN_1810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1812 = 7'h3e == r_count_16_io_out ? io_r_62_b : _GEN_1811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1813 = 7'h3f == r_count_16_io_out ? io_r_63_b : _GEN_1812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1814 = 7'h40 == r_count_16_io_out ? io_r_64_b : _GEN_1813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1815 = 7'h41 == r_count_16_io_out ? io_r_65_b : _GEN_1814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1816 = 7'h42 == r_count_16_io_out ? io_r_66_b : _GEN_1815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1817 = 7'h43 == r_count_16_io_out ? io_r_67_b : _GEN_1816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1818 = 7'h44 == r_count_16_io_out ? io_r_68_b : _GEN_1817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1819 = 7'h45 == r_count_16_io_out ? io_r_69_b : _GEN_1818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1820 = 7'h46 == r_count_16_io_out ? io_r_70_b : _GEN_1819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1821 = 7'h47 == r_count_16_io_out ? io_r_71_b : _GEN_1820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1822 = 7'h48 == r_count_16_io_out ? io_r_72_b : _GEN_1821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1823 = 7'h49 == r_count_16_io_out ? io_r_73_b : _GEN_1822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1824 = 7'h4a == r_count_16_io_out ? io_r_74_b : _GEN_1823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1825 = 7'h4b == r_count_16_io_out ? io_r_75_b : _GEN_1824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1826 = 7'h4c == r_count_16_io_out ? io_r_76_b : _GEN_1825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1827 = 7'h4d == r_count_16_io_out ? io_r_77_b : _GEN_1826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1828 = 7'h4e == r_count_16_io_out ? io_r_78_b : _GEN_1827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1829 = 7'h4f == r_count_16_io_out ? io_r_79_b : _GEN_1828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1830 = 7'h50 == r_count_16_io_out ? io_r_80_b : _GEN_1829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1831 = 7'h51 == r_count_16_io_out ? io_r_81_b : _GEN_1830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1832 = 7'h52 == r_count_16_io_out ? io_r_82_b : _GEN_1831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1833 = 7'h53 == r_count_16_io_out ? io_r_83_b : _GEN_1832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1834 = 7'h54 == r_count_16_io_out ? io_r_84_b : _GEN_1833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1835 = 7'h55 == r_count_16_io_out ? io_r_85_b : _GEN_1834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1836 = 7'h56 == r_count_16_io_out ? io_r_86_b : _GEN_1835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1837 = 7'h57 == r_count_16_io_out ? io_r_87_b : _GEN_1836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1838 = 7'h58 == r_count_16_io_out ? io_r_88_b : _GEN_1837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1839 = 7'h59 == r_count_16_io_out ? io_r_89_b : _GEN_1838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1840 = 7'h5a == r_count_16_io_out ? io_r_90_b : _GEN_1839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1841 = 7'h5b == r_count_16_io_out ? io_r_91_b : _GEN_1840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1842 = 7'h5c == r_count_16_io_out ? io_r_92_b : _GEN_1841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1843 = 7'h5d == r_count_16_io_out ? io_r_93_b : _GEN_1842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1844 = 7'h5e == r_count_16_io_out ? io_r_94_b : _GEN_1843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1845 = 7'h5f == r_count_16_io_out ? io_r_95_b : _GEN_1844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1846 = 7'h60 == r_count_16_io_out ? io_r_96_b : _GEN_1845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1847 = 7'h61 == r_count_16_io_out ? io_r_97_b : _GEN_1846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1848 = 7'h62 == r_count_16_io_out ? io_r_98_b : _GEN_1847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1851 = 7'h1 == r_count_17_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1852 = 7'h2 == r_count_17_io_out ? io_r_2_b : _GEN_1851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1853 = 7'h3 == r_count_17_io_out ? io_r_3_b : _GEN_1852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1854 = 7'h4 == r_count_17_io_out ? io_r_4_b : _GEN_1853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1855 = 7'h5 == r_count_17_io_out ? io_r_5_b : _GEN_1854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1856 = 7'h6 == r_count_17_io_out ? io_r_6_b : _GEN_1855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1857 = 7'h7 == r_count_17_io_out ? io_r_7_b : _GEN_1856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1858 = 7'h8 == r_count_17_io_out ? io_r_8_b : _GEN_1857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1859 = 7'h9 == r_count_17_io_out ? io_r_9_b : _GEN_1858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1860 = 7'ha == r_count_17_io_out ? io_r_10_b : _GEN_1859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1861 = 7'hb == r_count_17_io_out ? io_r_11_b : _GEN_1860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1862 = 7'hc == r_count_17_io_out ? io_r_12_b : _GEN_1861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1863 = 7'hd == r_count_17_io_out ? io_r_13_b : _GEN_1862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1864 = 7'he == r_count_17_io_out ? io_r_14_b : _GEN_1863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1865 = 7'hf == r_count_17_io_out ? io_r_15_b : _GEN_1864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1866 = 7'h10 == r_count_17_io_out ? io_r_16_b : _GEN_1865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1867 = 7'h11 == r_count_17_io_out ? io_r_17_b : _GEN_1866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1868 = 7'h12 == r_count_17_io_out ? io_r_18_b : _GEN_1867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1869 = 7'h13 == r_count_17_io_out ? io_r_19_b : _GEN_1868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1870 = 7'h14 == r_count_17_io_out ? io_r_20_b : _GEN_1869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1871 = 7'h15 == r_count_17_io_out ? io_r_21_b : _GEN_1870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1872 = 7'h16 == r_count_17_io_out ? io_r_22_b : _GEN_1871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1873 = 7'h17 == r_count_17_io_out ? io_r_23_b : _GEN_1872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1874 = 7'h18 == r_count_17_io_out ? io_r_24_b : _GEN_1873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1875 = 7'h19 == r_count_17_io_out ? io_r_25_b : _GEN_1874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1876 = 7'h1a == r_count_17_io_out ? io_r_26_b : _GEN_1875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1877 = 7'h1b == r_count_17_io_out ? io_r_27_b : _GEN_1876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1878 = 7'h1c == r_count_17_io_out ? io_r_28_b : _GEN_1877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1879 = 7'h1d == r_count_17_io_out ? io_r_29_b : _GEN_1878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1880 = 7'h1e == r_count_17_io_out ? io_r_30_b : _GEN_1879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1881 = 7'h1f == r_count_17_io_out ? io_r_31_b : _GEN_1880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1882 = 7'h20 == r_count_17_io_out ? io_r_32_b : _GEN_1881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1883 = 7'h21 == r_count_17_io_out ? io_r_33_b : _GEN_1882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1884 = 7'h22 == r_count_17_io_out ? io_r_34_b : _GEN_1883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1885 = 7'h23 == r_count_17_io_out ? io_r_35_b : _GEN_1884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1886 = 7'h24 == r_count_17_io_out ? io_r_36_b : _GEN_1885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1887 = 7'h25 == r_count_17_io_out ? io_r_37_b : _GEN_1886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1888 = 7'h26 == r_count_17_io_out ? io_r_38_b : _GEN_1887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1889 = 7'h27 == r_count_17_io_out ? io_r_39_b : _GEN_1888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1890 = 7'h28 == r_count_17_io_out ? io_r_40_b : _GEN_1889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1891 = 7'h29 == r_count_17_io_out ? io_r_41_b : _GEN_1890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1892 = 7'h2a == r_count_17_io_out ? io_r_42_b : _GEN_1891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1893 = 7'h2b == r_count_17_io_out ? io_r_43_b : _GEN_1892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1894 = 7'h2c == r_count_17_io_out ? io_r_44_b : _GEN_1893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1895 = 7'h2d == r_count_17_io_out ? io_r_45_b : _GEN_1894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1896 = 7'h2e == r_count_17_io_out ? io_r_46_b : _GEN_1895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1897 = 7'h2f == r_count_17_io_out ? io_r_47_b : _GEN_1896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1898 = 7'h30 == r_count_17_io_out ? io_r_48_b : _GEN_1897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1899 = 7'h31 == r_count_17_io_out ? io_r_49_b : _GEN_1898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1900 = 7'h32 == r_count_17_io_out ? io_r_50_b : _GEN_1899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1901 = 7'h33 == r_count_17_io_out ? io_r_51_b : _GEN_1900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1902 = 7'h34 == r_count_17_io_out ? io_r_52_b : _GEN_1901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1903 = 7'h35 == r_count_17_io_out ? io_r_53_b : _GEN_1902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1904 = 7'h36 == r_count_17_io_out ? io_r_54_b : _GEN_1903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1905 = 7'h37 == r_count_17_io_out ? io_r_55_b : _GEN_1904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1906 = 7'h38 == r_count_17_io_out ? io_r_56_b : _GEN_1905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1907 = 7'h39 == r_count_17_io_out ? io_r_57_b : _GEN_1906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1908 = 7'h3a == r_count_17_io_out ? io_r_58_b : _GEN_1907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1909 = 7'h3b == r_count_17_io_out ? io_r_59_b : _GEN_1908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1910 = 7'h3c == r_count_17_io_out ? io_r_60_b : _GEN_1909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1911 = 7'h3d == r_count_17_io_out ? io_r_61_b : _GEN_1910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1912 = 7'h3e == r_count_17_io_out ? io_r_62_b : _GEN_1911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1913 = 7'h3f == r_count_17_io_out ? io_r_63_b : _GEN_1912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1914 = 7'h40 == r_count_17_io_out ? io_r_64_b : _GEN_1913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1915 = 7'h41 == r_count_17_io_out ? io_r_65_b : _GEN_1914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1916 = 7'h42 == r_count_17_io_out ? io_r_66_b : _GEN_1915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1917 = 7'h43 == r_count_17_io_out ? io_r_67_b : _GEN_1916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1918 = 7'h44 == r_count_17_io_out ? io_r_68_b : _GEN_1917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1919 = 7'h45 == r_count_17_io_out ? io_r_69_b : _GEN_1918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1920 = 7'h46 == r_count_17_io_out ? io_r_70_b : _GEN_1919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1921 = 7'h47 == r_count_17_io_out ? io_r_71_b : _GEN_1920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1922 = 7'h48 == r_count_17_io_out ? io_r_72_b : _GEN_1921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1923 = 7'h49 == r_count_17_io_out ? io_r_73_b : _GEN_1922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1924 = 7'h4a == r_count_17_io_out ? io_r_74_b : _GEN_1923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1925 = 7'h4b == r_count_17_io_out ? io_r_75_b : _GEN_1924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1926 = 7'h4c == r_count_17_io_out ? io_r_76_b : _GEN_1925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1927 = 7'h4d == r_count_17_io_out ? io_r_77_b : _GEN_1926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1928 = 7'h4e == r_count_17_io_out ? io_r_78_b : _GEN_1927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1929 = 7'h4f == r_count_17_io_out ? io_r_79_b : _GEN_1928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1930 = 7'h50 == r_count_17_io_out ? io_r_80_b : _GEN_1929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1931 = 7'h51 == r_count_17_io_out ? io_r_81_b : _GEN_1930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1932 = 7'h52 == r_count_17_io_out ? io_r_82_b : _GEN_1931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1933 = 7'h53 == r_count_17_io_out ? io_r_83_b : _GEN_1932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1934 = 7'h54 == r_count_17_io_out ? io_r_84_b : _GEN_1933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1935 = 7'h55 == r_count_17_io_out ? io_r_85_b : _GEN_1934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1936 = 7'h56 == r_count_17_io_out ? io_r_86_b : _GEN_1935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1937 = 7'h57 == r_count_17_io_out ? io_r_87_b : _GEN_1936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1938 = 7'h58 == r_count_17_io_out ? io_r_88_b : _GEN_1937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1939 = 7'h59 == r_count_17_io_out ? io_r_89_b : _GEN_1938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1940 = 7'h5a == r_count_17_io_out ? io_r_90_b : _GEN_1939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1941 = 7'h5b == r_count_17_io_out ? io_r_91_b : _GEN_1940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1942 = 7'h5c == r_count_17_io_out ? io_r_92_b : _GEN_1941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1943 = 7'h5d == r_count_17_io_out ? io_r_93_b : _GEN_1942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1944 = 7'h5e == r_count_17_io_out ? io_r_94_b : _GEN_1943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1945 = 7'h5f == r_count_17_io_out ? io_r_95_b : _GEN_1944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1946 = 7'h60 == r_count_17_io_out ? io_r_96_b : _GEN_1945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1947 = 7'h61 == r_count_17_io_out ? io_r_97_b : _GEN_1946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1948 = 7'h62 == r_count_17_io_out ? io_r_98_b : _GEN_1947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1951 = 7'h1 == r_count_18_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1952 = 7'h2 == r_count_18_io_out ? io_r_2_b : _GEN_1951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1953 = 7'h3 == r_count_18_io_out ? io_r_3_b : _GEN_1952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1954 = 7'h4 == r_count_18_io_out ? io_r_4_b : _GEN_1953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1955 = 7'h5 == r_count_18_io_out ? io_r_5_b : _GEN_1954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1956 = 7'h6 == r_count_18_io_out ? io_r_6_b : _GEN_1955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1957 = 7'h7 == r_count_18_io_out ? io_r_7_b : _GEN_1956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1958 = 7'h8 == r_count_18_io_out ? io_r_8_b : _GEN_1957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1959 = 7'h9 == r_count_18_io_out ? io_r_9_b : _GEN_1958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1960 = 7'ha == r_count_18_io_out ? io_r_10_b : _GEN_1959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1961 = 7'hb == r_count_18_io_out ? io_r_11_b : _GEN_1960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1962 = 7'hc == r_count_18_io_out ? io_r_12_b : _GEN_1961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1963 = 7'hd == r_count_18_io_out ? io_r_13_b : _GEN_1962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1964 = 7'he == r_count_18_io_out ? io_r_14_b : _GEN_1963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1965 = 7'hf == r_count_18_io_out ? io_r_15_b : _GEN_1964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1966 = 7'h10 == r_count_18_io_out ? io_r_16_b : _GEN_1965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1967 = 7'h11 == r_count_18_io_out ? io_r_17_b : _GEN_1966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1968 = 7'h12 == r_count_18_io_out ? io_r_18_b : _GEN_1967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1969 = 7'h13 == r_count_18_io_out ? io_r_19_b : _GEN_1968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1970 = 7'h14 == r_count_18_io_out ? io_r_20_b : _GEN_1969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1971 = 7'h15 == r_count_18_io_out ? io_r_21_b : _GEN_1970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1972 = 7'h16 == r_count_18_io_out ? io_r_22_b : _GEN_1971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1973 = 7'h17 == r_count_18_io_out ? io_r_23_b : _GEN_1972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1974 = 7'h18 == r_count_18_io_out ? io_r_24_b : _GEN_1973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1975 = 7'h19 == r_count_18_io_out ? io_r_25_b : _GEN_1974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1976 = 7'h1a == r_count_18_io_out ? io_r_26_b : _GEN_1975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1977 = 7'h1b == r_count_18_io_out ? io_r_27_b : _GEN_1976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1978 = 7'h1c == r_count_18_io_out ? io_r_28_b : _GEN_1977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1979 = 7'h1d == r_count_18_io_out ? io_r_29_b : _GEN_1978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1980 = 7'h1e == r_count_18_io_out ? io_r_30_b : _GEN_1979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1981 = 7'h1f == r_count_18_io_out ? io_r_31_b : _GEN_1980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1982 = 7'h20 == r_count_18_io_out ? io_r_32_b : _GEN_1981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1983 = 7'h21 == r_count_18_io_out ? io_r_33_b : _GEN_1982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1984 = 7'h22 == r_count_18_io_out ? io_r_34_b : _GEN_1983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1985 = 7'h23 == r_count_18_io_out ? io_r_35_b : _GEN_1984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1986 = 7'h24 == r_count_18_io_out ? io_r_36_b : _GEN_1985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1987 = 7'h25 == r_count_18_io_out ? io_r_37_b : _GEN_1986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1988 = 7'h26 == r_count_18_io_out ? io_r_38_b : _GEN_1987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1989 = 7'h27 == r_count_18_io_out ? io_r_39_b : _GEN_1988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1990 = 7'h28 == r_count_18_io_out ? io_r_40_b : _GEN_1989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1991 = 7'h29 == r_count_18_io_out ? io_r_41_b : _GEN_1990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1992 = 7'h2a == r_count_18_io_out ? io_r_42_b : _GEN_1991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1993 = 7'h2b == r_count_18_io_out ? io_r_43_b : _GEN_1992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1994 = 7'h2c == r_count_18_io_out ? io_r_44_b : _GEN_1993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1995 = 7'h2d == r_count_18_io_out ? io_r_45_b : _GEN_1994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1996 = 7'h2e == r_count_18_io_out ? io_r_46_b : _GEN_1995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1997 = 7'h2f == r_count_18_io_out ? io_r_47_b : _GEN_1996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1998 = 7'h30 == r_count_18_io_out ? io_r_48_b : _GEN_1997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_1999 = 7'h31 == r_count_18_io_out ? io_r_49_b : _GEN_1998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2000 = 7'h32 == r_count_18_io_out ? io_r_50_b : _GEN_1999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2001 = 7'h33 == r_count_18_io_out ? io_r_51_b : _GEN_2000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2002 = 7'h34 == r_count_18_io_out ? io_r_52_b : _GEN_2001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2003 = 7'h35 == r_count_18_io_out ? io_r_53_b : _GEN_2002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2004 = 7'h36 == r_count_18_io_out ? io_r_54_b : _GEN_2003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2005 = 7'h37 == r_count_18_io_out ? io_r_55_b : _GEN_2004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2006 = 7'h38 == r_count_18_io_out ? io_r_56_b : _GEN_2005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2007 = 7'h39 == r_count_18_io_out ? io_r_57_b : _GEN_2006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2008 = 7'h3a == r_count_18_io_out ? io_r_58_b : _GEN_2007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2009 = 7'h3b == r_count_18_io_out ? io_r_59_b : _GEN_2008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2010 = 7'h3c == r_count_18_io_out ? io_r_60_b : _GEN_2009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2011 = 7'h3d == r_count_18_io_out ? io_r_61_b : _GEN_2010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2012 = 7'h3e == r_count_18_io_out ? io_r_62_b : _GEN_2011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2013 = 7'h3f == r_count_18_io_out ? io_r_63_b : _GEN_2012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2014 = 7'h40 == r_count_18_io_out ? io_r_64_b : _GEN_2013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2015 = 7'h41 == r_count_18_io_out ? io_r_65_b : _GEN_2014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2016 = 7'h42 == r_count_18_io_out ? io_r_66_b : _GEN_2015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2017 = 7'h43 == r_count_18_io_out ? io_r_67_b : _GEN_2016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2018 = 7'h44 == r_count_18_io_out ? io_r_68_b : _GEN_2017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2019 = 7'h45 == r_count_18_io_out ? io_r_69_b : _GEN_2018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2020 = 7'h46 == r_count_18_io_out ? io_r_70_b : _GEN_2019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2021 = 7'h47 == r_count_18_io_out ? io_r_71_b : _GEN_2020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2022 = 7'h48 == r_count_18_io_out ? io_r_72_b : _GEN_2021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2023 = 7'h49 == r_count_18_io_out ? io_r_73_b : _GEN_2022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2024 = 7'h4a == r_count_18_io_out ? io_r_74_b : _GEN_2023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2025 = 7'h4b == r_count_18_io_out ? io_r_75_b : _GEN_2024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2026 = 7'h4c == r_count_18_io_out ? io_r_76_b : _GEN_2025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2027 = 7'h4d == r_count_18_io_out ? io_r_77_b : _GEN_2026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2028 = 7'h4e == r_count_18_io_out ? io_r_78_b : _GEN_2027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2029 = 7'h4f == r_count_18_io_out ? io_r_79_b : _GEN_2028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2030 = 7'h50 == r_count_18_io_out ? io_r_80_b : _GEN_2029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2031 = 7'h51 == r_count_18_io_out ? io_r_81_b : _GEN_2030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2032 = 7'h52 == r_count_18_io_out ? io_r_82_b : _GEN_2031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2033 = 7'h53 == r_count_18_io_out ? io_r_83_b : _GEN_2032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2034 = 7'h54 == r_count_18_io_out ? io_r_84_b : _GEN_2033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2035 = 7'h55 == r_count_18_io_out ? io_r_85_b : _GEN_2034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2036 = 7'h56 == r_count_18_io_out ? io_r_86_b : _GEN_2035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2037 = 7'h57 == r_count_18_io_out ? io_r_87_b : _GEN_2036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2038 = 7'h58 == r_count_18_io_out ? io_r_88_b : _GEN_2037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2039 = 7'h59 == r_count_18_io_out ? io_r_89_b : _GEN_2038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2040 = 7'h5a == r_count_18_io_out ? io_r_90_b : _GEN_2039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2041 = 7'h5b == r_count_18_io_out ? io_r_91_b : _GEN_2040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2042 = 7'h5c == r_count_18_io_out ? io_r_92_b : _GEN_2041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2043 = 7'h5d == r_count_18_io_out ? io_r_93_b : _GEN_2042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2044 = 7'h5e == r_count_18_io_out ? io_r_94_b : _GEN_2043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2045 = 7'h5f == r_count_18_io_out ? io_r_95_b : _GEN_2044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2046 = 7'h60 == r_count_18_io_out ? io_r_96_b : _GEN_2045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2047 = 7'h61 == r_count_18_io_out ? io_r_97_b : _GEN_2046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2048 = 7'h62 == r_count_18_io_out ? io_r_98_b : _GEN_2047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2051 = 7'h1 == r_count_19_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2052 = 7'h2 == r_count_19_io_out ? io_r_2_b : _GEN_2051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2053 = 7'h3 == r_count_19_io_out ? io_r_3_b : _GEN_2052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2054 = 7'h4 == r_count_19_io_out ? io_r_4_b : _GEN_2053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2055 = 7'h5 == r_count_19_io_out ? io_r_5_b : _GEN_2054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2056 = 7'h6 == r_count_19_io_out ? io_r_6_b : _GEN_2055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2057 = 7'h7 == r_count_19_io_out ? io_r_7_b : _GEN_2056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2058 = 7'h8 == r_count_19_io_out ? io_r_8_b : _GEN_2057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2059 = 7'h9 == r_count_19_io_out ? io_r_9_b : _GEN_2058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2060 = 7'ha == r_count_19_io_out ? io_r_10_b : _GEN_2059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2061 = 7'hb == r_count_19_io_out ? io_r_11_b : _GEN_2060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2062 = 7'hc == r_count_19_io_out ? io_r_12_b : _GEN_2061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2063 = 7'hd == r_count_19_io_out ? io_r_13_b : _GEN_2062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2064 = 7'he == r_count_19_io_out ? io_r_14_b : _GEN_2063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2065 = 7'hf == r_count_19_io_out ? io_r_15_b : _GEN_2064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2066 = 7'h10 == r_count_19_io_out ? io_r_16_b : _GEN_2065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2067 = 7'h11 == r_count_19_io_out ? io_r_17_b : _GEN_2066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2068 = 7'h12 == r_count_19_io_out ? io_r_18_b : _GEN_2067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2069 = 7'h13 == r_count_19_io_out ? io_r_19_b : _GEN_2068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2070 = 7'h14 == r_count_19_io_out ? io_r_20_b : _GEN_2069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2071 = 7'h15 == r_count_19_io_out ? io_r_21_b : _GEN_2070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2072 = 7'h16 == r_count_19_io_out ? io_r_22_b : _GEN_2071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2073 = 7'h17 == r_count_19_io_out ? io_r_23_b : _GEN_2072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2074 = 7'h18 == r_count_19_io_out ? io_r_24_b : _GEN_2073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2075 = 7'h19 == r_count_19_io_out ? io_r_25_b : _GEN_2074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2076 = 7'h1a == r_count_19_io_out ? io_r_26_b : _GEN_2075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2077 = 7'h1b == r_count_19_io_out ? io_r_27_b : _GEN_2076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2078 = 7'h1c == r_count_19_io_out ? io_r_28_b : _GEN_2077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2079 = 7'h1d == r_count_19_io_out ? io_r_29_b : _GEN_2078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2080 = 7'h1e == r_count_19_io_out ? io_r_30_b : _GEN_2079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2081 = 7'h1f == r_count_19_io_out ? io_r_31_b : _GEN_2080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2082 = 7'h20 == r_count_19_io_out ? io_r_32_b : _GEN_2081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2083 = 7'h21 == r_count_19_io_out ? io_r_33_b : _GEN_2082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2084 = 7'h22 == r_count_19_io_out ? io_r_34_b : _GEN_2083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2085 = 7'h23 == r_count_19_io_out ? io_r_35_b : _GEN_2084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2086 = 7'h24 == r_count_19_io_out ? io_r_36_b : _GEN_2085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2087 = 7'h25 == r_count_19_io_out ? io_r_37_b : _GEN_2086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2088 = 7'h26 == r_count_19_io_out ? io_r_38_b : _GEN_2087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2089 = 7'h27 == r_count_19_io_out ? io_r_39_b : _GEN_2088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2090 = 7'h28 == r_count_19_io_out ? io_r_40_b : _GEN_2089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2091 = 7'h29 == r_count_19_io_out ? io_r_41_b : _GEN_2090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2092 = 7'h2a == r_count_19_io_out ? io_r_42_b : _GEN_2091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2093 = 7'h2b == r_count_19_io_out ? io_r_43_b : _GEN_2092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2094 = 7'h2c == r_count_19_io_out ? io_r_44_b : _GEN_2093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2095 = 7'h2d == r_count_19_io_out ? io_r_45_b : _GEN_2094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2096 = 7'h2e == r_count_19_io_out ? io_r_46_b : _GEN_2095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2097 = 7'h2f == r_count_19_io_out ? io_r_47_b : _GEN_2096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2098 = 7'h30 == r_count_19_io_out ? io_r_48_b : _GEN_2097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2099 = 7'h31 == r_count_19_io_out ? io_r_49_b : _GEN_2098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2100 = 7'h32 == r_count_19_io_out ? io_r_50_b : _GEN_2099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2101 = 7'h33 == r_count_19_io_out ? io_r_51_b : _GEN_2100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2102 = 7'h34 == r_count_19_io_out ? io_r_52_b : _GEN_2101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2103 = 7'h35 == r_count_19_io_out ? io_r_53_b : _GEN_2102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2104 = 7'h36 == r_count_19_io_out ? io_r_54_b : _GEN_2103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2105 = 7'h37 == r_count_19_io_out ? io_r_55_b : _GEN_2104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2106 = 7'h38 == r_count_19_io_out ? io_r_56_b : _GEN_2105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2107 = 7'h39 == r_count_19_io_out ? io_r_57_b : _GEN_2106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2108 = 7'h3a == r_count_19_io_out ? io_r_58_b : _GEN_2107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2109 = 7'h3b == r_count_19_io_out ? io_r_59_b : _GEN_2108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2110 = 7'h3c == r_count_19_io_out ? io_r_60_b : _GEN_2109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2111 = 7'h3d == r_count_19_io_out ? io_r_61_b : _GEN_2110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2112 = 7'h3e == r_count_19_io_out ? io_r_62_b : _GEN_2111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2113 = 7'h3f == r_count_19_io_out ? io_r_63_b : _GEN_2112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2114 = 7'h40 == r_count_19_io_out ? io_r_64_b : _GEN_2113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2115 = 7'h41 == r_count_19_io_out ? io_r_65_b : _GEN_2114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2116 = 7'h42 == r_count_19_io_out ? io_r_66_b : _GEN_2115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2117 = 7'h43 == r_count_19_io_out ? io_r_67_b : _GEN_2116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2118 = 7'h44 == r_count_19_io_out ? io_r_68_b : _GEN_2117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2119 = 7'h45 == r_count_19_io_out ? io_r_69_b : _GEN_2118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2120 = 7'h46 == r_count_19_io_out ? io_r_70_b : _GEN_2119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2121 = 7'h47 == r_count_19_io_out ? io_r_71_b : _GEN_2120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2122 = 7'h48 == r_count_19_io_out ? io_r_72_b : _GEN_2121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2123 = 7'h49 == r_count_19_io_out ? io_r_73_b : _GEN_2122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2124 = 7'h4a == r_count_19_io_out ? io_r_74_b : _GEN_2123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2125 = 7'h4b == r_count_19_io_out ? io_r_75_b : _GEN_2124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2126 = 7'h4c == r_count_19_io_out ? io_r_76_b : _GEN_2125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2127 = 7'h4d == r_count_19_io_out ? io_r_77_b : _GEN_2126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2128 = 7'h4e == r_count_19_io_out ? io_r_78_b : _GEN_2127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2129 = 7'h4f == r_count_19_io_out ? io_r_79_b : _GEN_2128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2130 = 7'h50 == r_count_19_io_out ? io_r_80_b : _GEN_2129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2131 = 7'h51 == r_count_19_io_out ? io_r_81_b : _GEN_2130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2132 = 7'h52 == r_count_19_io_out ? io_r_82_b : _GEN_2131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2133 = 7'h53 == r_count_19_io_out ? io_r_83_b : _GEN_2132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2134 = 7'h54 == r_count_19_io_out ? io_r_84_b : _GEN_2133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2135 = 7'h55 == r_count_19_io_out ? io_r_85_b : _GEN_2134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2136 = 7'h56 == r_count_19_io_out ? io_r_86_b : _GEN_2135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2137 = 7'h57 == r_count_19_io_out ? io_r_87_b : _GEN_2136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2138 = 7'h58 == r_count_19_io_out ? io_r_88_b : _GEN_2137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2139 = 7'h59 == r_count_19_io_out ? io_r_89_b : _GEN_2138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2140 = 7'h5a == r_count_19_io_out ? io_r_90_b : _GEN_2139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2141 = 7'h5b == r_count_19_io_out ? io_r_91_b : _GEN_2140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2142 = 7'h5c == r_count_19_io_out ? io_r_92_b : _GEN_2141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2143 = 7'h5d == r_count_19_io_out ? io_r_93_b : _GEN_2142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2144 = 7'h5e == r_count_19_io_out ? io_r_94_b : _GEN_2143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2145 = 7'h5f == r_count_19_io_out ? io_r_95_b : _GEN_2144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2146 = 7'h60 == r_count_19_io_out ? io_r_96_b : _GEN_2145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2147 = 7'h61 == r_count_19_io_out ? io_r_97_b : _GEN_2146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2148 = 7'h62 == r_count_19_io_out ? io_r_98_b : _GEN_2147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2151 = 7'h1 == r_count_20_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2152 = 7'h2 == r_count_20_io_out ? io_r_2_b : _GEN_2151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2153 = 7'h3 == r_count_20_io_out ? io_r_3_b : _GEN_2152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2154 = 7'h4 == r_count_20_io_out ? io_r_4_b : _GEN_2153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2155 = 7'h5 == r_count_20_io_out ? io_r_5_b : _GEN_2154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2156 = 7'h6 == r_count_20_io_out ? io_r_6_b : _GEN_2155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2157 = 7'h7 == r_count_20_io_out ? io_r_7_b : _GEN_2156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2158 = 7'h8 == r_count_20_io_out ? io_r_8_b : _GEN_2157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2159 = 7'h9 == r_count_20_io_out ? io_r_9_b : _GEN_2158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2160 = 7'ha == r_count_20_io_out ? io_r_10_b : _GEN_2159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2161 = 7'hb == r_count_20_io_out ? io_r_11_b : _GEN_2160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2162 = 7'hc == r_count_20_io_out ? io_r_12_b : _GEN_2161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2163 = 7'hd == r_count_20_io_out ? io_r_13_b : _GEN_2162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2164 = 7'he == r_count_20_io_out ? io_r_14_b : _GEN_2163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2165 = 7'hf == r_count_20_io_out ? io_r_15_b : _GEN_2164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2166 = 7'h10 == r_count_20_io_out ? io_r_16_b : _GEN_2165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2167 = 7'h11 == r_count_20_io_out ? io_r_17_b : _GEN_2166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2168 = 7'h12 == r_count_20_io_out ? io_r_18_b : _GEN_2167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2169 = 7'h13 == r_count_20_io_out ? io_r_19_b : _GEN_2168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2170 = 7'h14 == r_count_20_io_out ? io_r_20_b : _GEN_2169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2171 = 7'h15 == r_count_20_io_out ? io_r_21_b : _GEN_2170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2172 = 7'h16 == r_count_20_io_out ? io_r_22_b : _GEN_2171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2173 = 7'h17 == r_count_20_io_out ? io_r_23_b : _GEN_2172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2174 = 7'h18 == r_count_20_io_out ? io_r_24_b : _GEN_2173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2175 = 7'h19 == r_count_20_io_out ? io_r_25_b : _GEN_2174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2176 = 7'h1a == r_count_20_io_out ? io_r_26_b : _GEN_2175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2177 = 7'h1b == r_count_20_io_out ? io_r_27_b : _GEN_2176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2178 = 7'h1c == r_count_20_io_out ? io_r_28_b : _GEN_2177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2179 = 7'h1d == r_count_20_io_out ? io_r_29_b : _GEN_2178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2180 = 7'h1e == r_count_20_io_out ? io_r_30_b : _GEN_2179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2181 = 7'h1f == r_count_20_io_out ? io_r_31_b : _GEN_2180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2182 = 7'h20 == r_count_20_io_out ? io_r_32_b : _GEN_2181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2183 = 7'h21 == r_count_20_io_out ? io_r_33_b : _GEN_2182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2184 = 7'h22 == r_count_20_io_out ? io_r_34_b : _GEN_2183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2185 = 7'h23 == r_count_20_io_out ? io_r_35_b : _GEN_2184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2186 = 7'h24 == r_count_20_io_out ? io_r_36_b : _GEN_2185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2187 = 7'h25 == r_count_20_io_out ? io_r_37_b : _GEN_2186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2188 = 7'h26 == r_count_20_io_out ? io_r_38_b : _GEN_2187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2189 = 7'h27 == r_count_20_io_out ? io_r_39_b : _GEN_2188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2190 = 7'h28 == r_count_20_io_out ? io_r_40_b : _GEN_2189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2191 = 7'h29 == r_count_20_io_out ? io_r_41_b : _GEN_2190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2192 = 7'h2a == r_count_20_io_out ? io_r_42_b : _GEN_2191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2193 = 7'h2b == r_count_20_io_out ? io_r_43_b : _GEN_2192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2194 = 7'h2c == r_count_20_io_out ? io_r_44_b : _GEN_2193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2195 = 7'h2d == r_count_20_io_out ? io_r_45_b : _GEN_2194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2196 = 7'h2e == r_count_20_io_out ? io_r_46_b : _GEN_2195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2197 = 7'h2f == r_count_20_io_out ? io_r_47_b : _GEN_2196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2198 = 7'h30 == r_count_20_io_out ? io_r_48_b : _GEN_2197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2199 = 7'h31 == r_count_20_io_out ? io_r_49_b : _GEN_2198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2200 = 7'h32 == r_count_20_io_out ? io_r_50_b : _GEN_2199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2201 = 7'h33 == r_count_20_io_out ? io_r_51_b : _GEN_2200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2202 = 7'h34 == r_count_20_io_out ? io_r_52_b : _GEN_2201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2203 = 7'h35 == r_count_20_io_out ? io_r_53_b : _GEN_2202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2204 = 7'h36 == r_count_20_io_out ? io_r_54_b : _GEN_2203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2205 = 7'h37 == r_count_20_io_out ? io_r_55_b : _GEN_2204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2206 = 7'h38 == r_count_20_io_out ? io_r_56_b : _GEN_2205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2207 = 7'h39 == r_count_20_io_out ? io_r_57_b : _GEN_2206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2208 = 7'h3a == r_count_20_io_out ? io_r_58_b : _GEN_2207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2209 = 7'h3b == r_count_20_io_out ? io_r_59_b : _GEN_2208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2210 = 7'h3c == r_count_20_io_out ? io_r_60_b : _GEN_2209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2211 = 7'h3d == r_count_20_io_out ? io_r_61_b : _GEN_2210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2212 = 7'h3e == r_count_20_io_out ? io_r_62_b : _GEN_2211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2213 = 7'h3f == r_count_20_io_out ? io_r_63_b : _GEN_2212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2214 = 7'h40 == r_count_20_io_out ? io_r_64_b : _GEN_2213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2215 = 7'h41 == r_count_20_io_out ? io_r_65_b : _GEN_2214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2216 = 7'h42 == r_count_20_io_out ? io_r_66_b : _GEN_2215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2217 = 7'h43 == r_count_20_io_out ? io_r_67_b : _GEN_2216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2218 = 7'h44 == r_count_20_io_out ? io_r_68_b : _GEN_2217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2219 = 7'h45 == r_count_20_io_out ? io_r_69_b : _GEN_2218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2220 = 7'h46 == r_count_20_io_out ? io_r_70_b : _GEN_2219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2221 = 7'h47 == r_count_20_io_out ? io_r_71_b : _GEN_2220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2222 = 7'h48 == r_count_20_io_out ? io_r_72_b : _GEN_2221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2223 = 7'h49 == r_count_20_io_out ? io_r_73_b : _GEN_2222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2224 = 7'h4a == r_count_20_io_out ? io_r_74_b : _GEN_2223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2225 = 7'h4b == r_count_20_io_out ? io_r_75_b : _GEN_2224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2226 = 7'h4c == r_count_20_io_out ? io_r_76_b : _GEN_2225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2227 = 7'h4d == r_count_20_io_out ? io_r_77_b : _GEN_2226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2228 = 7'h4e == r_count_20_io_out ? io_r_78_b : _GEN_2227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2229 = 7'h4f == r_count_20_io_out ? io_r_79_b : _GEN_2228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2230 = 7'h50 == r_count_20_io_out ? io_r_80_b : _GEN_2229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2231 = 7'h51 == r_count_20_io_out ? io_r_81_b : _GEN_2230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2232 = 7'h52 == r_count_20_io_out ? io_r_82_b : _GEN_2231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2233 = 7'h53 == r_count_20_io_out ? io_r_83_b : _GEN_2232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2234 = 7'h54 == r_count_20_io_out ? io_r_84_b : _GEN_2233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2235 = 7'h55 == r_count_20_io_out ? io_r_85_b : _GEN_2234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2236 = 7'h56 == r_count_20_io_out ? io_r_86_b : _GEN_2235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2237 = 7'h57 == r_count_20_io_out ? io_r_87_b : _GEN_2236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2238 = 7'h58 == r_count_20_io_out ? io_r_88_b : _GEN_2237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2239 = 7'h59 == r_count_20_io_out ? io_r_89_b : _GEN_2238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2240 = 7'h5a == r_count_20_io_out ? io_r_90_b : _GEN_2239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2241 = 7'h5b == r_count_20_io_out ? io_r_91_b : _GEN_2240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2242 = 7'h5c == r_count_20_io_out ? io_r_92_b : _GEN_2241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2243 = 7'h5d == r_count_20_io_out ? io_r_93_b : _GEN_2242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2244 = 7'h5e == r_count_20_io_out ? io_r_94_b : _GEN_2243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2245 = 7'h5f == r_count_20_io_out ? io_r_95_b : _GEN_2244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2246 = 7'h60 == r_count_20_io_out ? io_r_96_b : _GEN_2245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2247 = 7'h61 == r_count_20_io_out ? io_r_97_b : _GEN_2246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2248 = 7'h62 == r_count_20_io_out ? io_r_98_b : _GEN_2247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2251 = 7'h1 == r_count_21_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2252 = 7'h2 == r_count_21_io_out ? io_r_2_b : _GEN_2251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2253 = 7'h3 == r_count_21_io_out ? io_r_3_b : _GEN_2252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2254 = 7'h4 == r_count_21_io_out ? io_r_4_b : _GEN_2253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2255 = 7'h5 == r_count_21_io_out ? io_r_5_b : _GEN_2254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2256 = 7'h6 == r_count_21_io_out ? io_r_6_b : _GEN_2255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2257 = 7'h7 == r_count_21_io_out ? io_r_7_b : _GEN_2256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2258 = 7'h8 == r_count_21_io_out ? io_r_8_b : _GEN_2257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2259 = 7'h9 == r_count_21_io_out ? io_r_9_b : _GEN_2258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2260 = 7'ha == r_count_21_io_out ? io_r_10_b : _GEN_2259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2261 = 7'hb == r_count_21_io_out ? io_r_11_b : _GEN_2260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2262 = 7'hc == r_count_21_io_out ? io_r_12_b : _GEN_2261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2263 = 7'hd == r_count_21_io_out ? io_r_13_b : _GEN_2262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2264 = 7'he == r_count_21_io_out ? io_r_14_b : _GEN_2263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2265 = 7'hf == r_count_21_io_out ? io_r_15_b : _GEN_2264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2266 = 7'h10 == r_count_21_io_out ? io_r_16_b : _GEN_2265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2267 = 7'h11 == r_count_21_io_out ? io_r_17_b : _GEN_2266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2268 = 7'h12 == r_count_21_io_out ? io_r_18_b : _GEN_2267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2269 = 7'h13 == r_count_21_io_out ? io_r_19_b : _GEN_2268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2270 = 7'h14 == r_count_21_io_out ? io_r_20_b : _GEN_2269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2271 = 7'h15 == r_count_21_io_out ? io_r_21_b : _GEN_2270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2272 = 7'h16 == r_count_21_io_out ? io_r_22_b : _GEN_2271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2273 = 7'h17 == r_count_21_io_out ? io_r_23_b : _GEN_2272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2274 = 7'h18 == r_count_21_io_out ? io_r_24_b : _GEN_2273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2275 = 7'h19 == r_count_21_io_out ? io_r_25_b : _GEN_2274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2276 = 7'h1a == r_count_21_io_out ? io_r_26_b : _GEN_2275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2277 = 7'h1b == r_count_21_io_out ? io_r_27_b : _GEN_2276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2278 = 7'h1c == r_count_21_io_out ? io_r_28_b : _GEN_2277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2279 = 7'h1d == r_count_21_io_out ? io_r_29_b : _GEN_2278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2280 = 7'h1e == r_count_21_io_out ? io_r_30_b : _GEN_2279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2281 = 7'h1f == r_count_21_io_out ? io_r_31_b : _GEN_2280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2282 = 7'h20 == r_count_21_io_out ? io_r_32_b : _GEN_2281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2283 = 7'h21 == r_count_21_io_out ? io_r_33_b : _GEN_2282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2284 = 7'h22 == r_count_21_io_out ? io_r_34_b : _GEN_2283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2285 = 7'h23 == r_count_21_io_out ? io_r_35_b : _GEN_2284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2286 = 7'h24 == r_count_21_io_out ? io_r_36_b : _GEN_2285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2287 = 7'h25 == r_count_21_io_out ? io_r_37_b : _GEN_2286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2288 = 7'h26 == r_count_21_io_out ? io_r_38_b : _GEN_2287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2289 = 7'h27 == r_count_21_io_out ? io_r_39_b : _GEN_2288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2290 = 7'h28 == r_count_21_io_out ? io_r_40_b : _GEN_2289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2291 = 7'h29 == r_count_21_io_out ? io_r_41_b : _GEN_2290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2292 = 7'h2a == r_count_21_io_out ? io_r_42_b : _GEN_2291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2293 = 7'h2b == r_count_21_io_out ? io_r_43_b : _GEN_2292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2294 = 7'h2c == r_count_21_io_out ? io_r_44_b : _GEN_2293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2295 = 7'h2d == r_count_21_io_out ? io_r_45_b : _GEN_2294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2296 = 7'h2e == r_count_21_io_out ? io_r_46_b : _GEN_2295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2297 = 7'h2f == r_count_21_io_out ? io_r_47_b : _GEN_2296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2298 = 7'h30 == r_count_21_io_out ? io_r_48_b : _GEN_2297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2299 = 7'h31 == r_count_21_io_out ? io_r_49_b : _GEN_2298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2300 = 7'h32 == r_count_21_io_out ? io_r_50_b : _GEN_2299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2301 = 7'h33 == r_count_21_io_out ? io_r_51_b : _GEN_2300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2302 = 7'h34 == r_count_21_io_out ? io_r_52_b : _GEN_2301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2303 = 7'h35 == r_count_21_io_out ? io_r_53_b : _GEN_2302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2304 = 7'h36 == r_count_21_io_out ? io_r_54_b : _GEN_2303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2305 = 7'h37 == r_count_21_io_out ? io_r_55_b : _GEN_2304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2306 = 7'h38 == r_count_21_io_out ? io_r_56_b : _GEN_2305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2307 = 7'h39 == r_count_21_io_out ? io_r_57_b : _GEN_2306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2308 = 7'h3a == r_count_21_io_out ? io_r_58_b : _GEN_2307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2309 = 7'h3b == r_count_21_io_out ? io_r_59_b : _GEN_2308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2310 = 7'h3c == r_count_21_io_out ? io_r_60_b : _GEN_2309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2311 = 7'h3d == r_count_21_io_out ? io_r_61_b : _GEN_2310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2312 = 7'h3e == r_count_21_io_out ? io_r_62_b : _GEN_2311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2313 = 7'h3f == r_count_21_io_out ? io_r_63_b : _GEN_2312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2314 = 7'h40 == r_count_21_io_out ? io_r_64_b : _GEN_2313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2315 = 7'h41 == r_count_21_io_out ? io_r_65_b : _GEN_2314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2316 = 7'h42 == r_count_21_io_out ? io_r_66_b : _GEN_2315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2317 = 7'h43 == r_count_21_io_out ? io_r_67_b : _GEN_2316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2318 = 7'h44 == r_count_21_io_out ? io_r_68_b : _GEN_2317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2319 = 7'h45 == r_count_21_io_out ? io_r_69_b : _GEN_2318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2320 = 7'h46 == r_count_21_io_out ? io_r_70_b : _GEN_2319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2321 = 7'h47 == r_count_21_io_out ? io_r_71_b : _GEN_2320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2322 = 7'h48 == r_count_21_io_out ? io_r_72_b : _GEN_2321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2323 = 7'h49 == r_count_21_io_out ? io_r_73_b : _GEN_2322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2324 = 7'h4a == r_count_21_io_out ? io_r_74_b : _GEN_2323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2325 = 7'h4b == r_count_21_io_out ? io_r_75_b : _GEN_2324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2326 = 7'h4c == r_count_21_io_out ? io_r_76_b : _GEN_2325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2327 = 7'h4d == r_count_21_io_out ? io_r_77_b : _GEN_2326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2328 = 7'h4e == r_count_21_io_out ? io_r_78_b : _GEN_2327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2329 = 7'h4f == r_count_21_io_out ? io_r_79_b : _GEN_2328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2330 = 7'h50 == r_count_21_io_out ? io_r_80_b : _GEN_2329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2331 = 7'h51 == r_count_21_io_out ? io_r_81_b : _GEN_2330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2332 = 7'h52 == r_count_21_io_out ? io_r_82_b : _GEN_2331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2333 = 7'h53 == r_count_21_io_out ? io_r_83_b : _GEN_2332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2334 = 7'h54 == r_count_21_io_out ? io_r_84_b : _GEN_2333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2335 = 7'h55 == r_count_21_io_out ? io_r_85_b : _GEN_2334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2336 = 7'h56 == r_count_21_io_out ? io_r_86_b : _GEN_2335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2337 = 7'h57 == r_count_21_io_out ? io_r_87_b : _GEN_2336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2338 = 7'h58 == r_count_21_io_out ? io_r_88_b : _GEN_2337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2339 = 7'h59 == r_count_21_io_out ? io_r_89_b : _GEN_2338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2340 = 7'h5a == r_count_21_io_out ? io_r_90_b : _GEN_2339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2341 = 7'h5b == r_count_21_io_out ? io_r_91_b : _GEN_2340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2342 = 7'h5c == r_count_21_io_out ? io_r_92_b : _GEN_2341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2343 = 7'h5d == r_count_21_io_out ? io_r_93_b : _GEN_2342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2344 = 7'h5e == r_count_21_io_out ? io_r_94_b : _GEN_2343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2345 = 7'h5f == r_count_21_io_out ? io_r_95_b : _GEN_2344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2346 = 7'h60 == r_count_21_io_out ? io_r_96_b : _GEN_2345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2347 = 7'h61 == r_count_21_io_out ? io_r_97_b : _GEN_2346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2348 = 7'h62 == r_count_21_io_out ? io_r_98_b : _GEN_2347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2351 = 7'h1 == r_count_22_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2352 = 7'h2 == r_count_22_io_out ? io_r_2_b : _GEN_2351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2353 = 7'h3 == r_count_22_io_out ? io_r_3_b : _GEN_2352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2354 = 7'h4 == r_count_22_io_out ? io_r_4_b : _GEN_2353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2355 = 7'h5 == r_count_22_io_out ? io_r_5_b : _GEN_2354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2356 = 7'h6 == r_count_22_io_out ? io_r_6_b : _GEN_2355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2357 = 7'h7 == r_count_22_io_out ? io_r_7_b : _GEN_2356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2358 = 7'h8 == r_count_22_io_out ? io_r_8_b : _GEN_2357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2359 = 7'h9 == r_count_22_io_out ? io_r_9_b : _GEN_2358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2360 = 7'ha == r_count_22_io_out ? io_r_10_b : _GEN_2359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2361 = 7'hb == r_count_22_io_out ? io_r_11_b : _GEN_2360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2362 = 7'hc == r_count_22_io_out ? io_r_12_b : _GEN_2361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2363 = 7'hd == r_count_22_io_out ? io_r_13_b : _GEN_2362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2364 = 7'he == r_count_22_io_out ? io_r_14_b : _GEN_2363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2365 = 7'hf == r_count_22_io_out ? io_r_15_b : _GEN_2364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2366 = 7'h10 == r_count_22_io_out ? io_r_16_b : _GEN_2365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2367 = 7'h11 == r_count_22_io_out ? io_r_17_b : _GEN_2366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2368 = 7'h12 == r_count_22_io_out ? io_r_18_b : _GEN_2367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2369 = 7'h13 == r_count_22_io_out ? io_r_19_b : _GEN_2368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2370 = 7'h14 == r_count_22_io_out ? io_r_20_b : _GEN_2369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2371 = 7'h15 == r_count_22_io_out ? io_r_21_b : _GEN_2370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2372 = 7'h16 == r_count_22_io_out ? io_r_22_b : _GEN_2371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2373 = 7'h17 == r_count_22_io_out ? io_r_23_b : _GEN_2372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2374 = 7'h18 == r_count_22_io_out ? io_r_24_b : _GEN_2373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2375 = 7'h19 == r_count_22_io_out ? io_r_25_b : _GEN_2374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2376 = 7'h1a == r_count_22_io_out ? io_r_26_b : _GEN_2375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2377 = 7'h1b == r_count_22_io_out ? io_r_27_b : _GEN_2376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2378 = 7'h1c == r_count_22_io_out ? io_r_28_b : _GEN_2377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2379 = 7'h1d == r_count_22_io_out ? io_r_29_b : _GEN_2378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2380 = 7'h1e == r_count_22_io_out ? io_r_30_b : _GEN_2379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2381 = 7'h1f == r_count_22_io_out ? io_r_31_b : _GEN_2380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2382 = 7'h20 == r_count_22_io_out ? io_r_32_b : _GEN_2381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2383 = 7'h21 == r_count_22_io_out ? io_r_33_b : _GEN_2382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2384 = 7'h22 == r_count_22_io_out ? io_r_34_b : _GEN_2383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2385 = 7'h23 == r_count_22_io_out ? io_r_35_b : _GEN_2384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2386 = 7'h24 == r_count_22_io_out ? io_r_36_b : _GEN_2385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2387 = 7'h25 == r_count_22_io_out ? io_r_37_b : _GEN_2386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2388 = 7'h26 == r_count_22_io_out ? io_r_38_b : _GEN_2387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2389 = 7'h27 == r_count_22_io_out ? io_r_39_b : _GEN_2388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2390 = 7'h28 == r_count_22_io_out ? io_r_40_b : _GEN_2389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2391 = 7'h29 == r_count_22_io_out ? io_r_41_b : _GEN_2390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2392 = 7'h2a == r_count_22_io_out ? io_r_42_b : _GEN_2391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2393 = 7'h2b == r_count_22_io_out ? io_r_43_b : _GEN_2392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2394 = 7'h2c == r_count_22_io_out ? io_r_44_b : _GEN_2393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2395 = 7'h2d == r_count_22_io_out ? io_r_45_b : _GEN_2394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2396 = 7'h2e == r_count_22_io_out ? io_r_46_b : _GEN_2395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2397 = 7'h2f == r_count_22_io_out ? io_r_47_b : _GEN_2396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2398 = 7'h30 == r_count_22_io_out ? io_r_48_b : _GEN_2397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2399 = 7'h31 == r_count_22_io_out ? io_r_49_b : _GEN_2398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2400 = 7'h32 == r_count_22_io_out ? io_r_50_b : _GEN_2399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2401 = 7'h33 == r_count_22_io_out ? io_r_51_b : _GEN_2400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2402 = 7'h34 == r_count_22_io_out ? io_r_52_b : _GEN_2401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2403 = 7'h35 == r_count_22_io_out ? io_r_53_b : _GEN_2402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2404 = 7'h36 == r_count_22_io_out ? io_r_54_b : _GEN_2403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2405 = 7'h37 == r_count_22_io_out ? io_r_55_b : _GEN_2404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2406 = 7'h38 == r_count_22_io_out ? io_r_56_b : _GEN_2405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2407 = 7'h39 == r_count_22_io_out ? io_r_57_b : _GEN_2406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2408 = 7'h3a == r_count_22_io_out ? io_r_58_b : _GEN_2407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2409 = 7'h3b == r_count_22_io_out ? io_r_59_b : _GEN_2408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2410 = 7'h3c == r_count_22_io_out ? io_r_60_b : _GEN_2409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2411 = 7'h3d == r_count_22_io_out ? io_r_61_b : _GEN_2410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2412 = 7'h3e == r_count_22_io_out ? io_r_62_b : _GEN_2411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2413 = 7'h3f == r_count_22_io_out ? io_r_63_b : _GEN_2412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2414 = 7'h40 == r_count_22_io_out ? io_r_64_b : _GEN_2413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2415 = 7'h41 == r_count_22_io_out ? io_r_65_b : _GEN_2414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2416 = 7'h42 == r_count_22_io_out ? io_r_66_b : _GEN_2415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2417 = 7'h43 == r_count_22_io_out ? io_r_67_b : _GEN_2416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2418 = 7'h44 == r_count_22_io_out ? io_r_68_b : _GEN_2417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2419 = 7'h45 == r_count_22_io_out ? io_r_69_b : _GEN_2418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2420 = 7'h46 == r_count_22_io_out ? io_r_70_b : _GEN_2419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2421 = 7'h47 == r_count_22_io_out ? io_r_71_b : _GEN_2420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2422 = 7'h48 == r_count_22_io_out ? io_r_72_b : _GEN_2421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2423 = 7'h49 == r_count_22_io_out ? io_r_73_b : _GEN_2422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2424 = 7'h4a == r_count_22_io_out ? io_r_74_b : _GEN_2423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2425 = 7'h4b == r_count_22_io_out ? io_r_75_b : _GEN_2424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2426 = 7'h4c == r_count_22_io_out ? io_r_76_b : _GEN_2425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2427 = 7'h4d == r_count_22_io_out ? io_r_77_b : _GEN_2426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2428 = 7'h4e == r_count_22_io_out ? io_r_78_b : _GEN_2427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2429 = 7'h4f == r_count_22_io_out ? io_r_79_b : _GEN_2428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2430 = 7'h50 == r_count_22_io_out ? io_r_80_b : _GEN_2429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2431 = 7'h51 == r_count_22_io_out ? io_r_81_b : _GEN_2430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2432 = 7'h52 == r_count_22_io_out ? io_r_82_b : _GEN_2431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2433 = 7'h53 == r_count_22_io_out ? io_r_83_b : _GEN_2432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2434 = 7'h54 == r_count_22_io_out ? io_r_84_b : _GEN_2433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2435 = 7'h55 == r_count_22_io_out ? io_r_85_b : _GEN_2434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2436 = 7'h56 == r_count_22_io_out ? io_r_86_b : _GEN_2435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2437 = 7'h57 == r_count_22_io_out ? io_r_87_b : _GEN_2436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2438 = 7'h58 == r_count_22_io_out ? io_r_88_b : _GEN_2437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2439 = 7'h59 == r_count_22_io_out ? io_r_89_b : _GEN_2438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2440 = 7'h5a == r_count_22_io_out ? io_r_90_b : _GEN_2439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2441 = 7'h5b == r_count_22_io_out ? io_r_91_b : _GEN_2440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2442 = 7'h5c == r_count_22_io_out ? io_r_92_b : _GEN_2441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2443 = 7'h5d == r_count_22_io_out ? io_r_93_b : _GEN_2442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2444 = 7'h5e == r_count_22_io_out ? io_r_94_b : _GEN_2443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2445 = 7'h5f == r_count_22_io_out ? io_r_95_b : _GEN_2444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2446 = 7'h60 == r_count_22_io_out ? io_r_96_b : _GEN_2445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2447 = 7'h61 == r_count_22_io_out ? io_r_97_b : _GEN_2446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2448 = 7'h62 == r_count_22_io_out ? io_r_98_b : _GEN_2447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2451 = 7'h1 == r_count_23_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2452 = 7'h2 == r_count_23_io_out ? io_r_2_b : _GEN_2451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2453 = 7'h3 == r_count_23_io_out ? io_r_3_b : _GEN_2452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2454 = 7'h4 == r_count_23_io_out ? io_r_4_b : _GEN_2453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2455 = 7'h5 == r_count_23_io_out ? io_r_5_b : _GEN_2454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2456 = 7'h6 == r_count_23_io_out ? io_r_6_b : _GEN_2455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2457 = 7'h7 == r_count_23_io_out ? io_r_7_b : _GEN_2456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2458 = 7'h8 == r_count_23_io_out ? io_r_8_b : _GEN_2457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2459 = 7'h9 == r_count_23_io_out ? io_r_9_b : _GEN_2458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2460 = 7'ha == r_count_23_io_out ? io_r_10_b : _GEN_2459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2461 = 7'hb == r_count_23_io_out ? io_r_11_b : _GEN_2460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2462 = 7'hc == r_count_23_io_out ? io_r_12_b : _GEN_2461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2463 = 7'hd == r_count_23_io_out ? io_r_13_b : _GEN_2462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2464 = 7'he == r_count_23_io_out ? io_r_14_b : _GEN_2463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2465 = 7'hf == r_count_23_io_out ? io_r_15_b : _GEN_2464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2466 = 7'h10 == r_count_23_io_out ? io_r_16_b : _GEN_2465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2467 = 7'h11 == r_count_23_io_out ? io_r_17_b : _GEN_2466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2468 = 7'h12 == r_count_23_io_out ? io_r_18_b : _GEN_2467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2469 = 7'h13 == r_count_23_io_out ? io_r_19_b : _GEN_2468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2470 = 7'h14 == r_count_23_io_out ? io_r_20_b : _GEN_2469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2471 = 7'h15 == r_count_23_io_out ? io_r_21_b : _GEN_2470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2472 = 7'h16 == r_count_23_io_out ? io_r_22_b : _GEN_2471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2473 = 7'h17 == r_count_23_io_out ? io_r_23_b : _GEN_2472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2474 = 7'h18 == r_count_23_io_out ? io_r_24_b : _GEN_2473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2475 = 7'h19 == r_count_23_io_out ? io_r_25_b : _GEN_2474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2476 = 7'h1a == r_count_23_io_out ? io_r_26_b : _GEN_2475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2477 = 7'h1b == r_count_23_io_out ? io_r_27_b : _GEN_2476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2478 = 7'h1c == r_count_23_io_out ? io_r_28_b : _GEN_2477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2479 = 7'h1d == r_count_23_io_out ? io_r_29_b : _GEN_2478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2480 = 7'h1e == r_count_23_io_out ? io_r_30_b : _GEN_2479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2481 = 7'h1f == r_count_23_io_out ? io_r_31_b : _GEN_2480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2482 = 7'h20 == r_count_23_io_out ? io_r_32_b : _GEN_2481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2483 = 7'h21 == r_count_23_io_out ? io_r_33_b : _GEN_2482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2484 = 7'h22 == r_count_23_io_out ? io_r_34_b : _GEN_2483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2485 = 7'h23 == r_count_23_io_out ? io_r_35_b : _GEN_2484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2486 = 7'h24 == r_count_23_io_out ? io_r_36_b : _GEN_2485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2487 = 7'h25 == r_count_23_io_out ? io_r_37_b : _GEN_2486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2488 = 7'h26 == r_count_23_io_out ? io_r_38_b : _GEN_2487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2489 = 7'h27 == r_count_23_io_out ? io_r_39_b : _GEN_2488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2490 = 7'h28 == r_count_23_io_out ? io_r_40_b : _GEN_2489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2491 = 7'h29 == r_count_23_io_out ? io_r_41_b : _GEN_2490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2492 = 7'h2a == r_count_23_io_out ? io_r_42_b : _GEN_2491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2493 = 7'h2b == r_count_23_io_out ? io_r_43_b : _GEN_2492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2494 = 7'h2c == r_count_23_io_out ? io_r_44_b : _GEN_2493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2495 = 7'h2d == r_count_23_io_out ? io_r_45_b : _GEN_2494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2496 = 7'h2e == r_count_23_io_out ? io_r_46_b : _GEN_2495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2497 = 7'h2f == r_count_23_io_out ? io_r_47_b : _GEN_2496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2498 = 7'h30 == r_count_23_io_out ? io_r_48_b : _GEN_2497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2499 = 7'h31 == r_count_23_io_out ? io_r_49_b : _GEN_2498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2500 = 7'h32 == r_count_23_io_out ? io_r_50_b : _GEN_2499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2501 = 7'h33 == r_count_23_io_out ? io_r_51_b : _GEN_2500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2502 = 7'h34 == r_count_23_io_out ? io_r_52_b : _GEN_2501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2503 = 7'h35 == r_count_23_io_out ? io_r_53_b : _GEN_2502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2504 = 7'h36 == r_count_23_io_out ? io_r_54_b : _GEN_2503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2505 = 7'h37 == r_count_23_io_out ? io_r_55_b : _GEN_2504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2506 = 7'h38 == r_count_23_io_out ? io_r_56_b : _GEN_2505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2507 = 7'h39 == r_count_23_io_out ? io_r_57_b : _GEN_2506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2508 = 7'h3a == r_count_23_io_out ? io_r_58_b : _GEN_2507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2509 = 7'h3b == r_count_23_io_out ? io_r_59_b : _GEN_2508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2510 = 7'h3c == r_count_23_io_out ? io_r_60_b : _GEN_2509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2511 = 7'h3d == r_count_23_io_out ? io_r_61_b : _GEN_2510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2512 = 7'h3e == r_count_23_io_out ? io_r_62_b : _GEN_2511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2513 = 7'h3f == r_count_23_io_out ? io_r_63_b : _GEN_2512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2514 = 7'h40 == r_count_23_io_out ? io_r_64_b : _GEN_2513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2515 = 7'h41 == r_count_23_io_out ? io_r_65_b : _GEN_2514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2516 = 7'h42 == r_count_23_io_out ? io_r_66_b : _GEN_2515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2517 = 7'h43 == r_count_23_io_out ? io_r_67_b : _GEN_2516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2518 = 7'h44 == r_count_23_io_out ? io_r_68_b : _GEN_2517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2519 = 7'h45 == r_count_23_io_out ? io_r_69_b : _GEN_2518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2520 = 7'h46 == r_count_23_io_out ? io_r_70_b : _GEN_2519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2521 = 7'h47 == r_count_23_io_out ? io_r_71_b : _GEN_2520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2522 = 7'h48 == r_count_23_io_out ? io_r_72_b : _GEN_2521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2523 = 7'h49 == r_count_23_io_out ? io_r_73_b : _GEN_2522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2524 = 7'h4a == r_count_23_io_out ? io_r_74_b : _GEN_2523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2525 = 7'h4b == r_count_23_io_out ? io_r_75_b : _GEN_2524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2526 = 7'h4c == r_count_23_io_out ? io_r_76_b : _GEN_2525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2527 = 7'h4d == r_count_23_io_out ? io_r_77_b : _GEN_2526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2528 = 7'h4e == r_count_23_io_out ? io_r_78_b : _GEN_2527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2529 = 7'h4f == r_count_23_io_out ? io_r_79_b : _GEN_2528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2530 = 7'h50 == r_count_23_io_out ? io_r_80_b : _GEN_2529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2531 = 7'h51 == r_count_23_io_out ? io_r_81_b : _GEN_2530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2532 = 7'h52 == r_count_23_io_out ? io_r_82_b : _GEN_2531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2533 = 7'h53 == r_count_23_io_out ? io_r_83_b : _GEN_2532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2534 = 7'h54 == r_count_23_io_out ? io_r_84_b : _GEN_2533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2535 = 7'h55 == r_count_23_io_out ? io_r_85_b : _GEN_2534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2536 = 7'h56 == r_count_23_io_out ? io_r_86_b : _GEN_2535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2537 = 7'h57 == r_count_23_io_out ? io_r_87_b : _GEN_2536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2538 = 7'h58 == r_count_23_io_out ? io_r_88_b : _GEN_2537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2539 = 7'h59 == r_count_23_io_out ? io_r_89_b : _GEN_2538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2540 = 7'h5a == r_count_23_io_out ? io_r_90_b : _GEN_2539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2541 = 7'h5b == r_count_23_io_out ? io_r_91_b : _GEN_2540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2542 = 7'h5c == r_count_23_io_out ? io_r_92_b : _GEN_2541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2543 = 7'h5d == r_count_23_io_out ? io_r_93_b : _GEN_2542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2544 = 7'h5e == r_count_23_io_out ? io_r_94_b : _GEN_2543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2545 = 7'h5f == r_count_23_io_out ? io_r_95_b : _GEN_2544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2546 = 7'h60 == r_count_23_io_out ? io_r_96_b : _GEN_2545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2547 = 7'h61 == r_count_23_io_out ? io_r_97_b : _GEN_2546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2548 = 7'h62 == r_count_23_io_out ? io_r_98_b : _GEN_2547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2551 = 7'h1 == r_count_24_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2552 = 7'h2 == r_count_24_io_out ? io_r_2_b : _GEN_2551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2553 = 7'h3 == r_count_24_io_out ? io_r_3_b : _GEN_2552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2554 = 7'h4 == r_count_24_io_out ? io_r_4_b : _GEN_2553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2555 = 7'h5 == r_count_24_io_out ? io_r_5_b : _GEN_2554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2556 = 7'h6 == r_count_24_io_out ? io_r_6_b : _GEN_2555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2557 = 7'h7 == r_count_24_io_out ? io_r_7_b : _GEN_2556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2558 = 7'h8 == r_count_24_io_out ? io_r_8_b : _GEN_2557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2559 = 7'h9 == r_count_24_io_out ? io_r_9_b : _GEN_2558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2560 = 7'ha == r_count_24_io_out ? io_r_10_b : _GEN_2559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2561 = 7'hb == r_count_24_io_out ? io_r_11_b : _GEN_2560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2562 = 7'hc == r_count_24_io_out ? io_r_12_b : _GEN_2561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2563 = 7'hd == r_count_24_io_out ? io_r_13_b : _GEN_2562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2564 = 7'he == r_count_24_io_out ? io_r_14_b : _GEN_2563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2565 = 7'hf == r_count_24_io_out ? io_r_15_b : _GEN_2564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2566 = 7'h10 == r_count_24_io_out ? io_r_16_b : _GEN_2565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2567 = 7'h11 == r_count_24_io_out ? io_r_17_b : _GEN_2566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2568 = 7'h12 == r_count_24_io_out ? io_r_18_b : _GEN_2567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2569 = 7'h13 == r_count_24_io_out ? io_r_19_b : _GEN_2568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2570 = 7'h14 == r_count_24_io_out ? io_r_20_b : _GEN_2569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2571 = 7'h15 == r_count_24_io_out ? io_r_21_b : _GEN_2570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2572 = 7'h16 == r_count_24_io_out ? io_r_22_b : _GEN_2571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2573 = 7'h17 == r_count_24_io_out ? io_r_23_b : _GEN_2572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2574 = 7'h18 == r_count_24_io_out ? io_r_24_b : _GEN_2573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2575 = 7'h19 == r_count_24_io_out ? io_r_25_b : _GEN_2574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2576 = 7'h1a == r_count_24_io_out ? io_r_26_b : _GEN_2575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2577 = 7'h1b == r_count_24_io_out ? io_r_27_b : _GEN_2576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2578 = 7'h1c == r_count_24_io_out ? io_r_28_b : _GEN_2577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2579 = 7'h1d == r_count_24_io_out ? io_r_29_b : _GEN_2578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2580 = 7'h1e == r_count_24_io_out ? io_r_30_b : _GEN_2579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2581 = 7'h1f == r_count_24_io_out ? io_r_31_b : _GEN_2580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2582 = 7'h20 == r_count_24_io_out ? io_r_32_b : _GEN_2581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2583 = 7'h21 == r_count_24_io_out ? io_r_33_b : _GEN_2582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2584 = 7'h22 == r_count_24_io_out ? io_r_34_b : _GEN_2583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2585 = 7'h23 == r_count_24_io_out ? io_r_35_b : _GEN_2584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2586 = 7'h24 == r_count_24_io_out ? io_r_36_b : _GEN_2585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2587 = 7'h25 == r_count_24_io_out ? io_r_37_b : _GEN_2586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2588 = 7'h26 == r_count_24_io_out ? io_r_38_b : _GEN_2587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2589 = 7'h27 == r_count_24_io_out ? io_r_39_b : _GEN_2588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2590 = 7'h28 == r_count_24_io_out ? io_r_40_b : _GEN_2589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2591 = 7'h29 == r_count_24_io_out ? io_r_41_b : _GEN_2590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2592 = 7'h2a == r_count_24_io_out ? io_r_42_b : _GEN_2591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2593 = 7'h2b == r_count_24_io_out ? io_r_43_b : _GEN_2592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2594 = 7'h2c == r_count_24_io_out ? io_r_44_b : _GEN_2593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2595 = 7'h2d == r_count_24_io_out ? io_r_45_b : _GEN_2594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2596 = 7'h2e == r_count_24_io_out ? io_r_46_b : _GEN_2595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2597 = 7'h2f == r_count_24_io_out ? io_r_47_b : _GEN_2596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2598 = 7'h30 == r_count_24_io_out ? io_r_48_b : _GEN_2597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2599 = 7'h31 == r_count_24_io_out ? io_r_49_b : _GEN_2598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2600 = 7'h32 == r_count_24_io_out ? io_r_50_b : _GEN_2599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2601 = 7'h33 == r_count_24_io_out ? io_r_51_b : _GEN_2600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2602 = 7'h34 == r_count_24_io_out ? io_r_52_b : _GEN_2601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2603 = 7'h35 == r_count_24_io_out ? io_r_53_b : _GEN_2602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2604 = 7'h36 == r_count_24_io_out ? io_r_54_b : _GEN_2603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2605 = 7'h37 == r_count_24_io_out ? io_r_55_b : _GEN_2604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2606 = 7'h38 == r_count_24_io_out ? io_r_56_b : _GEN_2605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2607 = 7'h39 == r_count_24_io_out ? io_r_57_b : _GEN_2606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2608 = 7'h3a == r_count_24_io_out ? io_r_58_b : _GEN_2607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2609 = 7'h3b == r_count_24_io_out ? io_r_59_b : _GEN_2608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2610 = 7'h3c == r_count_24_io_out ? io_r_60_b : _GEN_2609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2611 = 7'h3d == r_count_24_io_out ? io_r_61_b : _GEN_2610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2612 = 7'h3e == r_count_24_io_out ? io_r_62_b : _GEN_2611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2613 = 7'h3f == r_count_24_io_out ? io_r_63_b : _GEN_2612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2614 = 7'h40 == r_count_24_io_out ? io_r_64_b : _GEN_2613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2615 = 7'h41 == r_count_24_io_out ? io_r_65_b : _GEN_2614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2616 = 7'h42 == r_count_24_io_out ? io_r_66_b : _GEN_2615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2617 = 7'h43 == r_count_24_io_out ? io_r_67_b : _GEN_2616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2618 = 7'h44 == r_count_24_io_out ? io_r_68_b : _GEN_2617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2619 = 7'h45 == r_count_24_io_out ? io_r_69_b : _GEN_2618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2620 = 7'h46 == r_count_24_io_out ? io_r_70_b : _GEN_2619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2621 = 7'h47 == r_count_24_io_out ? io_r_71_b : _GEN_2620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2622 = 7'h48 == r_count_24_io_out ? io_r_72_b : _GEN_2621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2623 = 7'h49 == r_count_24_io_out ? io_r_73_b : _GEN_2622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2624 = 7'h4a == r_count_24_io_out ? io_r_74_b : _GEN_2623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2625 = 7'h4b == r_count_24_io_out ? io_r_75_b : _GEN_2624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2626 = 7'h4c == r_count_24_io_out ? io_r_76_b : _GEN_2625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2627 = 7'h4d == r_count_24_io_out ? io_r_77_b : _GEN_2626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2628 = 7'h4e == r_count_24_io_out ? io_r_78_b : _GEN_2627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2629 = 7'h4f == r_count_24_io_out ? io_r_79_b : _GEN_2628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2630 = 7'h50 == r_count_24_io_out ? io_r_80_b : _GEN_2629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2631 = 7'h51 == r_count_24_io_out ? io_r_81_b : _GEN_2630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2632 = 7'h52 == r_count_24_io_out ? io_r_82_b : _GEN_2631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2633 = 7'h53 == r_count_24_io_out ? io_r_83_b : _GEN_2632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2634 = 7'h54 == r_count_24_io_out ? io_r_84_b : _GEN_2633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2635 = 7'h55 == r_count_24_io_out ? io_r_85_b : _GEN_2634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2636 = 7'h56 == r_count_24_io_out ? io_r_86_b : _GEN_2635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2637 = 7'h57 == r_count_24_io_out ? io_r_87_b : _GEN_2636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2638 = 7'h58 == r_count_24_io_out ? io_r_88_b : _GEN_2637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2639 = 7'h59 == r_count_24_io_out ? io_r_89_b : _GEN_2638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2640 = 7'h5a == r_count_24_io_out ? io_r_90_b : _GEN_2639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2641 = 7'h5b == r_count_24_io_out ? io_r_91_b : _GEN_2640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2642 = 7'h5c == r_count_24_io_out ? io_r_92_b : _GEN_2641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2643 = 7'h5d == r_count_24_io_out ? io_r_93_b : _GEN_2642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2644 = 7'h5e == r_count_24_io_out ? io_r_94_b : _GEN_2643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2645 = 7'h5f == r_count_24_io_out ? io_r_95_b : _GEN_2644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2646 = 7'h60 == r_count_24_io_out ? io_r_96_b : _GEN_2645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2647 = 7'h61 == r_count_24_io_out ? io_r_97_b : _GEN_2646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2648 = 7'h62 == r_count_24_io_out ? io_r_98_b : _GEN_2647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2651 = 7'h1 == r_count_25_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2652 = 7'h2 == r_count_25_io_out ? io_r_2_b : _GEN_2651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2653 = 7'h3 == r_count_25_io_out ? io_r_3_b : _GEN_2652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2654 = 7'h4 == r_count_25_io_out ? io_r_4_b : _GEN_2653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2655 = 7'h5 == r_count_25_io_out ? io_r_5_b : _GEN_2654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2656 = 7'h6 == r_count_25_io_out ? io_r_6_b : _GEN_2655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2657 = 7'h7 == r_count_25_io_out ? io_r_7_b : _GEN_2656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2658 = 7'h8 == r_count_25_io_out ? io_r_8_b : _GEN_2657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2659 = 7'h9 == r_count_25_io_out ? io_r_9_b : _GEN_2658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2660 = 7'ha == r_count_25_io_out ? io_r_10_b : _GEN_2659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2661 = 7'hb == r_count_25_io_out ? io_r_11_b : _GEN_2660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2662 = 7'hc == r_count_25_io_out ? io_r_12_b : _GEN_2661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2663 = 7'hd == r_count_25_io_out ? io_r_13_b : _GEN_2662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2664 = 7'he == r_count_25_io_out ? io_r_14_b : _GEN_2663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2665 = 7'hf == r_count_25_io_out ? io_r_15_b : _GEN_2664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2666 = 7'h10 == r_count_25_io_out ? io_r_16_b : _GEN_2665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2667 = 7'h11 == r_count_25_io_out ? io_r_17_b : _GEN_2666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2668 = 7'h12 == r_count_25_io_out ? io_r_18_b : _GEN_2667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2669 = 7'h13 == r_count_25_io_out ? io_r_19_b : _GEN_2668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2670 = 7'h14 == r_count_25_io_out ? io_r_20_b : _GEN_2669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2671 = 7'h15 == r_count_25_io_out ? io_r_21_b : _GEN_2670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2672 = 7'h16 == r_count_25_io_out ? io_r_22_b : _GEN_2671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2673 = 7'h17 == r_count_25_io_out ? io_r_23_b : _GEN_2672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2674 = 7'h18 == r_count_25_io_out ? io_r_24_b : _GEN_2673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2675 = 7'h19 == r_count_25_io_out ? io_r_25_b : _GEN_2674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2676 = 7'h1a == r_count_25_io_out ? io_r_26_b : _GEN_2675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2677 = 7'h1b == r_count_25_io_out ? io_r_27_b : _GEN_2676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2678 = 7'h1c == r_count_25_io_out ? io_r_28_b : _GEN_2677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2679 = 7'h1d == r_count_25_io_out ? io_r_29_b : _GEN_2678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2680 = 7'h1e == r_count_25_io_out ? io_r_30_b : _GEN_2679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2681 = 7'h1f == r_count_25_io_out ? io_r_31_b : _GEN_2680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2682 = 7'h20 == r_count_25_io_out ? io_r_32_b : _GEN_2681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2683 = 7'h21 == r_count_25_io_out ? io_r_33_b : _GEN_2682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2684 = 7'h22 == r_count_25_io_out ? io_r_34_b : _GEN_2683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2685 = 7'h23 == r_count_25_io_out ? io_r_35_b : _GEN_2684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2686 = 7'h24 == r_count_25_io_out ? io_r_36_b : _GEN_2685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2687 = 7'h25 == r_count_25_io_out ? io_r_37_b : _GEN_2686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2688 = 7'h26 == r_count_25_io_out ? io_r_38_b : _GEN_2687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2689 = 7'h27 == r_count_25_io_out ? io_r_39_b : _GEN_2688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2690 = 7'h28 == r_count_25_io_out ? io_r_40_b : _GEN_2689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2691 = 7'h29 == r_count_25_io_out ? io_r_41_b : _GEN_2690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2692 = 7'h2a == r_count_25_io_out ? io_r_42_b : _GEN_2691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2693 = 7'h2b == r_count_25_io_out ? io_r_43_b : _GEN_2692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2694 = 7'h2c == r_count_25_io_out ? io_r_44_b : _GEN_2693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2695 = 7'h2d == r_count_25_io_out ? io_r_45_b : _GEN_2694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2696 = 7'h2e == r_count_25_io_out ? io_r_46_b : _GEN_2695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2697 = 7'h2f == r_count_25_io_out ? io_r_47_b : _GEN_2696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2698 = 7'h30 == r_count_25_io_out ? io_r_48_b : _GEN_2697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2699 = 7'h31 == r_count_25_io_out ? io_r_49_b : _GEN_2698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2700 = 7'h32 == r_count_25_io_out ? io_r_50_b : _GEN_2699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2701 = 7'h33 == r_count_25_io_out ? io_r_51_b : _GEN_2700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2702 = 7'h34 == r_count_25_io_out ? io_r_52_b : _GEN_2701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2703 = 7'h35 == r_count_25_io_out ? io_r_53_b : _GEN_2702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2704 = 7'h36 == r_count_25_io_out ? io_r_54_b : _GEN_2703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2705 = 7'h37 == r_count_25_io_out ? io_r_55_b : _GEN_2704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2706 = 7'h38 == r_count_25_io_out ? io_r_56_b : _GEN_2705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2707 = 7'h39 == r_count_25_io_out ? io_r_57_b : _GEN_2706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2708 = 7'h3a == r_count_25_io_out ? io_r_58_b : _GEN_2707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2709 = 7'h3b == r_count_25_io_out ? io_r_59_b : _GEN_2708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2710 = 7'h3c == r_count_25_io_out ? io_r_60_b : _GEN_2709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2711 = 7'h3d == r_count_25_io_out ? io_r_61_b : _GEN_2710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2712 = 7'h3e == r_count_25_io_out ? io_r_62_b : _GEN_2711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2713 = 7'h3f == r_count_25_io_out ? io_r_63_b : _GEN_2712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2714 = 7'h40 == r_count_25_io_out ? io_r_64_b : _GEN_2713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2715 = 7'h41 == r_count_25_io_out ? io_r_65_b : _GEN_2714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2716 = 7'h42 == r_count_25_io_out ? io_r_66_b : _GEN_2715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2717 = 7'h43 == r_count_25_io_out ? io_r_67_b : _GEN_2716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2718 = 7'h44 == r_count_25_io_out ? io_r_68_b : _GEN_2717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2719 = 7'h45 == r_count_25_io_out ? io_r_69_b : _GEN_2718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2720 = 7'h46 == r_count_25_io_out ? io_r_70_b : _GEN_2719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2721 = 7'h47 == r_count_25_io_out ? io_r_71_b : _GEN_2720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2722 = 7'h48 == r_count_25_io_out ? io_r_72_b : _GEN_2721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2723 = 7'h49 == r_count_25_io_out ? io_r_73_b : _GEN_2722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2724 = 7'h4a == r_count_25_io_out ? io_r_74_b : _GEN_2723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2725 = 7'h4b == r_count_25_io_out ? io_r_75_b : _GEN_2724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2726 = 7'h4c == r_count_25_io_out ? io_r_76_b : _GEN_2725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2727 = 7'h4d == r_count_25_io_out ? io_r_77_b : _GEN_2726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2728 = 7'h4e == r_count_25_io_out ? io_r_78_b : _GEN_2727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2729 = 7'h4f == r_count_25_io_out ? io_r_79_b : _GEN_2728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2730 = 7'h50 == r_count_25_io_out ? io_r_80_b : _GEN_2729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2731 = 7'h51 == r_count_25_io_out ? io_r_81_b : _GEN_2730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2732 = 7'h52 == r_count_25_io_out ? io_r_82_b : _GEN_2731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2733 = 7'h53 == r_count_25_io_out ? io_r_83_b : _GEN_2732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2734 = 7'h54 == r_count_25_io_out ? io_r_84_b : _GEN_2733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2735 = 7'h55 == r_count_25_io_out ? io_r_85_b : _GEN_2734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2736 = 7'h56 == r_count_25_io_out ? io_r_86_b : _GEN_2735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2737 = 7'h57 == r_count_25_io_out ? io_r_87_b : _GEN_2736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2738 = 7'h58 == r_count_25_io_out ? io_r_88_b : _GEN_2737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2739 = 7'h59 == r_count_25_io_out ? io_r_89_b : _GEN_2738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2740 = 7'h5a == r_count_25_io_out ? io_r_90_b : _GEN_2739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2741 = 7'h5b == r_count_25_io_out ? io_r_91_b : _GEN_2740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2742 = 7'h5c == r_count_25_io_out ? io_r_92_b : _GEN_2741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2743 = 7'h5d == r_count_25_io_out ? io_r_93_b : _GEN_2742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2744 = 7'h5e == r_count_25_io_out ? io_r_94_b : _GEN_2743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2745 = 7'h5f == r_count_25_io_out ? io_r_95_b : _GEN_2744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2746 = 7'h60 == r_count_25_io_out ? io_r_96_b : _GEN_2745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2747 = 7'h61 == r_count_25_io_out ? io_r_97_b : _GEN_2746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2748 = 7'h62 == r_count_25_io_out ? io_r_98_b : _GEN_2747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2751 = 7'h1 == r_count_26_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2752 = 7'h2 == r_count_26_io_out ? io_r_2_b : _GEN_2751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2753 = 7'h3 == r_count_26_io_out ? io_r_3_b : _GEN_2752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2754 = 7'h4 == r_count_26_io_out ? io_r_4_b : _GEN_2753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2755 = 7'h5 == r_count_26_io_out ? io_r_5_b : _GEN_2754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2756 = 7'h6 == r_count_26_io_out ? io_r_6_b : _GEN_2755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2757 = 7'h7 == r_count_26_io_out ? io_r_7_b : _GEN_2756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2758 = 7'h8 == r_count_26_io_out ? io_r_8_b : _GEN_2757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2759 = 7'h9 == r_count_26_io_out ? io_r_9_b : _GEN_2758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2760 = 7'ha == r_count_26_io_out ? io_r_10_b : _GEN_2759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2761 = 7'hb == r_count_26_io_out ? io_r_11_b : _GEN_2760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2762 = 7'hc == r_count_26_io_out ? io_r_12_b : _GEN_2761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2763 = 7'hd == r_count_26_io_out ? io_r_13_b : _GEN_2762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2764 = 7'he == r_count_26_io_out ? io_r_14_b : _GEN_2763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2765 = 7'hf == r_count_26_io_out ? io_r_15_b : _GEN_2764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2766 = 7'h10 == r_count_26_io_out ? io_r_16_b : _GEN_2765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2767 = 7'h11 == r_count_26_io_out ? io_r_17_b : _GEN_2766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2768 = 7'h12 == r_count_26_io_out ? io_r_18_b : _GEN_2767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2769 = 7'h13 == r_count_26_io_out ? io_r_19_b : _GEN_2768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2770 = 7'h14 == r_count_26_io_out ? io_r_20_b : _GEN_2769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2771 = 7'h15 == r_count_26_io_out ? io_r_21_b : _GEN_2770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2772 = 7'h16 == r_count_26_io_out ? io_r_22_b : _GEN_2771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2773 = 7'h17 == r_count_26_io_out ? io_r_23_b : _GEN_2772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2774 = 7'h18 == r_count_26_io_out ? io_r_24_b : _GEN_2773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2775 = 7'h19 == r_count_26_io_out ? io_r_25_b : _GEN_2774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2776 = 7'h1a == r_count_26_io_out ? io_r_26_b : _GEN_2775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2777 = 7'h1b == r_count_26_io_out ? io_r_27_b : _GEN_2776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2778 = 7'h1c == r_count_26_io_out ? io_r_28_b : _GEN_2777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2779 = 7'h1d == r_count_26_io_out ? io_r_29_b : _GEN_2778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2780 = 7'h1e == r_count_26_io_out ? io_r_30_b : _GEN_2779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2781 = 7'h1f == r_count_26_io_out ? io_r_31_b : _GEN_2780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2782 = 7'h20 == r_count_26_io_out ? io_r_32_b : _GEN_2781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2783 = 7'h21 == r_count_26_io_out ? io_r_33_b : _GEN_2782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2784 = 7'h22 == r_count_26_io_out ? io_r_34_b : _GEN_2783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2785 = 7'h23 == r_count_26_io_out ? io_r_35_b : _GEN_2784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2786 = 7'h24 == r_count_26_io_out ? io_r_36_b : _GEN_2785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2787 = 7'h25 == r_count_26_io_out ? io_r_37_b : _GEN_2786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2788 = 7'h26 == r_count_26_io_out ? io_r_38_b : _GEN_2787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2789 = 7'h27 == r_count_26_io_out ? io_r_39_b : _GEN_2788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2790 = 7'h28 == r_count_26_io_out ? io_r_40_b : _GEN_2789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2791 = 7'h29 == r_count_26_io_out ? io_r_41_b : _GEN_2790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2792 = 7'h2a == r_count_26_io_out ? io_r_42_b : _GEN_2791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2793 = 7'h2b == r_count_26_io_out ? io_r_43_b : _GEN_2792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2794 = 7'h2c == r_count_26_io_out ? io_r_44_b : _GEN_2793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2795 = 7'h2d == r_count_26_io_out ? io_r_45_b : _GEN_2794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2796 = 7'h2e == r_count_26_io_out ? io_r_46_b : _GEN_2795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2797 = 7'h2f == r_count_26_io_out ? io_r_47_b : _GEN_2796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2798 = 7'h30 == r_count_26_io_out ? io_r_48_b : _GEN_2797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2799 = 7'h31 == r_count_26_io_out ? io_r_49_b : _GEN_2798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2800 = 7'h32 == r_count_26_io_out ? io_r_50_b : _GEN_2799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2801 = 7'h33 == r_count_26_io_out ? io_r_51_b : _GEN_2800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2802 = 7'h34 == r_count_26_io_out ? io_r_52_b : _GEN_2801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2803 = 7'h35 == r_count_26_io_out ? io_r_53_b : _GEN_2802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2804 = 7'h36 == r_count_26_io_out ? io_r_54_b : _GEN_2803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2805 = 7'h37 == r_count_26_io_out ? io_r_55_b : _GEN_2804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2806 = 7'h38 == r_count_26_io_out ? io_r_56_b : _GEN_2805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2807 = 7'h39 == r_count_26_io_out ? io_r_57_b : _GEN_2806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2808 = 7'h3a == r_count_26_io_out ? io_r_58_b : _GEN_2807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2809 = 7'h3b == r_count_26_io_out ? io_r_59_b : _GEN_2808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2810 = 7'h3c == r_count_26_io_out ? io_r_60_b : _GEN_2809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2811 = 7'h3d == r_count_26_io_out ? io_r_61_b : _GEN_2810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2812 = 7'h3e == r_count_26_io_out ? io_r_62_b : _GEN_2811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2813 = 7'h3f == r_count_26_io_out ? io_r_63_b : _GEN_2812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2814 = 7'h40 == r_count_26_io_out ? io_r_64_b : _GEN_2813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2815 = 7'h41 == r_count_26_io_out ? io_r_65_b : _GEN_2814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2816 = 7'h42 == r_count_26_io_out ? io_r_66_b : _GEN_2815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2817 = 7'h43 == r_count_26_io_out ? io_r_67_b : _GEN_2816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2818 = 7'h44 == r_count_26_io_out ? io_r_68_b : _GEN_2817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2819 = 7'h45 == r_count_26_io_out ? io_r_69_b : _GEN_2818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2820 = 7'h46 == r_count_26_io_out ? io_r_70_b : _GEN_2819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2821 = 7'h47 == r_count_26_io_out ? io_r_71_b : _GEN_2820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2822 = 7'h48 == r_count_26_io_out ? io_r_72_b : _GEN_2821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2823 = 7'h49 == r_count_26_io_out ? io_r_73_b : _GEN_2822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2824 = 7'h4a == r_count_26_io_out ? io_r_74_b : _GEN_2823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2825 = 7'h4b == r_count_26_io_out ? io_r_75_b : _GEN_2824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2826 = 7'h4c == r_count_26_io_out ? io_r_76_b : _GEN_2825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2827 = 7'h4d == r_count_26_io_out ? io_r_77_b : _GEN_2826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2828 = 7'h4e == r_count_26_io_out ? io_r_78_b : _GEN_2827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2829 = 7'h4f == r_count_26_io_out ? io_r_79_b : _GEN_2828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2830 = 7'h50 == r_count_26_io_out ? io_r_80_b : _GEN_2829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2831 = 7'h51 == r_count_26_io_out ? io_r_81_b : _GEN_2830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2832 = 7'h52 == r_count_26_io_out ? io_r_82_b : _GEN_2831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2833 = 7'h53 == r_count_26_io_out ? io_r_83_b : _GEN_2832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2834 = 7'h54 == r_count_26_io_out ? io_r_84_b : _GEN_2833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2835 = 7'h55 == r_count_26_io_out ? io_r_85_b : _GEN_2834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2836 = 7'h56 == r_count_26_io_out ? io_r_86_b : _GEN_2835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2837 = 7'h57 == r_count_26_io_out ? io_r_87_b : _GEN_2836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2838 = 7'h58 == r_count_26_io_out ? io_r_88_b : _GEN_2837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2839 = 7'h59 == r_count_26_io_out ? io_r_89_b : _GEN_2838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2840 = 7'h5a == r_count_26_io_out ? io_r_90_b : _GEN_2839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2841 = 7'h5b == r_count_26_io_out ? io_r_91_b : _GEN_2840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2842 = 7'h5c == r_count_26_io_out ? io_r_92_b : _GEN_2841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2843 = 7'h5d == r_count_26_io_out ? io_r_93_b : _GEN_2842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2844 = 7'h5e == r_count_26_io_out ? io_r_94_b : _GEN_2843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2845 = 7'h5f == r_count_26_io_out ? io_r_95_b : _GEN_2844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2846 = 7'h60 == r_count_26_io_out ? io_r_96_b : _GEN_2845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2847 = 7'h61 == r_count_26_io_out ? io_r_97_b : _GEN_2846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2848 = 7'h62 == r_count_26_io_out ? io_r_98_b : _GEN_2847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2851 = 7'h1 == r_count_27_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2852 = 7'h2 == r_count_27_io_out ? io_r_2_b : _GEN_2851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2853 = 7'h3 == r_count_27_io_out ? io_r_3_b : _GEN_2852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2854 = 7'h4 == r_count_27_io_out ? io_r_4_b : _GEN_2853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2855 = 7'h5 == r_count_27_io_out ? io_r_5_b : _GEN_2854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2856 = 7'h6 == r_count_27_io_out ? io_r_6_b : _GEN_2855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2857 = 7'h7 == r_count_27_io_out ? io_r_7_b : _GEN_2856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2858 = 7'h8 == r_count_27_io_out ? io_r_8_b : _GEN_2857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2859 = 7'h9 == r_count_27_io_out ? io_r_9_b : _GEN_2858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2860 = 7'ha == r_count_27_io_out ? io_r_10_b : _GEN_2859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2861 = 7'hb == r_count_27_io_out ? io_r_11_b : _GEN_2860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2862 = 7'hc == r_count_27_io_out ? io_r_12_b : _GEN_2861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2863 = 7'hd == r_count_27_io_out ? io_r_13_b : _GEN_2862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2864 = 7'he == r_count_27_io_out ? io_r_14_b : _GEN_2863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2865 = 7'hf == r_count_27_io_out ? io_r_15_b : _GEN_2864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2866 = 7'h10 == r_count_27_io_out ? io_r_16_b : _GEN_2865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2867 = 7'h11 == r_count_27_io_out ? io_r_17_b : _GEN_2866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2868 = 7'h12 == r_count_27_io_out ? io_r_18_b : _GEN_2867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2869 = 7'h13 == r_count_27_io_out ? io_r_19_b : _GEN_2868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2870 = 7'h14 == r_count_27_io_out ? io_r_20_b : _GEN_2869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2871 = 7'h15 == r_count_27_io_out ? io_r_21_b : _GEN_2870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2872 = 7'h16 == r_count_27_io_out ? io_r_22_b : _GEN_2871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2873 = 7'h17 == r_count_27_io_out ? io_r_23_b : _GEN_2872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2874 = 7'h18 == r_count_27_io_out ? io_r_24_b : _GEN_2873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2875 = 7'h19 == r_count_27_io_out ? io_r_25_b : _GEN_2874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2876 = 7'h1a == r_count_27_io_out ? io_r_26_b : _GEN_2875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2877 = 7'h1b == r_count_27_io_out ? io_r_27_b : _GEN_2876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2878 = 7'h1c == r_count_27_io_out ? io_r_28_b : _GEN_2877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2879 = 7'h1d == r_count_27_io_out ? io_r_29_b : _GEN_2878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2880 = 7'h1e == r_count_27_io_out ? io_r_30_b : _GEN_2879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2881 = 7'h1f == r_count_27_io_out ? io_r_31_b : _GEN_2880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2882 = 7'h20 == r_count_27_io_out ? io_r_32_b : _GEN_2881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2883 = 7'h21 == r_count_27_io_out ? io_r_33_b : _GEN_2882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2884 = 7'h22 == r_count_27_io_out ? io_r_34_b : _GEN_2883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2885 = 7'h23 == r_count_27_io_out ? io_r_35_b : _GEN_2884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2886 = 7'h24 == r_count_27_io_out ? io_r_36_b : _GEN_2885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2887 = 7'h25 == r_count_27_io_out ? io_r_37_b : _GEN_2886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2888 = 7'h26 == r_count_27_io_out ? io_r_38_b : _GEN_2887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2889 = 7'h27 == r_count_27_io_out ? io_r_39_b : _GEN_2888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2890 = 7'h28 == r_count_27_io_out ? io_r_40_b : _GEN_2889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2891 = 7'h29 == r_count_27_io_out ? io_r_41_b : _GEN_2890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2892 = 7'h2a == r_count_27_io_out ? io_r_42_b : _GEN_2891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2893 = 7'h2b == r_count_27_io_out ? io_r_43_b : _GEN_2892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2894 = 7'h2c == r_count_27_io_out ? io_r_44_b : _GEN_2893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2895 = 7'h2d == r_count_27_io_out ? io_r_45_b : _GEN_2894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2896 = 7'h2e == r_count_27_io_out ? io_r_46_b : _GEN_2895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2897 = 7'h2f == r_count_27_io_out ? io_r_47_b : _GEN_2896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2898 = 7'h30 == r_count_27_io_out ? io_r_48_b : _GEN_2897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2899 = 7'h31 == r_count_27_io_out ? io_r_49_b : _GEN_2898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2900 = 7'h32 == r_count_27_io_out ? io_r_50_b : _GEN_2899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2901 = 7'h33 == r_count_27_io_out ? io_r_51_b : _GEN_2900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2902 = 7'h34 == r_count_27_io_out ? io_r_52_b : _GEN_2901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2903 = 7'h35 == r_count_27_io_out ? io_r_53_b : _GEN_2902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2904 = 7'h36 == r_count_27_io_out ? io_r_54_b : _GEN_2903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2905 = 7'h37 == r_count_27_io_out ? io_r_55_b : _GEN_2904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2906 = 7'h38 == r_count_27_io_out ? io_r_56_b : _GEN_2905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2907 = 7'h39 == r_count_27_io_out ? io_r_57_b : _GEN_2906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2908 = 7'h3a == r_count_27_io_out ? io_r_58_b : _GEN_2907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2909 = 7'h3b == r_count_27_io_out ? io_r_59_b : _GEN_2908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2910 = 7'h3c == r_count_27_io_out ? io_r_60_b : _GEN_2909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2911 = 7'h3d == r_count_27_io_out ? io_r_61_b : _GEN_2910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2912 = 7'h3e == r_count_27_io_out ? io_r_62_b : _GEN_2911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2913 = 7'h3f == r_count_27_io_out ? io_r_63_b : _GEN_2912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2914 = 7'h40 == r_count_27_io_out ? io_r_64_b : _GEN_2913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2915 = 7'h41 == r_count_27_io_out ? io_r_65_b : _GEN_2914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2916 = 7'h42 == r_count_27_io_out ? io_r_66_b : _GEN_2915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2917 = 7'h43 == r_count_27_io_out ? io_r_67_b : _GEN_2916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2918 = 7'h44 == r_count_27_io_out ? io_r_68_b : _GEN_2917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2919 = 7'h45 == r_count_27_io_out ? io_r_69_b : _GEN_2918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2920 = 7'h46 == r_count_27_io_out ? io_r_70_b : _GEN_2919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2921 = 7'h47 == r_count_27_io_out ? io_r_71_b : _GEN_2920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2922 = 7'h48 == r_count_27_io_out ? io_r_72_b : _GEN_2921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2923 = 7'h49 == r_count_27_io_out ? io_r_73_b : _GEN_2922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2924 = 7'h4a == r_count_27_io_out ? io_r_74_b : _GEN_2923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2925 = 7'h4b == r_count_27_io_out ? io_r_75_b : _GEN_2924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2926 = 7'h4c == r_count_27_io_out ? io_r_76_b : _GEN_2925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2927 = 7'h4d == r_count_27_io_out ? io_r_77_b : _GEN_2926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2928 = 7'h4e == r_count_27_io_out ? io_r_78_b : _GEN_2927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2929 = 7'h4f == r_count_27_io_out ? io_r_79_b : _GEN_2928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2930 = 7'h50 == r_count_27_io_out ? io_r_80_b : _GEN_2929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2931 = 7'h51 == r_count_27_io_out ? io_r_81_b : _GEN_2930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2932 = 7'h52 == r_count_27_io_out ? io_r_82_b : _GEN_2931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2933 = 7'h53 == r_count_27_io_out ? io_r_83_b : _GEN_2932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2934 = 7'h54 == r_count_27_io_out ? io_r_84_b : _GEN_2933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2935 = 7'h55 == r_count_27_io_out ? io_r_85_b : _GEN_2934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2936 = 7'h56 == r_count_27_io_out ? io_r_86_b : _GEN_2935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2937 = 7'h57 == r_count_27_io_out ? io_r_87_b : _GEN_2936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2938 = 7'h58 == r_count_27_io_out ? io_r_88_b : _GEN_2937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2939 = 7'h59 == r_count_27_io_out ? io_r_89_b : _GEN_2938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2940 = 7'h5a == r_count_27_io_out ? io_r_90_b : _GEN_2939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2941 = 7'h5b == r_count_27_io_out ? io_r_91_b : _GEN_2940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2942 = 7'h5c == r_count_27_io_out ? io_r_92_b : _GEN_2941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2943 = 7'h5d == r_count_27_io_out ? io_r_93_b : _GEN_2942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2944 = 7'h5e == r_count_27_io_out ? io_r_94_b : _GEN_2943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2945 = 7'h5f == r_count_27_io_out ? io_r_95_b : _GEN_2944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2946 = 7'h60 == r_count_27_io_out ? io_r_96_b : _GEN_2945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2947 = 7'h61 == r_count_27_io_out ? io_r_97_b : _GEN_2946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2948 = 7'h62 == r_count_27_io_out ? io_r_98_b : _GEN_2947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2951 = 7'h1 == r_count_28_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2952 = 7'h2 == r_count_28_io_out ? io_r_2_b : _GEN_2951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2953 = 7'h3 == r_count_28_io_out ? io_r_3_b : _GEN_2952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2954 = 7'h4 == r_count_28_io_out ? io_r_4_b : _GEN_2953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2955 = 7'h5 == r_count_28_io_out ? io_r_5_b : _GEN_2954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2956 = 7'h6 == r_count_28_io_out ? io_r_6_b : _GEN_2955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2957 = 7'h7 == r_count_28_io_out ? io_r_7_b : _GEN_2956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2958 = 7'h8 == r_count_28_io_out ? io_r_8_b : _GEN_2957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2959 = 7'h9 == r_count_28_io_out ? io_r_9_b : _GEN_2958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2960 = 7'ha == r_count_28_io_out ? io_r_10_b : _GEN_2959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2961 = 7'hb == r_count_28_io_out ? io_r_11_b : _GEN_2960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2962 = 7'hc == r_count_28_io_out ? io_r_12_b : _GEN_2961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2963 = 7'hd == r_count_28_io_out ? io_r_13_b : _GEN_2962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2964 = 7'he == r_count_28_io_out ? io_r_14_b : _GEN_2963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2965 = 7'hf == r_count_28_io_out ? io_r_15_b : _GEN_2964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2966 = 7'h10 == r_count_28_io_out ? io_r_16_b : _GEN_2965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2967 = 7'h11 == r_count_28_io_out ? io_r_17_b : _GEN_2966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2968 = 7'h12 == r_count_28_io_out ? io_r_18_b : _GEN_2967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2969 = 7'h13 == r_count_28_io_out ? io_r_19_b : _GEN_2968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2970 = 7'h14 == r_count_28_io_out ? io_r_20_b : _GEN_2969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2971 = 7'h15 == r_count_28_io_out ? io_r_21_b : _GEN_2970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2972 = 7'h16 == r_count_28_io_out ? io_r_22_b : _GEN_2971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2973 = 7'h17 == r_count_28_io_out ? io_r_23_b : _GEN_2972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2974 = 7'h18 == r_count_28_io_out ? io_r_24_b : _GEN_2973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2975 = 7'h19 == r_count_28_io_out ? io_r_25_b : _GEN_2974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2976 = 7'h1a == r_count_28_io_out ? io_r_26_b : _GEN_2975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2977 = 7'h1b == r_count_28_io_out ? io_r_27_b : _GEN_2976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2978 = 7'h1c == r_count_28_io_out ? io_r_28_b : _GEN_2977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2979 = 7'h1d == r_count_28_io_out ? io_r_29_b : _GEN_2978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2980 = 7'h1e == r_count_28_io_out ? io_r_30_b : _GEN_2979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2981 = 7'h1f == r_count_28_io_out ? io_r_31_b : _GEN_2980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2982 = 7'h20 == r_count_28_io_out ? io_r_32_b : _GEN_2981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2983 = 7'h21 == r_count_28_io_out ? io_r_33_b : _GEN_2982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2984 = 7'h22 == r_count_28_io_out ? io_r_34_b : _GEN_2983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2985 = 7'h23 == r_count_28_io_out ? io_r_35_b : _GEN_2984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2986 = 7'h24 == r_count_28_io_out ? io_r_36_b : _GEN_2985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2987 = 7'h25 == r_count_28_io_out ? io_r_37_b : _GEN_2986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2988 = 7'h26 == r_count_28_io_out ? io_r_38_b : _GEN_2987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2989 = 7'h27 == r_count_28_io_out ? io_r_39_b : _GEN_2988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2990 = 7'h28 == r_count_28_io_out ? io_r_40_b : _GEN_2989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2991 = 7'h29 == r_count_28_io_out ? io_r_41_b : _GEN_2990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2992 = 7'h2a == r_count_28_io_out ? io_r_42_b : _GEN_2991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2993 = 7'h2b == r_count_28_io_out ? io_r_43_b : _GEN_2992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2994 = 7'h2c == r_count_28_io_out ? io_r_44_b : _GEN_2993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2995 = 7'h2d == r_count_28_io_out ? io_r_45_b : _GEN_2994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2996 = 7'h2e == r_count_28_io_out ? io_r_46_b : _GEN_2995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2997 = 7'h2f == r_count_28_io_out ? io_r_47_b : _GEN_2996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2998 = 7'h30 == r_count_28_io_out ? io_r_48_b : _GEN_2997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_2999 = 7'h31 == r_count_28_io_out ? io_r_49_b : _GEN_2998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3000 = 7'h32 == r_count_28_io_out ? io_r_50_b : _GEN_2999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3001 = 7'h33 == r_count_28_io_out ? io_r_51_b : _GEN_3000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3002 = 7'h34 == r_count_28_io_out ? io_r_52_b : _GEN_3001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3003 = 7'h35 == r_count_28_io_out ? io_r_53_b : _GEN_3002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3004 = 7'h36 == r_count_28_io_out ? io_r_54_b : _GEN_3003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3005 = 7'h37 == r_count_28_io_out ? io_r_55_b : _GEN_3004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3006 = 7'h38 == r_count_28_io_out ? io_r_56_b : _GEN_3005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3007 = 7'h39 == r_count_28_io_out ? io_r_57_b : _GEN_3006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3008 = 7'h3a == r_count_28_io_out ? io_r_58_b : _GEN_3007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3009 = 7'h3b == r_count_28_io_out ? io_r_59_b : _GEN_3008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3010 = 7'h3c == r_count_28_io_out ? io_r_60_b : _GEN_3009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3011 = 7'h3d == r_count_28_io_out ? io_r_61_b : _GEN_3010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3012 = 7'h3e == r_count_28_io_out ? io_r_62_b : _GEN_3011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3013 = 7'h3f == r_count_28_io_out ? io_r_63_b : _GEN_3012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3014 = 7'h40 == r_count_28_io_out ? io_r_64_b : _GEN_3013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3015 = 7'h41 == r_count_28_io_out ? io_r_65_b : _GEN_3014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3016 = 7'h42 == r_count_28_io_out ? io_r_66_b : _GEN_3015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3017 = 7'h43 == r_count_28_io_out ? io_r_67_b : _GEN_3016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3018 = 7'h44 == r_count_28_io_out ? io_r_68_b : _GEN_3017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3019 = 7'h45 == r_count_28_io_out ? io_r_69_b : _GEN_3018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3020 = 7'h46 == r_count_28_io_out ? io_r_70_b : _GEN_3019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3021 = 7'h47 == r_count_28_io_out ? io_r_71_b : _GEN_3020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3022 = 7'h48 == r_count_28_io_out ? io_r_72_b : _GEN_3021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3023 = 7'h49 == r_count_28_io_out ? io_r_73_b : _GEN_3022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3024 = 7'h4a == r_count_28_io_out ? io_r_74_b : _GEN_3023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3025 = 7'h4b == r_count_28_io_out ? io_r_75_b : _GEN_3024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3026 = 7'h4c == r_count_28_io_out ? io_r_76_b : _GEN_3025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3027 = 7'h4d == r_count_28_io_out ? io_r_77_b : _GEN_3026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3028 = 7'h4e == r_count_28_io_out ? io_r_78_b : _GEN_3027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3029 = 7'h4f == r_count_28_io_out ? io_r_79_b : _GEN_3028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3030 = 7'h50 == r_count_28_io_out ? io_r_80_b : _GEN_3029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3031 = 7'h51 == r_count_28_io_out ? io_r_81_b : _GEN_3030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3032 = 7'h52 == r_count_28_io_out ? io_r_82_b : _GEN_3031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3033 = 7'h53 == r_count_28_io_out ? io_r_83_b : _GEN_3032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3034 = 7'h54 == r_count_28_io_out ? io_r_84_b : _GEN_3033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3035 = 7'h55 == r_count_28_io_out ? io_r_85_b : _GEN_3034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3036 = 7'h56 == r_count_28_io_out ? io_r_86_b : _GEN_3035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3037 = 7'h57 == r_count_28_io_out ? io_r_87_b : _GEN_3036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3038 = 7'h58 == r_count_28_io_out ? io_r_88_b : _GEN_3037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3039 = 7'h59 == r_count_28_io_out ? io_r_89_b : _GEN_3038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3040 = 7'h5a == r_count_28_io_out ? io_r_90_b : _GEN_3039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3041 = 7'h5b == r_count_28_io_out ? io_r_91_b : _GEN_3040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3042 = 7'h5c == r_count_28_io_out ? io_r_92_b : _GEN_3041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3043 = 7'h5d == r_count_28_io_out ? io_r_93_b : _GEN_3042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3044 = 7'h5e == r_count_28_io_out ? io_r_94_b : _GEN_3043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3045 = 7'h5f == r_count_28_io_out ? io_r_95_b : _GEN_3044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3046 = 7'h60 == r_count_28_io_out ? io_r_96_b : _GEN_3045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3047 = 7'h61 == r_count_28_io_out ? io_r_97_b : _GEN_3046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3048 = 7'h62 == r_count_28_io_out ? io_r_98_b : _GEN_3047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3051 = 7'h1 == r_count_29_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3052 = 7'h2 == r_count_29_io_out ? io_r_2_b : _GEN_3051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3053 = 7'h3 == r_count_29_io_out ? io_r_3_b : _GEN_3052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3054 = 7'h4 == r_count_29_io_out ? io_r_4_b : _GEN_3053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3055 = 7'h5 == r_count_29_io_out ? io_r_5_b : _GEN_3054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3056 = 7'h6 == r_count_29_io_out ? io_r_6_b : _GEN_3055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3057 = 7'h7 == r_count_29_io_out ? io_r_7_b : _GEN_3056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3058 = 7'h8 == r_count_29_io_out ? io_r_8_b : _GEN_3057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3059 = 7'h9 == r_count_29_io_out ? io_r_9_b : _GEN_3058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3060 = 7'ha == r_count_29_io_out ? io_r_10_b : _GEN_3059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3061 = 7'hb == r_count_29_io_out ? io_r_11_b : _GEN_3060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3062 = 7'hc == r_count_29_io_out ? io_r_12_b : _GEN_3061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3063 = 7'hd == r_count_29_io_out ? io_r_13_b : _GEN_3062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3064 = 7'he == r_count_29_io_out ? io_r_14_b : _GEN_3063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3065 = 7'hf == r_count_29_io_out ? io_r_15_b : _GEN_3064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3066 = 7'h10 == r_count_29_io_out ? io_r_16_b : _GEN_3065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3067 = 7'h11 == r_count_29_io_out ? io_r_17_b : _GEN_3066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3068 = 7'h12 == r_count_29_io_out ? io_r_18_b : _GEN_3067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3069 = 7'h13 == r_count_29_io_out ? io_r_19_b : _GEN_3068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3070 = 7'h14 == r_count_29_io_out ? io_r_20_b : _GEN_3069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3071 = 7'h15 == r_count_29_io_out ? io_r_21_b : _GEN_3070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3072 = 7'h16 == r_count_29_io_out ? io_r_22_b : _GEN_3071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3073 = 7'h17 == r_count_29_io_out ? io_r_23_b : _GEN_3072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3074 = 7'h18 == r_count_29_io_out ? io_r_24_b : _GEN_3073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3075 = 7'h19 == r_count_29_io_out ? io_r_25_b : _GEN_3074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3076 = 7'h1a == r_count_29_io_out ? io_r_26_b : _GEN_3075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3077 = 7'h1b == r_count_29_io_out ? io_r_27_b : _GEN_3076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3078 = 7'h1c == r_count_29_io_out ? io_r_28_b : _GEN_3077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3079 = 7'h1d == r_count_29_io_out ? io_r_29_b : _GEN_3078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3080 = 7'h1e == r_count_29_io_out ? io_r_30_b : _GEN_3079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3081 = 7'h1f == r_count_29_io_out ? io_r_31_b : _GEN_3080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3082 = 7'h20 == r_count_29_io_out ? io_r_32_b : _GEN_3081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3083 = 7'h21 == r_count_29_io_out ? io_r_33_b : _GEN_3082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3084 = 7'h22 == r_count_29_io_out ? io_r_34_b : _GEN_3083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3085 = 7'h23 == r_count_29_io_out ? io_r_35_b : _GEN_3084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3086 = 7'h24 == r_count_29_io_out ? io_r_36_b : _GEN_3085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3087 = 7'h25 == r_count_29_io_out ? io_r_37_b : _GEN_3086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3088 = 7'h26 == r_count_29_io_out ? io_r_38_b : _GEN_3087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3089 = 7'h27 == r_count_29_io_out ? io_r_39_b : _GEN_3088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3090 = 7'h28 == r_count_29_io_out ? io_r_40_b : _GEN_3089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3091 = 7'h29 == r_count_29_io_out ? io_r_41_b : _GEN_3090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3092 = 7'h2a == r_count_29_io_out ? io_r_42_b : _GEN_3091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3093 = 7'h2b == r_count_29_io_out ? io_r_43_b : _GEN_3092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3094 = 7'h2c == r_count_29_io_out ? io_r_44_b : _GEN_3093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3095 = 7'h2d == r_count_29_io_out ? io_r_45_b : _GEN_3094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3096 = 7'h2e == r_count_29_io_out ? io_r_46_b : _GEN_3095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3097 = 7'h2f == r_count_29_io_out ? io_r_47_b : _GEN_3096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3098 = 7'h30 == r_count_29_io_out ? io_r_48_b : _GEN_3097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3099 = 7'h31 == r_count_29_io_out ? io_r_49_b : _GEN_3098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3100 = 7'h32 == r_count_29_io_out ? io_r_50_b : _GEN_3099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3101 = 7'h33 == r_count_29_io_out ? io_r_51_b : _GEN_3100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3102 = 7'h34 == r_count_29_io_out ? io_r_52_b : _GEN_3101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3103 = 7'h35 == r_count_29_io_out ? io_r_53_b : _GEN_3102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3104 = 7'h36 == r_count_29_io_out ? io_r_54_b : _GEN_3103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3105 = 7'h37 == r_count_29_io_out ? io_r_55_b : _GEN_3104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3106 = 7'h38 == r_count_29_io_out ? io_r_56_b : _GEN_3105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3107 = 7'h39 == r_count_29_io_out ? io_r_57_b : _GEN_3106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3108 = 7'h3a == r_count_29_io_out ? io_r_58_b : _GEN_3107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3109 = 7'h3b == r_count_29_io_out ? io_r_59_b : _GEN_3108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3110 = 7'h3c == r_count_29_io_out ? io_r_60_b : _GEN_3109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3111 = 7'h3d == r_count_29_io_out ? io_r_61_b : _GEN_3110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3112 = 7'h3e == r_count_29_io_out ? io_r_62_b : _GEN_3111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3113 = 7'h3f == r_count_29_io_out ? io_r_63_b : _GEN_3112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3114 = 7'h40 == r_count_29_io_out ? io_r_64_b : _GEN_3113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3115 = 7'h41 == r_count_29_io_out ? io_r_65_b : _GEN_3114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3116 = 7'h42 == r_count_29_io_out ? io_r_66_b : _GEN_3115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3117 = 7'h43 == r_count_29_io_out ? io_r_67_b : _GEN_3116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3118 = 7'h44 == r_count_29_io_out ? io_r_68_b : _GEN_3117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3119 = 7'h45 == r_count_29_io_out ? io_r_69_b : _GEN_3118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3120 = 7'h46 == r_count_29_io_out ? io_r_70_b : _GEN_3119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3121 = 7'h47 == r_count_29_io_out ? io_r_71_b : _GEN_3120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3122 = 7'h48 == r_count_29_io_out ? io_r_72_b : _GEN_3121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3123 = 7'h49 == r_count_29_io_out ? io_r_73_b : _GEN_3122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3124 = 7'h4a == r_count_29_io_out ? io_r_74_b : _GEN_3123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3125 = 7'h4b == r_count_29_io_out ? io_r_75_b : _GEN_3124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3126 = 7'h4c == r_count_29_io_out ? io_r_76_b : _GEN_3125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3127 = 7'h4d == r_count_29_io_out ? io_r_77_b : _GEN_3126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3128 = 7'h4e == r_count_29_io_out ? io_r_78_b : _GEN_3127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3129 = 7'h4f == r_count_29_io_out ? io_r_79_b : _GEN_3128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3130 = 7'h50 == r_count_29_io_out ? io_r_80_b : _GEN_3129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3131 = 7'h51 == r_count_29_io_out ? io_r_81_b : _GEN_3130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3132 = 7'h52 == r_count_29_io_out ? io_r_82_b : _GEN_3131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3133 = 7'h53 == r_count_29_io_out ? io_r_83_b : _GEN_3132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3134 = 7'h54 == r_count_29_io_out ? io_r_84_b : _GEN_3133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3135 = 7'h55 == r_count_29_io_out ? io_r_85_b : _GEN_3134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3136 = 7'h56 == r_count_29_io_out ? io_r_86_b : _GEN_3135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3137 = 7'h57 == r_count_29_io_out ? io_r_87_b : _GEN_3136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3138 = 7'h58 == r_count_29_io_out ? io_r_88_b : _GEN_3137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3139 = 7'h59 == r_count_29_io_out ? io_r_89_b : _GEN_3138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3140 = 7'h5a == r_count_29_io_out ? io_r_90_b : _GEN_3139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3141 = 7'h5b == r_count_29_io_out ? io_r_91_b : _GEN_3140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3142 = 7'h5c == r_count_29_io_out ? io_r_92_b : _GEN_3141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3143 = 7'h5d == r_count_29_io_out ? io_r_93_b : _GEN_3142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3144 = 7'h5e == r_count_29_io_out ? io_r_94_b : _GEN_3143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3145 = 7'h5f == r_count_29_io_out ? io_r_95_b : _GEN_3144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3146 = 7'h60 == r_count_29_io_out ? io_r_96_b : _GEN_3145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3147 = 7'h61 == r_count_29_io_out ? io_r_97_b : _GEN_3146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3148 = 7'h62 == r_count_29_io_out ? io_r_98_b : _GEN_3147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3151 = 7'h1 == r_count_30_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3152 = 7'h2 == r_count_30_io_out ? io_r_2_b : _GEN_3151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3153 = 7'h3 == r_count_30_io_out ? io_r_3_b : _GEN_3152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3154 = 7'h4 == r_count_30_io_out ? io_r_4_b : _GEN_3153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3155 = 7'h5 == r_count_30_io_out ? io_r_5_b : _GEN_3154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3156 = 7'h6 == r_count_30_io_out ? io_r_6_b : _GEN_3155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3157 = 7'h7 == r_count_30_io_out ? io_r_7_b : _GEN_3156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3158 = 7'h8 == r_count_30_io_out ? io_r_8_b : _GEN_3157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3159 = 7'h9 == r_count_30_io_out ? io_r_9_b : _GEN_3158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3160 = 7'ha == r_count_30_io_out ? io_r_10_b : _GEN_3159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3161 = 7'hb == r_count_30_io_out ? io_r_11_b : _GEN_3160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3162 = 7'hc == r_count_30_io_out ? io_r_12_b : _GEN_3161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3163 = 7'hd == r_count_30_io_out ? io_r_13_b : _GEN_3162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3164 = 7'he == r_count_30_io_out ? io_r_14_b : _GEN_3163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3165 = 7'hf == r_count_30_io_out ? io_r_15_b : _GEN_3164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3166 = 7'h10 == r_count_30_io_out ? io_r_16_b : _GEN_3165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3167 = 7'h11 == r_count_30_io_out ? io_r_17_b : _GEN_3166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3168 = 7'h12 == r_count_30_io_out ? io_r_18_b : _GEN_3167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3169 = 7'h13 == r_count_30_io_out ? io_r_19_b : _GEN_3168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3170 = 7'h14 == r_count_30_io_out ? io_r_20_b : _GEN_3169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3171 = 7'h15 == r_count_30_io_out ? io_r_21_b : _GEN_3170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3172 = 7'h16 == r_count_30_io_out ? io_r_22_b : _GEN_3171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3173 = 7'h17 == r_count_30_io_out ? io_r_23_b : _GEN_3172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3174 = 7'h18 == r_count_30_io_out ? io_r_24_b : _GEN_3173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3175 = 7'h19 == r_count_30_io_out ? io_r_25_b : _GEN_3174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3176 = 7'h1a == r_count_30_io_out ? io_r_26_b : _GEN_3175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3177 = 7'h1b == r_count_30_io_out ? io_r_27_b : _GEN_3176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3178 = 7'h1c == r_count_30_io_out ? io_r_28_b : _GEN_3177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3179 = 7'h1d == r_count_30_io_out ? io_r_29_b : _GEN_3178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3180 = 7'h1e == r_count_30_io_out ? io_r_30_b : _GEN_3179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3181 = 7'h1f == r_count_30_io_out ? io_r_31_b : _GEN_3180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3182 = 7'h20 == r_count_30_io_out ? io_r_32_b : _GEN_3181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3183 = 7'h21 == r_count_30_io_out ? io_r_33_b : _GEN_3182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3184 = 7'h22 == r_count_30_io_out ? io_r_34_b : _GEN_3183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3185 = 7'h23 == r_count_30_io_out ? io_r_35_b : _GEN_3184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3186 = 7'h24 == r_count_30_io_out ? io_r_36_b : _GEN_3185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3187 = 7'h25 == r_count_30_io_out ? io_r_37_b : _GEN_3186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3188 = 7'h26 == r_count_30_io_out ? io_r_38_b : _GEN_3187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3189 = 7'h27 == r_count_30_io_out ? io_r_39_b : _GEN_3188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3190 = 7'h28 == r_count_30_io_out ? io_r_40_b : _GEN_3189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3191 = 7'h29 == r_count_30_io_out ? io_r_41_b : _GEN_3190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3192 = 7'h2a == r_count_30_io_out ? io_r_42_b : _GEN_3191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3193 = 7'h2b == r_count_30_io_out ? io_r_43_b : _GEN_3192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3194 = 7'h2c == r_count_30_io_out ? io_r_44_b : _GEN_3193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3195 = 7'h2d == r_count_30_io_out ? io_r_45_b : _GEN_3194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3196 = 7'h2e == r_count_30_io_out ? io_r_46_b : _GEN_3195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3197 = 7'h2f == r_count_30_io_out ? io_r_47_b : _GEN_3196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3198 = 7'h30 == r_count_30_io_out ? io_r_48_b : _GEN_3197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3199 = 7'h31 == r_count_30_io_out ? io_r_49_b : _GEN_3198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3200 = 7'h32 == r_count_30_io_out ? io_r_50_b : _GEN_3199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3201 = 7'h33 == r_count_30_io_out ? io_r_51_b : _GEN_3200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3202 = 7'h34 == r_count_30_io_out ? io_r_52_b : _GEN_3201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3203 = 7'h35 == r_count_30_io_out ? io_r_53_b : _GEN_3202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3204 = 7'h36 == r_count_30_io_out ? io_r_54_b : _GEN_3203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3205 = 7'h37 == r_count_30_io_out ? io_r_55_b : _GEN_3204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3206 = 7'h38 == r_count_30_io_out ? io_r_56_b : _GEN_3205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3207 = 7'h39 == r_count_30_io_out ? io_r_57_b : _GEN_3206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3208 = 7'h3a == r_count_30_io_out ? io_r_58_b : _GEN_3207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3209 = 7'h3b == r_count_30_io_out ? io_r_59_b : _GEN_3208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3210 = 7'h3c == r_count_30_io_out ? io_r_60_b : _GEN_3209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3211 = 7'h3d == r_count_30_io_out ? io_r_61_b : _GEN_3210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3212 = 7'h3e == r_count_30_io_out ? io_r_62_b : _GEN_3211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3213 = 7'h3f == r_count_30_io_out ? io_r_63_b : _GEN_3212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3214 = 7'h40 == r_count_30_io_out ? io_r_64_b : _GEN_3213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3215 = 7'h41 == r_count_30_io_out ? io_r_65_b : _GEN_3214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3216 = 7'h42 == r_count_30_io_out ? io_r_66_b : _GEN_3215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3217 = 7'h43 == r_count_30_io_out ? io_r_67_b : _GEN_3216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3218 = 7'h44 == r_count_30_io_out ? io_r_68_b : _GEN_3217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3219 = 7'h45 == r_count_30_io_out ? io_r_69_b : _GEN_3218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3220 = 7'h46 == r_count_30_io_out ? io_r_70_b : _GEN_3219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3221 = 7'h47 == r_count_30_io_out ? io_r_71_b : _GEN_3220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3222 = 7'h48 == r_count_30_io_out ? io_r_72_b : _GEN_3221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3223 = 7'h49 == r_count_30_io_out ? io_r_73_b : _GEN_3222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3224 = 7'h4a == r_count_30_io_out ? io_r_74_b : _GEN_3223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3225 = 7'h4b == r_count_30_io_out ? io_r_75_b : _GEN_3224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3226 = 7'h4c == r_count_30_io_out ? io_r_76_b : _GEN_3225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3227 = 7'h4d == r_count_30_io_out ? io_r_77_b : _GEN_3226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3228 = 7'h4e == r_count_30_io_out ? io_r_78_b : _GEN_3227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3229 = 7'h4f == r_count_30_io_out ? io_r_79_b : _GEN_3228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3230 = 7'h50 == r_count_30_io_out ? io_r_80_b : _GEN_3229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3231 = 7'h51 == r_count_30_io_out ? io_r_81_b : _GEN_3230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3232 = 7'h52 == r_count_30_io_out ? io_r_82_b : _GEN_3231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3233 = 7'h53 == r_count_30_io_out ? io_r_83_b : _GEN_3232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3234 = 7'h54 == r_count_30_io_out ? io_r_84_b : _GEN_3233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3235 = 7'h55 == r_count_30_io_out ? io_r_85_b : _GEN_3234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3236 = 7'h56 == r_count_30_io_out ? io_r_86_b : _GEN_3235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3237 = 7'h57 == r_count_30_io_out ? io_r_87_b : _GEN_3236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3238 = 7'h58 == r_count_30_io_out ? io_r_88_b : _GEN_3237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3239 = 7'h59 == r_count_30_io_out ? io_r_89_b : _GEN_3238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3240 = 7'h5a == r_count_30_io_out ? io_r_90_b : _GEN_3239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3241 = 7'h5b == r_count_30_io_out ? io_r_91_b : _GEN_3240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3242 = 7'h5c == r_count_30_io_out ? io_r_92_b : _GEN_3241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3243 = 7'h5d == r_count_30_io_out ? io_r_93_b : _GEN_3242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3244 = 7'h5e == r_count_30_io_out ? io_r_94_b : _GEN_3243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3245 = 7'h5f == r_count_30_io_out ? io_r_95_b : _GEN_3244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3246 = 7'h60 == r_count_30_io_out ? io_r_96_b : _GEN_3245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3247 = 7'h61 == r_count_30_io_out ? io_r_97_b : _GEN_3246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3248 = 7'h62 == r_count_30_io_out ? io_r_98_b : _GEN_3247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3251 = 7'h1 == r_count_31_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3252 = 7'h2 == r_count_31_io_out ? io_r_2_b : _GEN_3251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3253 = 7'h3 == r_count_31_io_out ? io_r_3_b : _GEN_3252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3254 = 7'h4 == r_count_31_io_out ? io_r_4_b : _GEN_3253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3255 = 7'h5 == r_count_31_io_out ? io_r_5_b : _GEN_3254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3256 = 7'h6 == r_count_31_io_out ? io_r_6_b : _GEN_3255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3257 = 7'h7 == r_count_31_io_out ? io_r_7_b : _GEN_3256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3258 = 7'h8 == r_count_31_io_out ? io_r_8_b : _GEN_3257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3259 = 7'h9 == r_count_31_io_out ? io_r_9_b : _GEN_3258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3260 = 7'ha == r_count_31_io_out ? io_r_10_b : _GEN_3259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3261 = 7'hb == r_count_31_io_out ? io_r_11_b : _GEN_3260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3262 = 7'hc == r_count_31_io_out ? io_r_12_b : _GEN_3261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3263 = 7'hd == r_count_31_io_out ? io_r_13_b : _GEN_3262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3264 = 7'he == r_count_31_io_out ? io_r_14_b : _GEN_3263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3265 = 7'hf == r_count_31_io_out ? io_r_15_b : _GEN_3264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3266 = 7'h10 == r_count_31_io_out ? io_r_16_b : _GEN_3265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3267 = 7'h11 == r_count_31_io_out ? io_r_17_b : _GEN_3266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3268 = 7'h12 == r_count_31_io_out ? io_r_18_b : _GEN_3267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3269 = 7'h13 == r_count_31_io_out ? io_r_19_b : _GEN_3268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3270 = 7'h14 == r_count_31_io_out ? io_r_20_b : _GEN_3269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3271 = 7'h15 == r_count_31_io_out ? io_r_21_b : _GEN_3270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3272 = 7'h16 == r_count_31_io_out ? io_r_22_b : _GEN_3271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3273 = 7'h17 == r_count_31_io_out ? io_r_23_b : _GEN_3272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3274 = 7'h18 == r_count_31_io_out ? io_r_24_b : _GEN_3273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3275 = 7'h19 == r_count_31_io_out ? io_r_25_b : _GEN_3274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3276 = 7'h1a == r_count_31_io_out ? io_r_26_b : _GEN_3275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3277 = 7'h1b == r_count_31_io_out ? io_r_27_b : _GEN_3276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3278 = 7'h1c == r_count_31_io_out ? io_r_28_b : _GEN_3277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3279 = 7'h1d == r_count_31_io_out ? io_r_29_b : _GEN_3278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3280 = 7'h1e == r_count_31_io_out ? io_r_30_b : _GEN_3279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3281 = 7'h1f == r_count_31_io_out ? io_r_31_b : _GEN_3280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3282 = 7'h20 == r_count_31_io_out ? io_r_32_b : _GEN_3281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3283 = 7'h21 == r_count_31_io_out ? io_r_33_b : _GEN_3282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3284 = 7'h22 == r_count_31_io_out ? io_r_34_b : _GEN_3283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3285 = 7'h23 == r_count_31_io_out ? io_r_35_b : _GEN_3284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3286 = 7'h24 == r_count_31_io_out ? io_r_36_b : _GEN_3285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3287 = 7'h25 == r_count_31_io_out ? io_r_37_b : _GEN_3286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3288 = 7'h26 == r_count_31_io_out ? io_r_38_b : _GEN_3287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3289 = 7'h27 == r_count_31_io_out ? io_r_39_b : _GEN_3288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3290 = 7'h28 == r_count_31_io_out ? io_r_40_b : _GEN_3289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3291 = 7'h29 == r_count_31_io_out ? io_r_41_b : _GEN_3290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3292 = 7'h2a == r_count_31_io_out ? io_r_42_b : _GEN_3291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3293 = 7'h2b == r_count_31_io_out ? io_r_43_b : _GEN_3292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3294 = 7'h2c == r_count_31_io_out ? io_r_44_b : _GEN_3293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3295 = 7'h2d == r_count_31_io_out ? io_r_45_b : _GEN_3294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3296 = 7'h2e == r_count_31_io_out ? io_r_46_b : _GEN_3295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3297 = 7'h2f == r_count_31_io_out ? io_r_47_b : _GEN_3296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3298 = 7'h30 == r_count_31_io_out ? io_r_48_b : _GEN_3297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3299 = 7'h31 == r_count_31_io_out ? io_r_49_b : _GEN_3298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3300 = 7'h32 == r_count_31_io_out ? io_r_50_b : _GEN_3299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3301 = 7'h33 == r_count_31_io_out ? io_r_51_b : _GEN_3300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3302 = 7'h34 == r_count_31_io_out ? io_r_52_b : _GEN_3301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3303 = 7'h35 == r_count_31_io_out ? io_r_53_b : _GEN_3302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3304 = 7'h36 == r_count_31_io_out ? io_r_54_b : _GEN_3303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3305 = 7'h37 == r_count_31_io_out ? io_r_55_b : _GEN_3304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3306 = 7'h38 == r_count_31_io_out ? io_r_56_b : _GEN_3305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3307 = 7'h39 == r_count_31_io_out ? io_r_57_b : _GEN_3306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3308 = 7'h3a == r_count_31_io_out ? io_r_58_b : _GEN_3307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3309 = 7'h3b == r_count_31_io_out ? io_r_59_b : _GEN_3308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3310 = 7'h3c == r_count_31_io_out ? io_r_60_b : _GEN_3309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3311 = 7'h3d == r_count_31_io_out ? io_r_61_b : _GEN_3310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3312 = 7'h3e == r_count_31_io_out ? io_r_62_b : _GEN_3311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3313 = 7'h3f == r_count_31_io_out ? io_r_63_b : _GEN_3312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3314 = 7'h40 == r_count_31_io_out ? io_r_64_b : _GEN_3313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3315 = 7'h41 == r_count_31_io_out ? io_r_65_b : _GEN_3314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3316 = 7'h42 == r_count_31_io_out ? io_r_66_b : _GEN_3315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3317 = 7'h43 == r_count_31_io_out ? io_r_67_b : _GEN_3316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3318 = 7'h44 == r_count_31_io_out ? io_r_68_b : _GEN_3317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3319 = 7'h45 == r_count_31_io_out ? io_r_69_b : _GEN_3318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3320 = 7'h46 == r_count_31_io_out ? io_r_70_b : _GEN_3319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3321 = 7'h47 == r_count_31_io_out ? io_r_71_b : _GEN_3320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3322 = 7'h48 == r_count_31_io_out ? io_r_72_b : _GEN_3321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3323 = 7'h49 == r_count_31_io_out ? io_r_73_b : _GEN_3322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3324 = 7'h4a == r_count_31_io_out ? io_r_74_b : _GEN_3323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3325 = 7'h4b == r_count_31_io_out ? io_r_75_b : _GEN_3324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3326 = 7'h4c == r_count_31_io_out ? io_r_76_b : _GEN_3325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3327 = 7'h4d == r_count_31_io_out ? io_r_77_b : _GEN_3326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3328 = 7'h4e == r_count_31_io_out ? io_r_78_b : _GEN_3327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3329 = 7'h4f == r_count_31_io_out ? io_r_79_b : _GEN_3328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3330 = 7'h50 == r_count_31_io_out ? io_r_80_b : _GEN_3329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3331 = 7'h51 == r_count_31_io_out ? io_r_81_b : _GEN_3330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3332 = 7'h52 == r_count_31_io_out ? io_r_82_b : _GEN_3331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3333 = 7'h53 == r_count_31_io_out ? io_r_83_b : _GEN_3332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3334 = 7'h54 == r_count_31_io_out ? io_r_84_b : _GEN_3333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3335 = 7'h55 == r_count_31_io_out ? io_r_85_b : _GEN_3334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3336 = 7'h56 == r_count_31_io_out ? io_r_86_b : _GEN_3335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3337 = 7'h57 == r_count_31_io_out ? io_r_87_b : _GEN_3336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3338 = 7'h58 == r_count_31_io_out ? io_r_88_b : _GEN_3337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3339 = 7'h59 == r_count_31_io_out ? io_r_89_b : _GEN_3338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3340 = 7'h5a == r_count_31_io_out ? io_r_90_b : _GEN_3339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3341 = 7'h5b == r_count_31_io_out ? io_r_91_b : _GEN_3340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3342 = 7'h5c == r_count_31_io_out ? io_r_92_b : _GEN_3341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3343 = 7'h5d == r_count_31_io_out ? io_r_93_b : _GEN_3342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3344 = 7'h5e == r_count_31_io_out ? io_r_94_b : _GEN_3343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3345 = 7'h5f == r_count_31_io_out ? io_r_95_b : _GEN_3344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3346 = 7'h60 == r_count_31_io_out ? io_r_96_b : _GEN_3345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3347 = 7'h61 == r_count_31_io_out ? io_r_97_b : _GEN_3346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3348 = 7'h62 == r_count_31_io_out ? io_r_98_b : _GEN_3347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3351 = 7'h1 == r_count_32_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3352 = 7'h2 == r_count_32_io_out ? io_r_2_b : _GEN_3351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3353 = 7'h3 == r_count_32_io_out ? io_r_3_b : _GEN_3352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3354 = 7'h4 == r_count_32_io_out ? io_r_4_b : _GEN_3353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3355 = 7'h5 == r_count_32_io_out ? io_r_5_b : _GEN_3354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3356 = 7'h6 == r_count_32_io_out ? io_r_6_b : _GEN_3355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3357 = 7'h7 == r_count_32_io_out ? io_r_7_b : _GEN_3356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3358 = 7'h8 == r_count_32_io_out ? io_r_8_b : _GEN_3357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3359 = 7'h9 == r_count_32_io_out ? io_r_9_b : _GEN_3358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3360 = 7'ha == r_count_32_io_out ? io_r_10_b : _GEN_3359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3361 = 7'hb == r_count_32_io_out ? io_r_11_b : _GEN_3360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3362 = 7'hc == r_count_32_io_out ? io_r_12_b : _GEN_3361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3363 = 7'hd == r_count_32_io_out ? io_r_13_b : _GEN_3362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3364 = 7'he == r_count_32_io_out ? io_r_14_b : _GEN_3363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3365 = 7'hf == r_count_32_io_out ? io_r_15_b : _GEN_3364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3366 = 7'h10 == r_count_32_io_out ? io_r_16_b : _GEN_3365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3367 = 7'h11 == r_count_32_io_out ? io_r_17_b : _GEN_3366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3368 = 7'h12 == r_count_32_io_out ? io_r_18_b : _GEN_3367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3369 = 7'h13 == r_count_32_io_out ? io_r_19_b : _GEN_3368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3370 = 7'h14 == r_count_32_io_out ? io_r_20_b : _GEN_3369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3371 = 7'h15 == r_count_32_io_out ? io_r_21_b : _GEN_3370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3372 = 7'h16 == r_count_32_io_out ? io_r_22_b : _GEN_3371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3373 = 7'h17 == r_count_32_io_out ? io_r_23_b : _GEN_3372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3374 = 7'h18 == r_count_32_io_out ? io_r_24_b : _GEN_3373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3375 = 7'h19 == r_count_32_io_out ? io_r_25_b : _GEN_3374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3376 = 7'h1a == r_count_32_io_out ? io_r_26_b : _GEN_3375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3377 = 7'h1b == r_count_32_io_out ? io_r_27_b : _GEN_3376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3378 = 7'h1c == r_count_32_io_out ? io_r_28_b : _GEN_3377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3379 = 7'h1d == r_count_32_io_out ? io_r_29_b : _GEN_3378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3380 = 7'h1e == r_count_32_io_out ? io_r_30_b : _GEN_3379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3381 = 7'h1f == r_count_32_io_out ? io_r_31_b : _GEN_3380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3382 = 7'h20 == r_count_32_io_out ? io_r_32_b : _GEN_3381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3383 = 7'h21 == r_count_32_io_out ? io_r_33_b : _GEN_3382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3384 = 7'h22 == r_count_32_io_out ? io_r_34_b : _GEN_3383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3385 = 7'h23 == r_count_32_io_out ? io_r_35_b : _GEN_3384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3386 = 7'h24 == r_count_32_io_out ? io_r_36_b : _GEN_3385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3387 = 7'h25 == r_count_32_io_out ? io_r_37_b : _GEN_3386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3388 = 7'h26 == r_count_32_io_out ? io_r_38_b : _GEN_3387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3389 = 7'h27 == r_count_32_io_out ? io_r_39_b : _GEN_3388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3390 = 7'h28 == r_count_32_io_out ? io_r_40_b : _GEN_3389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3391 = 7'h29 == r_count_32_io_out ? io_r_41_b : _GEN_3390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3392 = 7'h2a == r_count_32_io_out ? io_r_42_b : _GEN_3391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3393 = 7'h2b == r_count_32_io_out ? io_r_43_b : _GEN_3392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3394 = 7'h2c == r_count_32_io_out ? io_r_44_b : _GEN_3393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3395 = 7'h2d == r_count_32_io_out ? io_r_45_b : _GEN_3394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3396 = 7'h2e == r_count_32_io_out ? io_r_46_b : _GEN_3395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3397 = 7'h2f == r_count_32_io_out ? io_r_47_b : _GEN_3396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3398 = 7'h30 == r_count_32_io_out ? io_r_48_b : _GEN_3397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3399 = 7'h31 == r_count_32_io_out ? io_r_49_b : _GEN_3398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3400 = 7'h32 == r_count_32_io_out ? io_r_50_b : _GEN_3399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3401 = 7'h33 == r_count_32_io_out ? io_r_51_b : _GEN_3400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3402 = 7'h34 == r_count_32_io_out ? io_r_52_b : _GEN_3401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3403 = 7'h35 == r_count_32_io_out ? io_r_53_b : _GEN_3402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3404 = 7'h36 == r_count_32_io_out ? io_r_54_b : _GEN_3403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3405 = 7'h37 == r_count_32_io_out ? io_r_55_b : _GEN_3404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3406 = 7'h38 == r_count_32_io_out ? io_r_56_b : _GEN_3405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3407 = 7'h39 == r_count_32_io_out ? io_r_57_b : _GEN_3406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3408 = 7'h3a == r_count_32_io_out ? io_r_58_b : _GEN_3407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3409 = 7'h3b == r_count_32_io_out ? io_r_59_b : _GEN_3408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3410 = 7'h3c == r_count_32_io_out ? io_r_60_b : _GEN_3409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3411 = 7'h3d == r_count_32_io_out ? io_r_61_b : _GEN_3410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3412 = 7'h3e == r_count_32_io_out ? io_r_62_b : _GEN_3411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3413 = 7'h3f == r_count_32_io_out ? io_r_63_b : _GEN_3412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3414 = 7'h40 == r_count_32_io_out ? io_r_64_b : _GEN_3413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3415 = 7'h41 == r_count_32_io_out ? io_r_65_b : _GEN_3414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3416 = 7'h42 == r_count_32_io_out ? io_r_66_b : _GEN_3415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3417 = 7'h43 == r_count_32_io_out ? io_r_67_b : _GEN_3416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3418 = 7'h44 == r_count_32_io_out ? io_r_68_b : _GEN_3417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3419 = 7'h45 == r_count_32_io_out ? io_r_69_b : _GEN_3418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3420 = 7'h46 == r_count_32_io_out ? io_r_70_b : _GEN_3419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3421 = 7'h47 == r_count_32_io_out ? io_r_71_b : _GEN_3420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3422 = 7'h48 == r_count_32_io_out ? io_r_72_b : _GEN_3421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3423 = 7'h49 == r_count_32_io_out ? io_r_73_b : _GEN_3422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3424 = 7'h4a == r_count_32_io_out ? io_r_74_b : _GEN_3423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3425 = 7'h4b == r_count_32_io_out ? io_r_75_b : _GEN_3424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3426 = 7'h4c == r_count_32_io_out ? io_r_76_b : _GEN_3425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3427 = 7'h4d == r_count_32_io_out ? io_r_77_b : _GEN_3426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3428 = 7'h4e == r_count_32_io_out ? io_r_78_b : _GEN_3427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3429 = 7'h4f == r_count_32_io_out ? io_r_79_b : _GEN_3428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3430 = 7'h50 == r_count_32_io_out ? io_r_80_b : _GEN_3429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3431 = 7'h51 == r_count_32_io_out ? io_r_81_b : _GEN_3430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3432 = 7'h52 == r_count_32_io_out ? io_r_82_b : _GEN_3431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3433 = 7'h53 == r_count_32_io_out ? io_r_83_b : _GEN_3432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3434 = 7'h54 == r_count_32_io_out ? io_r_84_b : _GEN_3433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3435 = 7'h55 == r_count_32_io_out ? io_r_85_b : _GEN_3434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3436 = 7'h56 == r_count_32_io_out ? io_r_86_b : _GEN_3435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3437 = 7'h57 == r_count_32_io_out ? io_r_87_b : _GEN_3436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3438 = 7'h58 == r_count_32_io_out ? io_r_88_b : _GEN_3437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3439 = 7'h59 == r_count_32_io_out ? io_r_89_b : _GEN_3438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3440 = 7'h5a == r_count_32_io_out ? io_r_90_b : _GEN_3439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3441 = 7'h5b == r_count_32_io_out ? io_r_91_b : _GEN_3440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3442 = 7'h5c == r_count_32_io_out ? io_r_92_b : _GEN_3441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3443 = 7'h5d == r_count_32_io_out ? io_r_93_b : _GEN_3442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3444 = 7'h5e == r_count_32_io_out ? io_r_94_b : _GEN_3443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3445 = 7'h5f == r_count_32_io_out ? io_r_95_b : _GEN_3444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3446 = 7'h60 == r_count_32_io_out ? io_r_96_b : _GEN_3445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3447 = 7'h61 == r_count_32_io_out ? io_r_97_b : _GEN_3446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3448 = 7'h62 == r_count_32_io_out ? io_r_98_b : _GEN_3447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3451 = 7'h1 == r_count_33_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3452 = 7'h2 == r_count_33_io_out ? io_r_2_b : _GEN_3451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3453 = 7'h3 == r_count_33_io_out ? io_r_3_b : _GEN_3452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3454 = 7'h4 == r_count_33_io_out ? io_r_4_b : _GEN_3453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3455 = 7'h5 == r_count_33_io_out ? io_r_5_b : _GEN_3454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3456 = 7'h6 == r_count_33_io_out ? io_r_6_b : _GEN_3455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3457 = 7'h7 == r_count_33_io_out ? io_r_7_b : _GEN_3456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3458 = 7'h8 == r_count_33_io_out ? io_r_8_b : _GEN_3457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3459 = 7'h9 == r_count_33_io_out ? io_r_9_b : _GEN_3458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3460 = 7'ha == r_count_33_io_out ? io_r_10_b : _GEN_3459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3461 = 7'hb == r_count_33_io_out ? io_r_11_b : _GEN_3460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3462 = 7'hc == r_count_33_io_out ? io_r_12_b : _GEN_3461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3463 = 7'hd == r_count_33_io_out ? io_r_13_b : _GEN_3462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3464 = 7'he == r_count_33_io_out ? io_r_14_b : _GEN_3463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3465 = 7'hf == r_count_33_io_out ? io_r_15_b : _GEN_3464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3466 = 7'h10 == r_count_33_io_out ? io_r_16_b : _GEN_3465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3467 = 7'h11 == r_count_33_io_out ? io_r_17_b : _GEN_3466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3468 = 7'h12 == r_count_33_io_out ? io_r_18_b : _GEN_3467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3469 = 7'h13 == r_count_33_io_out ? io_r_19_b : _GEN_3468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3470 = 7'h14 == r_count_33_io_out ? io_r_20_b : _GEN_3469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3471 = 7'h15 == r_count_33_io_out ? io_r_21_b : _GEN_3470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3472 = 7'h16 == r_count_33_io_out ? io_r_22_b : _GEN_3471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3473 = 7'h17 == r_count_33_io_out ? io_r_23_b : _GEN_3472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3474 = 7'h18 == r_count_33_io_out ? io_r_24_b : _GEN_3473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3475 = 7'h19 == r_count_33_io_out ? io_r_25_b : _GEN_3474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3476 = 7'h1a == r_count_33_io_out ? io_r_26_b : _GEN_3475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3477 = 7'h1b == r_count_33_io_out ? io_r_27_b : _GEN_3476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3478 = 7'h1c == r_count_33_io_out ? io_r_28_b : _GEN_3477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3479 = 7'h1d == r_count_33_io_out ? io_r_29_b : _GEN_3478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3480 = 7'h1e == r_count_33_io_out ? io_r_30_b : _GEN_3479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3481 = 7'h1f == r_count_33_io_out ? io_r_31_b : _GEN_3480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3482 = 7'h20 == r_count_33_io_out ? io_r_32_b : _GEN_3481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3483 = 7'h21 == r_count_33_io_out ? io_r_33_b : _GEN_3482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3484 = 7'h22 == r_count_33_io_out ? io_r_34_b : _GEN_3483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3485 = 7'h23 == r_count_33_io_out ? io_r_35_b : _GEN_3484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3486 = 7'h24 == r_count_33_io_out ? io_r_36_b : _GEN_3485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3487 = 7'h25 == r_count_33_io_out ? io_r_37_b : _GEN_3486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3488 = 7'h26 == r_count_33_io_out ? io_r_38_b : _GEN_3487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3489 = 7'h27 == r_count_33_io_out ? io_r_39_b : _GEN_3488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3490 = 7'h28 == r_count_33_io_out ? io_r_40_b : _GEN_3489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3491 = 7'h29 == r_count_33_io_out ? io_r_41_b : _GEN_3490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3492 = 7'h2a == r_count_33_io_out ? io_r_42_b : _GEN_3491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3493 = 7'h2b == r_count_33_io_out ? io_r_43_b : _GEN_3492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3494 = 7'h2c == r_count_33_io_out ? io_r_44_b : _GEN_3493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3495 = 7'h2d == r_count_33_io_out ? io_r_45_b : _GEN_3494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3496 = 7'h2e == r_count_33_io_out ? io_r_46_b : _GEN_3495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3497 = 7'h2f == r_count_33_io_out ? io_r_47_b : _GEN_3496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3498 = 7'h30 == r_count_33_io_out ? io_r_48_b : _GEN_3497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3499 = 7'h31 == r_count_33_io_out ? io_r_49_b : _GEN_3498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3500 = 7'h32 == r_count_33_io_out ? io_r_50_b : _GEN_3499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3501 = 7'h33 == r_count_33_io_out ? io_r_51_b : _GEN_3500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3502 = 7'h34 == r_count_33_io_out ? io_r_52_b : _GEN_3501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3503 = 7'h35 == r_count_33_io_out ? io_r_53_b : _GEN_3502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3504 = 7'h36 == r_count_33_io_out ? io_r_54_b : _GEN_3503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3505 = 7'h37 == r_count_33_io_out ? io_r_55_b : _GEN_3504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3506 = 7'h38 == r_count_33_io_out ? io_r_56_b : _GEN_3505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3507 = 7'h39 == r_count_33_io_out ? io_r_57_b : _GEN_3506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3508 = 7'h3a == r_count_33_io_out ? io_r_58_b : _GEN_3507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3509 = 7'h3b == r_count_33_io_out ? io_r_59_b : _GEN_3508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3510 = 7'h3c == r_count_33_io_out ? io_r_60_b : _GEN_3509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3511 = 7'h3d == r_count_33_io_out ? io_r_61_b : _GEN_3510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3512 = 7'h3e == r_count_33_io_out ? io_r_62_b : _GEN_3511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3513 = 7'h3f == r_count_33_io_out ? io_r_63_b : _GEN_3512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3514 = 7'h40 == r_count_33_io_out ? io_r_64_b : _GEN_3513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3515 = 7'h41 == r_count_33_io_out ? io_r_65_b : _GEN_3514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3516 = 7'h42 == r_count_33_io_out ? io_r_66_b : _GEN_3515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3517 = 7'h43 == r_count_33_io_out ? io_r_67_b : _GEN_3516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3518 = 7'h44 == r_count_33_io_out ? io_r_68_b : _GEN_3517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3519 = 7'h45 == r_count_33_io_out ? io_r_69_b : _GEN_3518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3520 = 7'h46 == r_count_33_io_out ? io_r_70_b : _GEN_3519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3521 = 7'h47 == r_count_33_io_out ? io_r_71_b : _GEN_3520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3522 = 7'h48 == r_count_33_io_out ? io_r_72_b : _GEN_3521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3523 = 7'h49 == r_count_33_io_out ? io_r_73_b : _GEN_3522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3524 = 7'h4a == r_count_33_io_out ? io_r_74_b : _GEN_3523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3525 = 7'h4b == r_count_33_io_out ? io_r_75_b : _GEN_3524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3526 = 7'h4c == r_count_33_io_out ? io_r_76_b : _GEN_3525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3527 = 7'h4d == r_count_33_io_out ? io_r_77_b : _GEN_3526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3528 = 7'h4e == r_count_33_io_out ? io_r_78_b : _GEN_3527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3529 = 7'h4f == r_count_33_io_out ? io_r_79_b : _GEN_3528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3530 = 7'h50 == r_count_33_io_out ? io_r_80_b : _GEN_3529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3531 = 7'h51 == r_count_33_io_out ? io_r_81_b : _GEN_3530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3532 = 7'h52 == r_count_33_io_out ? io_r_82_b : _GEN_3531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3533 = 7'h53 == r_count_33_io_out ? io_r_83_b : _GEN_3532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3534 = 7'h54 == r_count_33_io_out ? io_r_84_b : _GEN_3533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3535 = 7'h55 == r_count_33_io_out ? io_r_85_b : _GEN_3534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3536 = 7'h56 == r_count_33_io_out ? io_r_86_b : _GEN_3535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3537 = 7'h57 == r_count_33_io_out ? io_r_87_b : _GEN_3536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3538 = 7'h58 == r_count_33_io_out ? io_r_88_b : _GEN_3537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3539 = 7'h59 == r_count_33_io_out ? io_r_89_b : _GEN_3538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3540 = 7'h5a == r_count_33_io_out ? io_r_90_b : _GEN_3539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3541 = 7'h5b == r_count_33_io_out ? io_r_91_b : _GEN_3540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3542 = 7'h5c == r_count_33_io_out ? io_r_92_b : _GEN_3541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3543 = 7'h5d == r_count_33_io_out ? io_r_93_b : _GEN_3542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3544 = 7'h5e == r_count_33_io_out ? io_r_94_b : _GEN_3543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3545 = 7'h5f == r_count_33_io_out ? io_r_95_b : _GEN_3544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3546 = 7'h60 == r_count_33_io_out ? io_r_96_b : _GEN_3545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3547 = 7'h61 == r_count_33_io_out ? io_r_97_b : _GEN_3546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3548 = 7'h62 == r_count_33_io_out ? io_r_98_b : _GEN_3547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3551 = 7'h1 == r_count_34_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3552 = 7'h2 == r_count_34_io_out ? io_r_2_b : _GEN_3551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3553 = 7'h3 == r_count_34_io_out ? io_r_3_b : _GEN_3552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3554 = 7'h4 == r_count_34_io_out ? io_r_4_b : _GEN_3553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3555 = 7'h5 == r_count_34_io_out ? io_r_5_b : _GEN_3554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3556 = 7'h6 == r_count_34_io_out ? io_r_6_b : _GEN_3555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3557 = 7'h7 == r_count_34_io_out ? io_r_7_b : _GEN_3556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3558 = 7'h8 == r_count_34_io_out ? io_r_8_b : _GEN_3557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3559 = 7'h9 == r_count_34_io_out ? io_r_9_b : _GEN_3558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3560 = 7'ha == r_count_34_io_out ? io_r_10_b : _GEN_3559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3561 = 7'hb == r_count_34_io_out ? io_r_11_b : _GEN_3560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3562 = 7'hc == r_count_34_io_out ? io_r_12_b : _GEN_3561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3563 = 7'hd == r_count_34_io_out ? io_r_13_b : _GEN_3562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3564 = 7'he == r_count_34_io_out ? io_r_14_b : _GEN_3563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3565 = 7'hf == r_count_34_io_out ? io_r_15_b : _GEN_3564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3566 = 7'h10 == r_count_34_io_out ? io_r_16_b : _GEN_3565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3567 = 7'h11 == r_count_34_io_out ? io_r_17_b : _GEN_3566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3568 = 7'h12 == r_count_34_io_out ? io_r_18_b : _GEN_3567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3569 = 7'h13 == r_count_34_io_out ? io_r_19_b : _GEN_3568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3570 = 7'h14 == r_count_34_io_out ? io_r_20_b : _GEN_3569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3571 = 7'h15 == r_count_34_io_out ? io_r_21_b : _GEN_3570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3572 = 7'h16 == r_count_34_io_out ? io_r_22_b : _GEN_3571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3573 = 7'h17 == r_count_34_io_out ? io_r_23_b : _GEN_3572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3574 = 7'h18 == r_count_34_io_out ? io_r_24_b : _GEN_3573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3575 = 7'h19 == r_count_34_io_out ? io_r_25_b : _GEN_3574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3576 = 7'h1a == r_count_34_io_out ? io_r_26_b : _GEN_3575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3577 = 7'h1b == r_count_34_io_out ? io_r_27_b : _GEN_3576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3578 = 7'h1c == r_count_34_io_out ? io_r_28_b : _GEN_3577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3579 = 7'h1d == r_count_34_io_out ? io_r_29_b : _GEN_3578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3580 = 7'h1e == r_count_34_io_out ? io_r_30_b : _GEN_3579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3581 = 7'h1f == r_count_34_io_out ? io_r_31_b : _GEN_3580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3582 = 7'h20 == r_count_34_io_out ? io_r_32_b : _GEN_3581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3583 = 7'h21 == r_count_34_io_out ? io_r_33_b : _GEN_3582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3584 = 7'h22 == r_count_34_io_out ? io_r_34_b : _GEN_3583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3585 = 7'h23 == r_count_34_io_out ? io_r_35_b : _GEN_3584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3586 = 7'h24 == r_count_34_io_out ? io_r_36_b : _GEN_3585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3587 = 7'h25 == r_count_34_io_out ? io_r_37_b : _GEN_3586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3588 = 7'h26 == r_count_34_io_out ? io_r_38_b : _GEN_3587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3589 = 7'h27 == r_count_34_io_out ? io_r_39_b : _GEN_3588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3590 = 7'h28 == r_count_34_io_out ? io_r_40_b : _GEN_3589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3591 = 7'h29 == r_count_34_io_out ? io_r_41_b : _GEN_3590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3592 = 7'h2a == r_count_34_io_out ? io_r_42_b : _GEN_3591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3593 = 7'h2b == r_count_34_io_out ? io_r_43_b : _GEN_3592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3594 = 7'h2c == r_count_34_io_out ? io_r_44_b : _GEN_3593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3595 = 7'h2d == r_count_34_io_out ? io_r_45_b : _GEN_3594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3596 = 7'h2e == r_count_34_io_out ? io_r_46_b : _GEN_3595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3597 = 7'h2f == r_count_34_io_out ? io_r_47_b : _GEN_3596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3598 = 7'h30 == r_count_34_io_out ? io_r_48_b : _GEN_3597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3599 = 7'h31 == r_count_34_io_out ? io_r_49_b : _GEN_3598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3600 = 7'h32 == r_count_34_io_out ? io_r_50_b : _GEN_3599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3601 = 7'h33 == r_count_34_io_out ? io_r_51_b : _GEN_3600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3602 = 7'h34 == r_count_34_io_out ? io_r_52_b : _GEN_3601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3603 = 7'h35 == r_count_34_io_out ? io_r_53_b : _GEN_3602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3604 = 7'h36 == r_count_34_io_out ? io_r_54_b : _GEN_3603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3605 = 7'h37 == r_count_34_io_out ? io_r_55_b : _GEN_3604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3606 = 7'h38 == r_count_34_io_out ? io_r_56_b : _GEN_3605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3607 = 7'h39 == r_count_34_io_out ? io_r_57_b : _GEN_3606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3608 = 7'h3a == r_count_34_io_out ? io_r_58_b : _GEN_3607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3609 = 7'h3b == r_count_34_io_out ? io_r_59_b : _GEN_3608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3610 = 7'h3c == r_count_34_io_out ? io_r_60_b : _GEN_3609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3611 = 7'h3d == r_count_34_io_out ? io_r_61_b : _GEN_3610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3612 = 7'h3e == r_count_34_io_out ? io_r_62_b : _GEN_3611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3613 = 7'h3f == r_count_34_io_out ? io_r_63_b : _GEN_3612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3614 = 7'h40 == r_count_34_io_out ? io_r_64_b : _GEN_3613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3615 = 7'h41 == r_count_34_io_out ? io_r_65_b : _GEN_3614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3616 = 7'h42 == r_count_34_io_out ? io_r_66_b : _GEN_3615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3617 = 7'h43 == r_count_34_io_out ? io_r_67_b : _GEN_3616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3618 = 7'h44 == r_count_34_io_out ? io_r_68_b : _GEN_3617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3619 = 7'h45 == r_count_34_io_out ? io_r_69_b : _GEN_3618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3620 = 7'h46 == r_count_34_io_out ? io_r_70_b : _GEN_3619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3621 = 7'h47 == r_count_34_io_out ? io_r_71_b : _GEN_3620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3622 = 7'h48 == r_count_34_io_out ? io_r_72_b : _GEN_3621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3623 = 7'h49 == r_count_34_io_out ? io_r_73_b : _GEN_3622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3624 = 7'h4a == r_count_34_io_out ? io_r_74_b : _GEN_3623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3625 = 7'h4b == r_count_34_io_out ? io_r_75_b : _GEN_3624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3626 = 7'h4c == r_count_34_io_out ? io_r_76_b : _GEN_3625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3627 = 7'h4d == r_count_34_io_out ? io_r_77_b : _GEN_3626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3628 = 7'h4e == r_count_34_io_out ? io_r_78_b : _GEN_3627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3629 = 7'h4f == r_count_34_io_out ? io_r_79_b : _GEN_3628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3630 = 7'h50 == r_count_34_io_out ? io_r_80_b : _GEN_3629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3631 = 7'h51 == r_count_34_io_out ? io_r_81_b : _GEN_3630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3632 = 7'h52 == r_count_34_io_out ? io_r_82_b : _GEN_3631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3633 = 7'h53 == r_count_34_io_out ? io_r_83_b : _GEN_3632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3634 = 7'h54 == r_count_34_io_out ? io_r_84_b : _GEN_3633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3635 = 7'h55 == r_count_34_io_out ? io_r_85_b : _GEN_3634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3636 = 7'h56 == r_count_34_io_out ? io_r_86_b : _GEN_3635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3637 = 7'h57 == r_count_34_io_out ? io_r_87_b : _GEN_3636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3638 = 7'h58 == r_count_34_io_out ? io_r_88_b : _GEN_3637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3639 = 7'h59 == r_count_34_io_out ? io_r_89_b : _GEN_3638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3640 = 7'h5a == r_count_34_io_out ? io_r_90_b : _GEN_3639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3641 = 7'h5b == r_count_34_io_out ? io_r_91_b : _GEN_3640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3642 = 7'h5c == r_count_34_io_out ? io_r_92_b : _GEN_3641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3643 = 7'h5d == r_count_34_io_out ? io_r_93_b : _GEN_3642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3644 = 7'h5e == r_count_34_io_out ? io_r_94_b : _GEN_3643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3645 = 7'h5f == r_count_34_io_out ? io_r_95_b : _GEN_3644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3646 = 7'h60 == r_count_34_io_out ? io_r_96_b : _GEN_3645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3647 = 7'h61 == r_count_34_io_out ? io_r_97_b : _GEN_3646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3648 = 7'h62 == r_count_34_io_out ? io_r_98_b : _GEN_3647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3651 = 7'h1 == r_count_35_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3652 = 7'h2 == r_count_35_io_out ? io_r_2_b : _GEN_3651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3653 = 7'h3 == r_count_35_io_out ? io_r_3_b : _GEN_3652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3654 = 7'h4 == r_count_35_io_out ? io_r_4_b : _GEN_3653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3655 = 7'h5 == r_count_35_io_out ? io_r_5_b : _GEN_3654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3656 = 7'h6 == r_count_35_io_out ? io_r_6_b : _GEN_3655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3657 = 7'h7 == r_count_35_io_out ? io_r_7_b : _GEN_3656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3658 = 7'h8 == r_count_35_io_out ? io_r_8_b : _GEN_3657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3659 = 7'h9 == r_count_35_io_out ? io_r_9_b : _GEN_3658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3660 = 7'ha == r_count_35_io_out ? io_r_10_b : _GEN_3659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3661 = 7'hb == r_count_35_io_out ? io_r_11_b : _GEN_3660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3662 = 7'hc == r_count_35_io_out ? io_r_12_b : _GEN_3661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3663 = 7'hd == r_count_35_io_out ? io_r_13_b : _GEN_3662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3664 = 7'he == r_count_35_io_out ? io_r_14_b : _GEN_3663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3665 = 7'hf == r_count_35_io_out ? io_r_15_b : _GEN_3664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3666 = 7'h10 == r_count_35_io_out ? io_r_16_b : _GEN_3665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3667 = 7'h11 == r_count_35_io_out ? io_r_17_b : _GEN_3666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3668 = 7'h12 == r_count_35_io_out ? io_r_18_b : _GEN_3667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3669 = 7'h13 == r_count_35_io_out ? io_r_19_b : _GEN_3668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3670 = 7'h14 == r_count_35_io_out ? io_r_20_b : _GEN_3669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3671 = 7'h15 == r_count_35_io_out ? io_r_21_b : _GEN_3670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3672 = 7'h16 == r_count_35_io_out ? io_r_22_b : _GEN_3671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3673 = 7'h17 == r_count_35_io_out ? io_r_23_b : _GEN_3672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3674 = 7'h18 == r_count_35_io_out ? io_r_24_b : _GEN_3673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3675 = 7'h19 == r_count_35_io_out ? io_r_25_b : _GEN_3674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3676 = 7'h1a == r_count_35_io_out ? io_r_26_b : _GEN_3675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3677 = 7'h1b == r_count_35_io_out ? io_r_27_b : _GEN_3676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3678 = 7'h1c == r_count_35_io_out ? io_r_28_b : _GEN_3677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3679 = 7'h1d == r_count_35_io_out ? io_r_29_b : _GEN_3678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3680 = 7'h1e == r_count_35_io_out ? io_r_30_b : _GEN_3679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3681 = 7'h1f == r_count_35_io_out ? io_r_31_b : _GEN_3680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3682 = 7'h20 == r_count_35_io_out ? io_r_32_b : _GEN_3681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3683 = 7'h21 == r_count_35_io_out ? io_r_33_b : _GEN_3682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3684 = 7'h22 == r_count_35_io_out ? io_r_34_b : _GEN_3683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3685 = 7'h23 == r_count_35_io_out ? io_r_35_b : _GEN_3684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3686 = 7'h24 == r_count_35_io_out ? io_r_36_b : _GEN_3685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3687 = 7'h25 == r_count_35_io_out ? io_r_37_b : _GEN_3686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3688 = 7'h26 == r_count_35_io_out ? io_r_38_b : _GEN_3687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3689 = 7'h27 == r_count_35_io_out ? io_r_39_b : _GEN_3688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3690 = 7'h28 == r_count_35_io_out ? io_r_40_b : _GEN_3689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3691 = 7'h29 == r_count_35_io_out ? io_r_41_b : _GEN_3690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3692 = 7'h2a == r_count_35_io_out ? io_r_42_b : _GEN_3691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3693 = 7'h2b == r_count_35_io_out ? io_r_43_b : _GEN_3692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3694 = 7'h2c == r_count_35_io_out ? io_r_44_b : _GEN_3693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3695 = 7'h2d == r_count_35_io_out ? io_r_45_b : _GEN_3694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3696 = 7'h2e == r_count_35_io_out ? io_r_46_b : _GEN_3695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3697 = 7'h2f == r_count_35_io_out ? io_r_47_b : _GEN_3696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3698 = 7'h30 == r_count_35_io_out ? io_r_48_b : _GEN_3697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3699 = 7'h31 == r_count_35_io_out ? io_r_49_b : _GEN_3698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3700 = 7'h32 == r_count_35_io_out ? io_r_50_b : _GEN_3699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3701 = 7'h33 == r_count_35_io_out ? io_r_51_b : _GEN_3700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3702 = 7'h34 == r_count_35_io_out ? io_r_52_b : _GEN_3701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3703 = 7'h35 == r_count_35_io_out ? io_r_53_b : _GEN_3702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3704 = 7'h36 == r_count_35_io_out ? io_r_54_b : _GEN_3703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3705 = 7'h37 == r_count_35_io_out ? io_r_55_b : _GEN_3704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3706 = 7'h38 == r_count_35_io_out ? io_r_56_b : _GEN_3705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3707 = 7'h39 == r_count_35_io_out ? io_r_57_b : _GEN_3706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3708 = 7'h3a == r_count_35_io_out ? io_r_58_b : _GEN_3707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3709 = 7'h3b == r_count_35_io_out ? io_r_59_b : _GEN_3708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3710 = 7'h3c == r_count_35_io_out ? io_r_60_b : _GEN_3709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3711 = 7'h3d == r_count_35_io_out ? io_r_61_b : _GEN_3710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3712 = 7'h3e == r_count_35_io_out ? io_r_62_b : _GEN_3711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3713 = 7'h3f == r_count_35_io_out ? io_r_63_b : _GEN_3712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3714 = 7'h40 == r_count_35_io_out ? io_r_64_b : _GEN_3713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3715 = 7'h41 == r_count_35_io_out ? io_r_65_b : _GEN_3714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3716 = 7'h42 == r_count_35_io_out ? io_r_66_b : _GEN_3715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3717 = 7'h43 == r_count_35_io_out ? io_r_67_b : _GEN_3716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3718 = 7'h44 == r_count_35_io_out ? io_r_68_b : _GEN_3717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3719 = 7'h45 == r_count_35_io_out ? io_r_69_b : _GEN_3718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3720 = 7'h46 == r_count_35_io_out ? io_r_70_b : _GEN_3719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3721 = 7'h47 == r_count_35_io_out ? io_r_71_b : _GEN_3720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3722 = 7'h48 == r_count_35_io_out ? io_r_72_b : _GEN_3721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3723 = 7'h49 == r_count_35_io_out ? io_r_73_b : _GEN_3722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3724 = 7'h4a == r_count_35_io_out ? io_r_74_b : _GEN_3723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3725 = 7'h4b == r_count_35_io_out ? io_r_75_b : _GEN_3724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3726 = 7'h4c == r_count_35_io_out ? io_r_76_b : _GEN_3725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3727 = 7'h4d == r_count_35_io_out ? io_r_77_b : _GEN_3726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3728 = 7'h4e == r_count_35_io_out ? io_r_78_b : _GEN_3727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3729 = 7'h4f == r_count_35_io_out ? io_r_79_b : _GEN_3728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3730 = 7'h50 == r_count_35_io_out ? io_r_80_b : _GEN_3729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3731 = 7'h51 == r_count_35_io_out ? io_r_81_b : _GEN_3730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3732 = 7'h52 == r_count_35_io_out ? io_r_82_b : _GEN_3731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3733 = 7'h53 == r_count_35_io_out ? io_r_83_b : _GEN_3732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3734 = 7'h54 == r_count_35_io_out ? io_r_84_b : _GEN_3733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3735 = 7'h55 == r_count_35_io_out ? io_r_85_b : _GEN_3734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3736 = 7'h56 == r_count_35_io_out ? io_r_86_b : _GEN_3735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3737 = 7'h57 == r_count_35_io_out ? io_r_87_b : _GEN_3736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3738 = 7'h58 == r_count_35_io_out ? io_r_88_b : _GEN_3737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3739 = 7'h59 == r_count_35_io_out ? io_r_89_b : _GEN_3738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3740 = 7'h5a == r_count_35_io_out ? io_r_90_b : _GEN_3739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3741 = 7'h5b == r_count_35_io_out ? io_r_91_b : _GEN_3740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3742 = 7'h5c == r_count_35_io_out ? io_r_92_b : _GEN_3741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3743 = 7'h5d == r_count_35_io_out ? io_r_93_b : _GEN_3742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3744 = 7'h5e == r_count_35_io_out ? io_r_94_b : _GEN_3743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3745 = 7'h5f == r_count_35_io_out ? io_r_95_b : _GEN_3744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3746 = 7'h60 == r_count_35_io_out ? io_r_96_b : _GEN_3745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3747 = 7'h61 == r_count_35_io_out ? io_r_97_b : _GEN_3746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3748 = 7'h62 == r_count_35_io_out ? io_r_98_b : _GEN_3747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3751 = 7'h1 == r_count_36_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3752 = 7'h2 == r_count_36_io_out ? io_r_2_b : _GEN_3751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3753 = 7'h3 == r_count_36_io_out ? io_r_3_b : _GEN_3752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3754 = 7'h4 == r_count_36_io_out ? io_r_4_b : _GEN_3753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3755 = 7'h5 == r_count_36_io_out ? io_r_5_b : _GEN_3754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3756 = 7'h6 == r_count_36_io_out ? io_r_6_b : _GEN_3755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3757 = 7'h7 == r_count_36_io_out ? io_r_7_b : _GEN_3756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3758 = 7'h8 == r_count_36_io_out ? io_r_8_b : _GEN_3757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3759 = 7'h9 == r_count_36_io_out ? io_r_9_b : _GEN_3758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3760 = 7'ha == r_count_36_io_out ? io_r_10_b : _GEN_3759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3761 = 7'hb == r_count_36_io_out ? io_r_11_b : _GEN_3760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3762 = 7'hc == r_count_36_io_out ? io_r_12_b : _GEN_3761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3763 = 7'hd == r_count_36_io_out ? io_r_13_b : _GEN_3762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3764 = 7'he == r_count_36_io_out ? io_r_14_b : _GEN_3763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3765 = 7'hf == r_count_36_io_out ? io_r_15_b : _GEN_3764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3766 = 7'h10 == r_count_36_io_out ? io_r_16_b : _GEN_3765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3767 = 7'h11 == r_count_36_io_out ? io_r_17_b : _GEN_3766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3768 = 7'h12 == r_count_36_io_out ? io_r_18_b : _GEN_3767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3769 = 7'h13 == r_count_36_io_out ? io_r_19_b : _GEN_3768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3770 = 7'h14 == r_count_36_io_out ? io_r_20_b : _GEN_3769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3771 = 7'h15 == r_count_36_io_out ? io_r_21_b : _GEN_3770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3772 = 7'h16 == r_count_36_io_out ? io_r_22_b : _GEN_3771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3773 = 7'h17 == r_count_36_io_out ? io_r_23_b : _GEN_3772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3774 = 7'h18 == r_count_36_io_out ? io_r_24_b : _GEN_3773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3775 = 7'h19 == r_count_36_io_out ? io_r_25_b : _GEN_3774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3776 = 7'h1a == r_count_36_io_out ? io_r_26_b : _GEN_3775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3777 = 7'h1b == r_count_36_io_out ? io_r_27_b : _GEN_3776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3778 = 7'h1c == r_count_36_io_out ? io_r_28_b : _GEN_3777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3779 = 7'h1d == r_count_36_io_out ? io_r_29_b : _GEN_3778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3780 = 7'h1e == r_count_36_io_out ? io_r_30_b : _GEN_3779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3781 = 7'h1f == r_count_36_io_out ? io_r_31_b : _GEN_3780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3782 = 7'h20 == r_count_36_io_out ? io_r_32_b : _GEN_3781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3783 = 7'h21 == r_count_36_io_out ? io_r_33_b : _GEN_3782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3784 = 7'h22 == r_count_36_io_out ? io_r_34_b : _GEN_3783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3785 = 7'h23 == r_count_36_io_out ? io_r_35_b : _GEN_3784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3786 = 7'h24 == r_count_36_io_out ? io_r_36_b : _GEN_3785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3787 = 7'h25 == r_count_36_io_out ? io_r_37_b : _GEN_3786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3788 = 7'h26 == r_count_36_io_out ? io_r_38_b : _GEN_3787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3789 = 7'h27 == r_count_36_io_out ? io_r_39_b : _GEN_3788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3790 = 7'h28 == r_count_36_io_out ? io_r_40_b : _GEN_3789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3791 = 7'h29 == r_count_36_io_out ? io_r_41_b : _GEN_3790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3792 = 7'h2a == r_count_36_io_out ? io_r_42_b : _GEN_3791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3793 = 7'h2b == r_count_36_io_out ? io_r_43_b : _GEN_3792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3794 = 7'h2c == r_count_36_io_out ? io_r_44_b : _GEN_3793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3795 = 7'h2d == r_count_36_io_out ? io_r_45_b : _GEN_3794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3796 = 7'h2e == r_count_36_io_out ? io_r_46_b : _GEN_3795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3797 = 7'h2f == r_count_36_io_out ? io_r_47_b : _GEN_3796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3798 = 7'h30 == r_count_36_io_out ? io_r_48_b : _GEN_3797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3799 = 7'h31 == r_count_36_io_out ? io_r_49_b : _GEN_3798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3800 = 7'h32 == r_count_36_io_out ? io_r_50_b : _GEN_3799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3801 = 7'h33 == r_count_36_io_out ? io_r_51_b : _GEN_3800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3802 = 7'h34 == r_count_36_io_out ? io_r_52_b : _GEN_3801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3803 = 7'h35 == r_count_36_io_out ? io_r_53_b : _GEN_3802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3804 = 7'h36 == r_count_36_io_out ? io_r_54_b : _GEN_3803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3805 = 7'h37 == r_count_36_io_out ? io_r_55_b : _GEN_3804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3806 = 7'h38 == r_count_36_io_out ? io_r_56_b : _GEN_3805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3807 = 7'h39 == r_count_36_io_out ? io_r_57_b : _GEN_3806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3808 = 7'h3a == r_count_36_io_out ? io_r_58_b : _GEN_3807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3809 = 7'h3b == r_count_36_io_out ? io_r_59_b : _GEN_3808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3810 = 7'h3c == r_count_36_io_out ? io_r_60_b : _GEN_3809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3811 = 7'h3d == r_count_36_io_out ? io_r_61_b : _GEN_3810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3812 = 7'h3e == r_count_36_io_out ? io_r_62_b : _GEN_3811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3813 = 7'h3f == r_count_36_io_out ? io_r_63_b : _GEN_3812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3814 = 7'h40 == r_count_36_io_out ? io_r_64_b : _GEN_3813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3815 = 7'h41 == r_count_36_io_out ? io_r_65_b : _GEN_3814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3816 = 7'h42 == r_count_36_io_out ? io_r_66_b : _GEN_3815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3817 = 7'h43 == r_count_36_io_out ? io_r_67_b : _GEN_3816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3818 = 7'h44 == r_count_36_io_out ? io_r_68_b : _GEN_3817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3819 = 7'h45 == r_count_36_io_out ? io_r_69_b : _GEN_3818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3820 = 7'h46 == r_count_36_io_out ? io_r_70_b : _GEN_3819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3821 = 7'h47 == r_count_36_io_out ? io_r_71_b : _GEN_3820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3822 = 7'h48 == r_count_36_io_out ? io_r_72_b : _GEN_3821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3823 = 7'h49 == r_count_36_io_out ? io_r_73_b : _GEN_3822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3824 = 7'h4a == r_count_36_io_out ? io_r_74_b : _GEN_3823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3825 = 7'h4b == r_count_36_io_out ? io_r_75_b : _GEN_3824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3826 = 7'h4c == r_count_36_io_out ? io_r_76_b : _GEN_3825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3827 = 7'h4d == r_count_36_io_out ? io_r_77_b : _GEN_3826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3828 = 7'h4e == r_count_36_io_out ? io_r_78_b : _GEN_3827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3829 = 7'h4f == r_count_36_io_out ? io_r_79_b : _GEN_3828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3830 = 7'h50 == r_count_36_io_out ? io_r_80_b : _GEN_3829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3831 = 7'h51 == r_count_36_io_out ? io_r_81_b : _GEN_3830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3832 = 7'h52 == r_count_36_io_out ? io_r_82_b : _GEN_3831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3833 = 7'h53 == r_count_36_io_out ? io_r_83_b : _GEN_3832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3834 = 7'h54 == r_count_36_io_out ? io_r_84_b : _GEN_3833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3835 = 7'h55 == r_count_36_io_out ? io_r_85_b : _GEN_3834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3836 = 7'h56 == r_count_36_io_out ? io_r_86_b : _GEN_3835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3837 = 7'h57 == r_count_36_io_out ? io_r_87_b : _GEN_3836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3838 = 7'h58 == r_count_36_io_out ? io_r_88_b : _GEN_3837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3839 = 7'h59 == r_count_36_io_out ? io_r_89_b : _GEN_3838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3840 = 7'h5a == r_count_36_io_out ? io_r_90_b : _GEN_3839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3841 = 7'h5b == r_count_36_io_out ? io_r_91_b : _GEN_3840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3842 = 7'h5c == r_count_36_io_out ? io_r_92_b : _GEN_3841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3843 = 7'h5d == r_count_36_io_out ? io_r_93_b : _GEN_3842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3844 = 7'h5e == r_count_36_io_out ? io_r_94_b : _GEN_3843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3845 = 7'h5f == r_count_36_io_out ? io_r_95_b : _GEN_3844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3846 = 7'h60 == r_count_36_io_out ? io_r_96_b : _GEN_3845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3847 = 7'h61 == r_count_36_io_out ? io_r_97_b : _GEN_3846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3848 = 7'h62 == r_count_36_io_out ? io_r_98_b : _GEN_3847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3851 = 7'h1 == r_count_37_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3852 = 7'h2 == r_count_37_io_out ? io_r_2_b : _GEN_3851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3853 = 7'h3 == r_count_37_io_out ? io_r_3_b : _GEN_3852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3854 = 7'h4 == r_count_37_io_out ? io_r_4_b : _GEN_3853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3855 = 7'h5 == r_count_37_io_out ? io_r_5_b : _GEN_3854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3856 = 7'h6 == r_count_37_io_out ? io_r_6_b : _GEN_3855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3857 = 7'h7 == r_count_37_io_out ? io_r_7_b : _GEN_3856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3858 = 7'h8 == r_count_37_io_out ? io_r_8_b : _GEN_3857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3859 = 7'h9 == r_count_37_io_out ? io_r_9_b : _GEN_3858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3860 = 7'ha == r_count_37_io_out ? io_r_10_b : _GEN_3859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3861 = 7'hb == r_count_37_io_out ? io_r_11_b : _GEN_3860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3862 = 7'hc == r_count_37_io_out ? io_r_12_b : _GEN_3861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3863 = 7'hd == r_count_37_io_out ? io_r_13_b : _GEN_3862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3864 = 7'he == r_count_37_io_out ? io_r_14_b : _GEN_3863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3865 = 7'hf == r_count_37_io_out ? io_r_15_b : _GEN_3864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3866 = 7'h10 == r_count_37_io_out ? io_r_16_b : _GEN_3865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3867 = 7'h11 == r_count_37_io_out ? io_r_17_b : _GEN_3866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3868 = 7'h12 == r_count_37_io_out ? io_r_18_b : _GEN_3867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3869 = 7'h13 == r_count_37_io_out ? io_r_19_b : _GEN_3868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3870 = 7'h14 == r_count_37_io_out ? io_r_20_b : _GEN_3869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3871 = 7'h15 == r_count_37_io_out ? io_r_21_b : _GEN_3870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3872 = 7'h16 == r_count_37_io_out ? io_r_22_b : _GEN_3871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3873 = 7'h17 == r_count_37_io_out ? io_r_23_b : _GEN_3872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3874 = 7'h18 == r_count_37_io_out ? io_r_24_b : _GEN_3873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3875 = 7'h19 == r_count_37_io_out ? io_r_25_b : _GEN_3874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3876 = 7'h1a == r_count_37_io_out ? io_r_26_b : _GEN_3875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3877 = 7'h1b == r_count_37_io_out ? io_r_27_b : _GEN_3876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3878 = 7'h1c == r_count_37_io_out ? io_r_28_b : _GEN_3877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3879 = 7'h1d == r_count_37_io_out ? io_r_29_b : _GEN_3878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3880 = 7'h1e == r_count_37_io_out ? io_r_30_b : _GEN_3879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3881 = 7'h1f == r_count_37_io_out ? io_r_31_b : _GEN_3880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3882 = 7'h20 == r_count_37_io_out ? io_r_32_b : _GEN_3881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3883 = 7'h21 == r_count_37_io_out ? io_r_33_b : _GEN_3882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3884 = 7'h22 == r_count_37_io_out ? io_r_34_b : _GEN_3883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3885 = 7'h23 == r_count_37_io_out ? io_r_35_b : _GEN_3884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3886 = 7'h24 == r_count_37_io_out ? io_r_36_b : _GEN_3885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3887 = 7'h25 == r_count_37_io_out ? io_r_37_b : _GEN_3886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3888 = 7'h26 == r_count_37_io_out ? io_r_38_b : _GEN_3887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3889 = 7'h27 == r_count_37_io_out ? io_r_39_b : _GEN_3888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3890 = 7'h28 == r_count_37_io_out ? io_r_40_b : _GEN_3889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3891 = 7'h29 == r_count_37_io_out ? io_r_41_b : _GEN_3890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3892 = 7'h2a == r_count_37_io_out ? io_r_42_b : _GEN_3891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3893 = 7'h2b == r_count_37_io_out ? io_r_43_b : _GEN_3892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3894 = 7'h2c == r_count_37_io_out ? io_r_44_b : _GEN_3893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3895 = 7'h2d == r_count_37_io_out ? io_r_45_b : _GEN_3894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3896 = 7'h2e == r_count_37_io_out ? io_r_46_b : _GEN_3895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3897 = 7'h2f == r_count_37_io_out ? io_r_47_b : _GEN_3896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3898 = 7'h30 == r_count_37_io_out ? io_r_48_b : _GEN_3897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3899 = 7'h31 == r_count_37_io_out ? io_r_49_b : _GEN_3898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3900 = 7'h32 == r_count_37_io_out ? io_r_50_b : _GEN_3899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3901 = 7'h33 == r_count_37_io_out ? io_r_51_b : _GEN_3900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3902 = 7'h34 == r_count_37_io_out ? io_r_52_b : _GEN_3901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3903 = 7'h35 == r_count_37_io_out ? io_r_53_b : _GEN_3902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3904 = 7'h36 == r_count_37_io_out ? io_r_54_b : _GEN_3903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3905 = 7'h37 == r_count_37_io_out ? io_r_55_b : _GEN_3904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3906 = 7'h38 == r_count_37_io_out ? io_r_56_b : _GEN_3905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3907 = 7'h39 == r_count_37_io_out ? io_r_57_b : _GEN_3906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3908 = 7'h3a == r_count_37_io_out ? io_r_58_b : _GEN_3907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3909 = 7'h3b == r_count_37_io_out ? io_r_59_b : _GEN_3908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3910 = 7'h3c == r_count_37_io_out ? io_r_60_b : _GEN_3909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3911 = 7'h3d == r_count_37_io_out ? io_r_61_b : _GEN_3910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3912 = 7'h3e == r_count_37_io_out ? io_r_62_b : _GEN_3911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3913 = 7'h3f == r_count_37_io_out ? io_r_63_b : _GEN_3912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3914 = 7'h40 == r_count_37_io_out ? io_r_64_b : _GEN_3913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3915 = 7'h41 == r_count_37_io_out ? io_r_65_b : _GEN_3914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3916 = 7'h42 == r_count_37_io_out ? io_r_66_b : _GEN_3915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3917 = 7'h43 == r_count_37_io_out ? io_r_67_b : _GEN_3916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3918 = 7'h44 == r_count_37_io_out ? io_r_68_b : _GEN_3917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3919 = 7'h45 == r_count_37_io_out ? io_r_69_b : _GEN_3918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3920 = 7'h46 == r_count_37_io_out ? io_r_70_b : _GEN_3919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3921 = 7'h47 == r_count_37_io_out ? io_r_71_b : _GEN_3920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3922 = 7'h48 == r_count_37_io_out ? io_r_72_b : _GEN_3921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3923 = 7'h49 == r_count_37_io_out ? io_r_73_b : _GEN_3922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3924 = 7'h4a == r_count_37_io_out ? io_r_74_b : _GEN_3923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3925 = 7'h4b == r_count_37_io_out ? io_r_75_b : _GEN_3924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3926 = 7'h4c == r_count_37_io_out ? io_r_76_b : _GEN_3925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3927 = 7'h4d == r_count_37_io_out ? io_r_77_b : _GEN_3926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3928 = 7'h4e == r_count_37_io_out ? io_r_78_b : _GEN_3927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3929 = 7'h4f == r_count_37_io_out ? io_r_79_b : _GEN_3928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3930 = 7'h50 == r_count_37_io_out ? io_r_80_b : _GEN_3929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3931 = 7'h51 == r_count_37_io_out ? io_r_81_b : _GEN_3930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3932 = 7'h52 == r_count_37_io_out ? io_r_82_b : _GEN_3931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3933 = 7'h53 == r_count_37_io_out ? io_r_83_b : _GEN_3932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3934 = 7'h54 == r_count_37_io_out ? io_r_84_b : _GEN_3933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3935 = 7'h55 == r_count_37_io_out ? io_r_85_b : _GEN_3934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3936 = 7'h56 == r_count_37_io_out ? io_r_86_b : _GEN_3935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3937 = 7'h57 == r_count_37_io_out ? io_r_87_b : _GEN_3936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3938 = 7'h58 == r_count_37_io_out ? io_r_88_b : _GEN_3937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3939 = 7'h59 == r_count_37_io_out ? io_r_89_b : _GEN_3938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3940 = 7'h5a == r_count_37_io_out ? io_r_90_b : _GEN_3939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3941 = 7'h5b == r_count_37_io_out ? io_r_91_b : _GEN_3940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3942 = 7'h5c == r_count_37_io_out ? io_r_92_b : _GEN_3941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3943 = 7'h5d == r_count_37_io_out ? io_r_93_b : _GEN_3942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3944 = 7'h5e == r_count_37_io_out ? io_r_94_b : _GEN_3943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3945 = 7'h5f == r_count_37_io_out ? io_r_95_b : _GEN_3944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3946 = 7'h60 == r_count_37_io_out ? io_r_96_b : _GEN_3945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3947 = 7'h61 == r_count_37_io_out ? io_r_97_b : _GEN_3946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3948 = 7'h62 == r_count_37_io_out ? io_r_98_b : _GEN_3947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3951 = 7'h1 == r_count_38_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3952 = 7'h2 == r_count_38_io_out ? io_r_2_b : _GEN_3951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3953 = 7'h3 == r_count_38_io_out ? io_r_3_b : _GEN_3952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3954 = 7'h4 == r_count_38_io_out ? io_r_4_b : _GEN_3953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3955 = 7'h5 == r_count_38_io_out ? io_r_5_b : _GEN_3954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3956 = 7'h6 == r_count_38_io_out ? io_r_6_b : _GEN_3955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3957 = 7'h7 == r_count_38_io_out ? io_r_7_b : _GEN_3956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3958 = 7'h8 == r_count_38_io_out ? io_r_8_b : _GEN_3957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3959 = 7'h9 == r_count_38_io_out ? io_r_9_b : _GEN_3958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3960 = 7'ha == r_count_38_io_out ? io_r_10_b : _GEN_3959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3961 = 7'hb == r_count_38_io_out ? io_r_11_b : _GEN_3960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3962 = 7'hc == r_count_38_io_out ? io_r_12_b : _GEN_3961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3963 = 7'hd == r_count_38_io_out ? io_r_13_b : _GEN_3962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3964 = 7'he == r_count_38_io_out ? io_r_14_b : _GEN_3963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3965 = 7'hf == r_count_38_io_out ? io_r_15_b : _GEN_3964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3966 = 7'h10 == r_count_38_io_out ? io_r_16_b : _GEN_3965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3967 = 7'h11 == r_count_38_io_out ? io_r_17_b : _GEN_3966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3968 = 7'h12 == r_count_38_io_out ? io_r_18_b : _GEN_3967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3969 = 7'h13 == r_count_38_io_out ? io_r_19_b : _GEN_3968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3970 = 7'h14 == r_count_38_io_out ? io_r_20_b : _GEN_3969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3971 = 7'h15 == r_count_38_io_out ? io_r_21_b : _GEN_3970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3972 = 7'h16 == r_count_38_io_out ? io_r_22_b : _GEN_3971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3973 = 7'h17 == r_count_38_io_out ? io_r_23_b : _GEN_3972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3974 = 7'h18 == r_count_38_io_out ? io_r_24_b : _GEN_3973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3975 = 7'h19 == r_count_38_io_out ? io_r_25_b : _GEN_3974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3976 = 7'h1a == r_count_38_io_out ? io_r_26_b : _GEN_3975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3977 = 7'h1b == r_count_38_io_out ? io_r_27_b : _GEN_3976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3978 = 7'h1c == r_count_38_io_out ? io_r_28_b : _GEN_3977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3979 = 7'h1d == r_count_38_io_out ? io_r_29_b : _GEN_3978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3980 = 7'h1e == r_count_38_io_out ? io_r_30_b : _GEN_3979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3981 = 7'h1f == r_count_38_io_out ? io_r_31_b : _GEN_3980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3982 = 7'h20 == r_count_38_io_out ? io_r_32_b : _GEN_3981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3983 = 7'h21 == r_count_38_io_out ? io_r_33_b : _GEN_3982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3984 = 7'h22 == r_count_38_io_out ? io_r_34_b : _GEN_3983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3985 = 7'h23 == r_count_38_io_out ? io_r_35_b : _GEN_3984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3986 = 7'h24 == r_count_38_io_out ? io_r_36_b : _GEN_3985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3987 = 7'h25 == r_count_38_io_out ? io_r_37_b : _GEN_3986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3988 = 7'h26 == r_count_38_io_out ? io_r_38_b : _GEN_3987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3989 = 7'h27 == r_count_38_io_out ? io_r_39_b : _GEN_3988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3990 = 7'h28 == r_count_38_io_out ? io_r_40_b : _GEN_3989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3991 = 7'h29 == r_count_38_io_out ? io_r_41_b : _GEN_3990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3992 = 7'h2a == r_count_38_io_out ? io_r_42_b : _GEN_3991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3993 = 7'h2b == r_count_38_io_out ? io_r_43_b : _GEN_3992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3994 = 7'h2c == r_count_38_io_out ? io_r_44_b : _GEN_3993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3995 = 7'h2d == r_count_38_io_out ? io_r_45_b : _GEN_3994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3996 = 7'h2e == r_count_38_io_out ? io_r_46_b : _GEN_3995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3997 = 7'h2f == r_count_38_io_out ? io_r_47_b : _GEN_3996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3998 = 7'h30 == r_count_38_io_out ? io_r_48_b : _GEN_3997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_3999 = 7'h31 == r_count_38_io_out ? io_r_49_b : _GEN_3998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4000 = 7'h32 == r_count_38_io_out ? io_r_50_b : _GEN_3999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4001 = 7'h33 == r_count_38_io_out ? io_r_51_b : _GEN_4000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4002 = 7'h34 == r_count_38_io_out ? io_r_52_b : _GEN_4001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4003 = 7'h35 == r_count_38_io_out ? io_r_53_b : _GEN_4002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4004 = 7'h36 == r_count_38_io_out ? io_r_54_b : _GEN_4003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4005 = 7'h37 == r_count_38_io_out ? io_r_55_b : _GEN_4004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4006 = 7'h38 == r_count_38_io_out ? io_r_56_b : _GEN_4005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4007 = 7'h39 == r_count_38_io_out ? io_r_57_b : _GEN_4006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4008 = 7'h3a == r_count_38_io_out ? io_r_58_b : _GEN_4007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4009 = 7'h3b == r_count_38_io_out ? io_r_59_b : _GEN_4008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4010 = 7'h3c == r_count_38_io_out ? io_r_60_b : _GEN_4009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4011 = 7'h3d == r_count_38_io_out ? io_r_61_b : _GEN_4010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4012 = 7'h3e == r_count_38_io_out ? io_r_62_b : _GEN_4011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4013 = 7'h3f == r_count_38_io_out ? io_r_63_b : _GEN_4012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4014 = 7'h40 == r_count_38_io_out ? io_r_64_b : _GEN_4013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4015 = 7'h41 == r_count_38_io_out ? io_r_65_b : _GEN_4014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4016 = 7'h42 == r_count_38_io_out ? io_r_66_b : _GEN_4015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4017 = 7'h43 == r_count_38_io_out ? io_r_67_b : _GEN_4016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4018 = 7'h44 == r_count_38_io_out ? io_r_68_b : _GEN_4017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4019 = 7'h45 == r_count_38_io_out ? io_r_69_b : _GEN_4018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4020 = 7'h46 == r_count_38_io_out ? io_r_70_b : _GEN_4019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4021 = 7'h47 == r_count_38_io_out ? io_r_71_b : _GEN_4020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4022 = 7'h48 == r_count_38_io_out ? io_r_72_b : _GEN_4021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4023 = 7'h49 == r_count_38_io_out ? io_r_73_b : _GEN_4022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4024 = 7'h4a == r_count_38_io_out ? io_r_74_b : _GEN_4023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4025 = 7'h4b == r_count_38_io_out ? io_r_75_b : _GEN_4024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4026 = 7'h4c == r_count_38_io_out ? io_r_76_b : _GEN_4025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4027 = 7'h4d == r_count_38_io_out ? io_r_77_b : _GEN_4026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4028 = 7'h4e == r_count_38_io_out ? io_r_78_b : _GEN_4027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4029 = 7'h4f == r_count_38_io_out ? io_r_79_b : _GEN_4028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4030 = 7'h50 == r_count_38_io_out ? io_r_80_b : _GEN_4029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4031 = 7'h51 == r_count_38_io_out ? io_r_81_b : _GEN_4030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4032 = 7'h52 == r_count_38_io_out ? io_r_82_b : _GEN_4031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4033 = 7'h53 == r_count_38_io_out ? io_r_83_b : _GEN_4032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4034 = 7'h54 == r_count_38_io_out ? io_r_84_b : _GEN_4033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4035 = 7'h55 == r_count_38_io_out ? io_r_85_b : _GEN_4034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4036 = 7'h56 == r_count_38_io_out ? io_r_86_b : _GEN_4035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4037 = 7'h57 == r_count_38_io_out ? io_r_87_b : _GEN_4036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4038 = 7'h58 == r_count_38_io_out ? io_r_88_b : _GEN_4037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4039 = 7'h59 == r_count_38_io_out ? io_r_89_b : _GEN_4038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4040 = 7'h5a == r_count_38_io_out ? io_r_90_b : _GEN_4039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4041 = 7'h5b == r_count_38_io_out ? io_r_91_b : _GEN_4040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4042 = 7'h5c == r_count_38_io_out ? io_r_92_b : _GEN_4041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4043 = 7'h5d == r_count_38_io_out ? io_r_93_b : _GEN_4042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4044 = 7'h5e == r_count_38_io_out ? io_r_94_b : _GEN_4043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4045 = 7'h5f == r_count_38_io_out ? io_r_95_b : _GEN_4044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4046 = 7'h60 == r_count_38_io_out ? io_r_96_b : _GEN_4045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4047 = 7'h61 == r_count_38_io_out ? io_r_97_b : _GEN_4046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4048 = 7'h62 == r_count_38_io_out ? io_r_98_b : _GEN_4047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4051 = 7'h1 == r_count_39_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4052 = 7'h2 == r_count_39_io_out ? io_r_2_b : _GEN_4051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4053 = 7'h3 == r_count_39_io_out ? io_r_3_b : _GEN_4052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4054 = 7'h4 == r_count_39_io_out ? io_r_4_b : _GEN_4053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4055 = 7'h5 == r_count_39_io_out ? io_r_5_b : _GEN_4054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4056 = 7'h6 == r_count_39_io_out ? io_r_6_b : _GEN_4055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4057 = 7'h7 == r_count_39_io_out ? io_r_7_b : _GEN_4056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4058 = 7'h8 == r_count_39_io_out ? io_r_8_b : _GEN_4057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4059 = 7'h9 == r_count_39_io_out ? io_r_9_b : _GEN_4058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4060 = 7'ha == r_count_39_io_out ? io_r_10_b : _GEN_4059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4061 = 7'hb == r_count_39_io_out ? io_r_11_b : _GEN_4060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4062 = 7'hc == r_count_39_io_out ? io_r_12_b : _GEN_4061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4063 = 7'hd == r_count_39_io_out ? io_r_13_b : _GEN_4062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4064 = 7'he == r_count_39_io_out ? io_r_14_b : _GEN_4063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4065 = 7'hf == r_count_39_io_out ? io_r_15_b : _GEN_4064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4066 = 7'h10 == r_count_39_io_out ? io_r_16_b : _GEN_4065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4067 = 7'h11 == r_count_39_io_out ? io_r_17_b : _GEN_4066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4068 = 7'h12 == r_count_39_io_out ? io_r_18_b : _GEN_4067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4069 = 7'h13 == r_count_39_io_out ? io_r_19_b : _GEN_4068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4070 = 7'h14 == r_count_39_io_out ? io_r_20_b : _GEN_4069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4071 = 7'h15 == r_count_39_io_out ? io_r_21_b : _GEN_4070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4072 = 7'h16 == r_count_39_io_out ? io_r_22_b : _GEN_4071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4073 = 7'h17 == r_count_39_io_out ? io_r_23_b : _GEN_4072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4074 = 7'h18 == r_count_39_io_out ? io_r_24_b : _GEN_4073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4075 = 7'h19 == r_count_39_io_out ? io_r_25_b : _GEN_4074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4076 = 7'h1a == r_count_39_io_out ? io_r_26_b : _GEN_4075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4077 = 7'h1b == r_count_39_io_out ? io_r_27_b : _GEN_4076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4078 = 7'h1c == r_count_39_io_out ? io_r_28_b : _GEN_4077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4079 = 7'h1d == r_count_39_io_out ? io_r_29_b : _GEN_4078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4080 = 7'h1e == r_count_39_io_out ? io_r_30_b : _GEN_4079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4081 = 7'h1f == r_count_39_io_out ? io_r_31_b : _GEN_4080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4082 = 7'h20 == r_count_39_io_out ? io_r_32_b : _GEN_4081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4083 = 7'h21 == r_count_39_io_out ? io_r_33_b : _GEN_4082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4084 = 7'h22 == r_count_39_io_out ? io_r_34_b : _GEN_4083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4085 = 7'h23 == r_count_39_io_out ? io_r_35_b : _GEN_4084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4086 = 7'h24 == r_count_39_io_out ? io_r_36_b : _GEN_4085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4087 = 7'h25 == r_count_39_io_out ? io_r_37_b : _GEN_4086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4088 = 7'h26 == r_count_39_io_out ? io_r_38_b : _GEN_4087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4089 = 7'h27 == r_count_39_io_out ? io_r_39_b : _GEN_4088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4090 = 7'h28 == r_count_39_io_out ? io_r_40_b : _GEN_4089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4091 = 7'h29 == r_count_39_io_out ? io_r_41_b : _GEN_4090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4092 = 7'h2a == r_count_39_io_out ? io_r_42_b : _GEN_4091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4093 = 7'h2b == r_count_39_io_out ? io_r_43_b : _GEN_4092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4094 = 7'h2c == r_count_39_io_out ? io_r_44_b : _GEN_4093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4095 = 7'h2d == r_count_39_io_out ? io_r_45_b : _GEN_4094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4096 = 7'h2e == r_count_39_io_out ? io_r_46_b : _GEN_4095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4097 = 7'h2f == r_count_39_io_out ? io_r_47_b : _GEN_4096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4098 = 7'h30 == r_count_39_io_out ? io_r_48_b : _GEN_4097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4099 = 7'h31 == r_count_39_io_out ? io_r_49_b : _GEN_4098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4100 = 7'h32 == r_count_39_io_out ? io_r_50_b : _GEN_4099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4101 = 7'h33 == r_count_39_io_out ? io_r_51_b : _GEN_4100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4102 = 7'h34 == r_count_39_io_out ? io_r_52_b : _GEN_4101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4103 = 7'h35 == r_count_39_io_out ? io_r_53_b : _GEN_4102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4104 = 7'h36 == r_count_39_io_out ? io_r_54_b : _GEN_4103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4105 = 7'h37 == r_count_39_io_out ? io_r_55_b : _GEN_4104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4106 = 7'h38 == r_count_39_io_out ? io_r_56_b : _GEN_4105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4107 = 7'h39 == r_count_39_io_out ? io_r_57_b : _GEN_4106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4108 = 7'h3a == r_count_39_io_out ? io_r_58_b : _GEN_4107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4109 = 7'h3b == r_count_39_io_out ? io_r_59_b : _GEN_4108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4110 = 7'h3c == r_count_39_io_out ? io_r_60_b : _GEN_4109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4111 = 7'h3d == r_count_39_io_out ? io_r_61_b : _GEN_4110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4112 = 7'h3e == r_count_39_io_out ? io_r_62_b : _GEN_4111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4113 = 7'h3f == r_count_39_io_out ? io_r_63_b : _GEN_4112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4114 = 7'h40 == r_count_39_io_out ? io_r_64_b : _GEN_4113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4115 = 7'h41 == r_count_39_io_out ? io_r_65_b : _GEN_4114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4116 = 7'h42 == r_count_39_io_out ? io_r_66_b : _GEN_4115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4117 = 7'h43 == r_count_39_io_out ? io_r_67_b : _GEN_4116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4118 = 7'h44 == r_count_39_io_out ? io_r_68_b : _GEN_4117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4119 = 7'h45 == r_count_39_io_out ? io_r_69_b : _GEN_4118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4120 = 7'h46 == r_count_39_io_out ? io_r_70_b : _GEN_4119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4121 = 7'h47 == r_count_39_io_out ? io_r_71_b : _GEN_4120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4122 = 7'h48 == r_count_39_io_out ? io_r_72_b : _GEN_4121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4123 = 7'h49 == r_count_39_io_out ? io_r_73_b : _GEN_4122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4124 = 7'h4a == r_count_39_io_out ? io_r_74_b : _GEN_4123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4125 = 7'h4b == r_count_39_io_out ? io_r_75_b : _GEN_4124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4126 = 7'h4c == r_count_39_io_out ? io_r_76_b : _GEN_4125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4127 = 7'h4d == r_count_39_io_out ? io_r_77_b : _GEN_4126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4128 = 7'h4e == r_count_39_io_out ? io_r_78_b : _GEN_4127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4129 = 7'h4f == r_count_39_io_out ? io_r_79_b : _GEN_4128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4130 = 7'h50 == r_count_39_io_out ? io_r_80_b : _GEN_4129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4131 = 7'h51 == r_count_39_io_out ? io_r_81_b : _GEN_4130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4132 = 7'h52 == r_count_39_io_out ? io_r_82_b : _GEN_4131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4133 = 7'h53 == r_count_39_io_out ? io_r_83_b : _GEN_4132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4134 = 7'h54 == r_count_39_io_out ? io_r_84_b : _GEN_4133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4135 = 7'h55 == r_count_39_io_out ? io_r_85_b : _GEN_4134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4136 = 7'h56 == r_count_39_io_out ? io_r_86_b : _GEN_4135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4137 = 7'h57 == r_count_39_io_out ? io_r_87_b : _GEN_4136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4138 = 7'h58 == r_count_39_io_out ? io_r_88_b : _GEN_4137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4139 = 7'h59 == r_count_39_io_out ? io_r_89_b : _GEN_4138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4140 = 7'h5a == r_count_39_io_out ? io_r_90_b : _GEN_4139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4141 = 7'h5b == r_count_39_io_out ? io_r_91_b : _GEN_4140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4142 = 7'h5c == r_count_39_io_out ? io_r_92_b : _GEN_4141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4143 = 7'h5d == r_count_39_io_out ? io_r_93_b : _GEN_4142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4144 = 7'h5e == r_count_39_io_out ? io_r_94_b : _GEN_4143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4145 = 7'h5f == r_count_39_io_out ? io_r_95_b : _GEN_4144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4146 = 7'h60 == r_count_39_io_out ? io_r_96_b : _GEN_4145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4147 = 7'h61 == r_count_39_io_out ? io_r_97_b : _GEN_4146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4148 = 7'h62 == r_count_39_io_out ? io_r_98_b : _GEN_4147; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4151 = 7'h1 == r_count_40_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4152 = 7'h2 == r_count_40_io_out ? io_r_2_b : _GEN_4151; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4153 = 7'h3 == r_count_40_io_out ? io_r_3_b : _GEN_4152; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4154 = 7'h4 == r_count_40_io_out ? io_r_4_b : _GEN_4153; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4155 = 7'h5 == r_count_40_io_out ? io_r_5_b : _GEN_4154; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4156 = 7'h6 == r_count_40_io_out ? io_r_6_b : _GEN_4155; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4157 = 7'h7 == r_count_40_io_out ? io_r_7_b : _GEN_4156; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4158 = 7'h8 == r_count_40_io_out ? io_r_8_b : _GEN_4157; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4159 = 7'h9 == r_count_40_io_out ? io_r_9_b : _GEN_4158; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4160 = 7'ha == r_count_40_io_out ? io_r_10_b : _GEN_4159; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4161 = 7'hb == r_count_40_io_out ? io_r_11_b : _GEN_4160; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4162 = 7'hc == r_count_40_io_out ? io_r_12_b : _GEN_4161; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4163 = 7'hd == r_count_40_io_out ? io_r_13_b : _GEN_4162; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4164 = 7'he == r_count_40_io_out ? io_r_14_b : _GEN_4163; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4165 = 7'hf == r_count_40_io_out ? io_r_15_b : _GEN_4164; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4166 = 7'h10 == r_count_40_io_out ? io_r_16_b : _GEN_4165; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4167 = 7'h11 == r_count_40_io_out ? io_r_17_b : _GEN_4166; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4168 = 7'h12 == r_count_40_io_out ? io_r_18_b : _GEN_4167; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4169 = 7'h13 == r_count_40_io_out ? io_r_19_b : _GEN_4168; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4170 = 7'h14 == r_count_40_io_out ? io_r_20_b : _GEN_4169; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4171 = 7'h15 == r_count_40_io_out ? io_r_21_b : _GEN_4170; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4172 = 7'h16 == r_count_40_io_out ? io_r_22_b : _GEN_4171; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4173 = 7'h17 == r_count_40_io_out ? io_r_23_b : _GEN_4172; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4174 = 7'h18 == r_count_40_io_out ? io_r_24_b : _GEN_4173; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4175 = 7'h19 == r_count_40_io_out ? io_r_25_b : _GEN_4174; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4176 = 7'h1a == r_count_40_io_out ? io_r_26_b : _GEN_4175; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4177 = 7'h1b == r_count_40_io_out ? io_r_27_b : _GEN_4176; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4178 = 7'h1c == r_count_40_io_out ? io_r_28_b : _GEN_4177; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4179 = 7'h1d == r_count_40_io_out ? io_r_29_b : _GEN_4178; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4180 = 7'h1e == r_count_40_io_out ? io_r_30_b : _GEN_4179; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4181 = 7'h1f == r_count_40_io_out ? io_r_31_b : _GEN_4180; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4182 = 7'h20 == r_count_40_io_out ? io_r_32_b : _GEN_4181; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4183 = 7'h21 == r_count_40_io_out ? io_r_33_b : _GEN_4182; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4184 = 7'h22 == r_count_40_io_out ? io_r_34_b : _GEN_4183; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4185 = 7'h23 == r_count_40_io_out ? io_r_35_b : _GEN_4184; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4186 = 7'h24 == r_count_40_io_out ? io_r_36_b : _GEN_4185; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4187 = 7'h25 == r_count_40_io_out ? io_r_37_b : _GEN_4186; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4188 = 7'h26 == r_count_40_io_out ? io_r_38_b : _GEN_4187; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4189 = 7'h27 == r_count_40_io_out ? io_r_39_b : _GEN_4188; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4190 = 7'h28 == r_count_40_io_out ? io_r_40_b : _GEN_4189; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4191 = 7'h29 == r_count_40_io_out ? io_r_41_b : _GEN_4190; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4192 = 7'h2a == r_count_40_io_out ? io_r_42_b : _GEN_4191; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4193 = 7'h2b == r_count_40_io_out ? io_r_43_b : _GEN_4192; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4194 = 7'h2c == r_count_40_io_out ? io_r_44_b : _GEN_4193; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4195 = 7'h2d == r_count_40_io_out ? io_r_45_b : _GEN_4194; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4196 = 7'h2e == r_count_40_io_out ? io_r_46_b : _GEN_4195; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4197 = 7'h2f == r_count_40_io_out ? io_r_47_b : _GEN_4196; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4198 = 7'h30 == r_count_40_io_out ? io_r_48_b : _GEN_4197; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4199 = 7'h31 == r_count_40_io_out ? io_r_49_b : _GEN_4198; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4200 = 7'h32 == r_count_40_io_out ? io_r_50_b : _GEN_4199; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4201 = 7'h33 == r_count_40_io_out ? io_r_51_b : _GEN_4200; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4202 = 7'h34 == r_count_40_io_out ? io_r_52_b : _GEN_4201; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4203 = 7'h35 == r_count_40_io_out ? io_r_53_b : _GEN_4202; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4204 = 7'h36 == r_count_40_io_out ? io_r_54_b : _GEN_4203; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4205 = 7'h37 == r_count_40_io_out ? io_r_55_b : _GEN_4204; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4206 = 7'h38 == r_count_40_io_out ? io_r_56_b : _GEN_4205; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4207 = 7'h39 == r_count_40_io_out ? io_r_57_b : _GEN_4206; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4208 = 7'h3a == r_count_40_io_out ? io_r_58_b : _GEN_4207; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4209 = 7'h3b == r_count_40_io_out ? io_r_59_b : _GEN_4208; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4210 = 7'h3c == r_count_40_io_out ? io_r_60_b : _GEN_4209; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4211 = 7'h3d == r_count_40_io_out ? io_r_61_b : _GEN_4210; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4212 = 7'h3e == r_count_40_io_out ? io_r_62_b : _GEN_4211; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4213 = 7'h3f == r_count_40_io_out ? io_r_63_b : _GEN_4212; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4214 = 7'h40 == r_count_40_io_out ? io_r_64_b : _GEN_4213; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4215 = 7'h41 == r_count_40_io_out ? io_r_65_b : _GEN_4214; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4216 = 7'h42 == r_count_40_io_out ? io_r_66_b : _GEN_4215; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4217 = 7'h43 == r_count_40_io_out ? io_r_67_b : _GEN_4216; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4218 = 7'h44 == r_count_40_io_out ? io_r_68_b : _GEN_4217; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4219 = 7'h45 == r_count_40_io_out ? io_r_69_b : _GEN_4218; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4220 = 7'h46 == r_count_40_io_out ? io_r_70_b : _GEN_4219; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4221 = 7'h47 == r_count_40_io_out ? io_r_71_b : _GEN_4220; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4222 = 7'h48 == r_count_40_io_out ? io_r_72_b : _GEN_4221; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4223 = 7'h49 == r_count_40_io_out ? io_r_73_b : _GEN_4222; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4224 = 7'h4a == r_count_40_io_out ? io_r_74_b : _GEN_4223; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4225 = 7'h4b == r_count_40_io_out ? io_r_75_b : _GEN_4224; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4226 = 7'h4c == r_count_40_io_out ? io_r_76_b : _GEN_4225; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4227 = 7'h4d == r_count_40_io_out ? io_r_77_b : _GEN_4226; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4228 = 7'h4e == r_count_40_io_out ? io_r_78_b : _GEN_4227; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4229 = 7'h4f == r_count_40_io_out ? io_r_79_b : _GEN_4228; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4230 = 7'h50 == r_count_40_io_out ? io_r_80_b : _GEN_4229; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4231 = 7'h51 == r_count_40_io_out ? io_r_81_b : _GEN_4230; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4232 = 7'h52 == r_count_40_io_out ? io_r_82_b : _GEN_4231; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4233 = 7'h53 == r_count_40_io_out ? io_r_83_b : _GEN_4232; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4234 = 7'h54 == r_count_40_io_out ? io_r_84_b : _GEN_4233; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4235 = 7'h55 == r_count_40_io_out ? io_r_85_b : _GEN_4234; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4236 = 7'h56 == r_count_40_io_out ? io_r_86_b : _GEN_4235; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4237 = 7'h57 == r_count_40_io_out ? io_r_87_b : _GEN_4236; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4238 = 7'h58 == r_count_40_io_out ? io_r_88_b : _GEN_4237; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4239 = 7'h59 == r_count_40_io_out ? io_r_89_b : _GEN_4238; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4240 = 7'h5a == r_count_40_io_out ? io_r_90_b : _GEN_4239; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4241 = 7'h5b == r_count_40_io_out ? io_r_91_b : _GEN_4240; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4242 = 7'h5c == r_count_40_io_out ? io_r_92_b : _GEN_4241; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4243 = 7'h5d == r_count_40_io_out ? io_r_93_b : _GEN_4242; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4244 = 7'h5e == r_count_40_io_out ? io_r_94_b : _GEN_4243; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4245 = 7'h5f == r_count_40_io_out ? io_r_95_b : _GEN_4244; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4246 = 7'h60 == r_count_40_io_out ? io_r_96_b : _GEN_4245; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4247 = 7'h61 == r_count_40_io_out ? io_r_97_b : _GEN_4246; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4248 = 7'h62 == r_count_40_io_out ? io_r_98_b : _GEN_4247; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4251 = 7'h1 == r_count_41_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4252 = 7'h2 == r_count_41_io_out ? io_r_2_b : _GEN_4251; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4253 = 7'h3 == r_count_41_io_out ? io_r_3_b : _GEN_4252; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4254 = 7'h4 == r_count_41_io_out ? io_r_4_b : _GEN_4253; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4255 = 7'h5 == r_count_41_io_out ? io_r_5_b : _GEN_4254; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4256 = 7'h6 == r_count_41_io_out ? io_r_6_b : _GEN_4255; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4257 = 7'h7 == r_count_41_io_out ? io_r_7_b : _GEN_4256; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4258 = 7'h8 == r_count_41_io_out ? io_r_8_b : _GEN_4257; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4259 = 7'h9 == r_count_41_io_out ? io_r_9_b : _GEN_4258; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4260 = 7'ha == r_count_41_io_out ? io_r_10_b : _GEN_4259; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4261 = 7'hb == r_count_41_io_out ? io_r_11_b : _GEN_4260; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4262 = 7'hc == r_count_41_io_out ? io_r_12_b : _GEN_4261; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4263 = 7'hd == r_count_41_io_out ? io_r_13_b : _GEN_4262; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4264 = 7'he == r_count_41_io_out ? io_r_14_b : _GEN_4263; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4265 = 7'hf == r_count_41_io_out ? io_r_15_b : _GEN_4264; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4266 = 7'h10 == r_count_41_io_out ? io_r_16_b : _GEN_4265; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4267 = 7'h11 == r_count_41_io_out ? io_r_17_b : _GEN_4266; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4268 = 7'h12 == r_count_41_io_out ? io_r_18_b : _GEN_4267; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4269 = 7'h13 == r_count_41_io_out ? io_r_19_b : _GEN_4268; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4270 = 7'h14 == r_count_41_io_out ? io_r_20_b : _GEN_4269; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4271 = 7'h15 == r_count_41_io_out ? io_r_21_b : _GEN_4270; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4272 = 7'h16 == r_count_41_io_out ? io_r_22_b : _GEN_4271; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4273 = 7'h17 == r_count_41_io_out ? io_r_23_b : _GEN_4272; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4274 = 7'h18 == r_count_41_io_out ? io_r_24_b : _GEN_4273; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4275 = 7'h19 == r_count_41_io_out ? io_r_25_b : _GEN_4274; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4276 = 7'h1a == r_count_41_io_out ? io_r_26_b : _GEN_4275; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4277 = 7'h1b == r_count_41_io_out ? io_r_27_b : _GEN_4276; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4278 = 7'h1c == r_count_41_io_out ? io_r_28_b : _GEN_4277; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4279 = 7'h1d == r_count_41_io_out ? io_r_29_b : _GEN_4278; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4280 = 7'h1e == r_count_41_io_out ? io_r_30_b : _GEN_4279; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4281 = 7'h1f == r_count_41_io_out ? io_r_31_b : _GEN_4280; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4282 = 7'h20 == r_count_41_io_out ? io_r_32_b : _GEN_4281; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4283 = 7'h21 == r_count_41_io_out ? io_r_33_b : _GEN_4282; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4284 = 7'h22 == r_count_41_io_out ? io_r_34_b : _GEN_4283; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4285 = 7'h23 == r_count_41_io_out ? io_r_35_b : _GEN_4284; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4286 = 7'h24 == r_count_41_io_out ? io_r_36_b : _GEN_4285; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4287 = 7'h25 == r_count_41_io_out ? io_r_37_b : _GEN_4286; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4288 = 7'h26 == r_count_41_io_out ? io_r_38_b : _GEN_4287; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4289 = 7'h27 == r_count_41_io_out ? io_r_39_b : _GEN_4288; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4290 = 7'h28 == r_count_41_io_out ? io_r_40_b : _GEN_4289; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4291 = 7'h29 == r_count_41_io_out ? io_r_41_b : _GEN_4290; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4292 = 7'h2a == r_count_41_io_out ? io_r_42_b : _GEN_4291; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4293 = 7'h2b == r_count_41_io_out ? io_r_43_b : _GEN_4292; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4294 = 7'h2c == r_count_41_io_out ? io_r_44_b : _GEN_4293; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4295 = 7'h2d == r_count_41_io_out ? io_r_45_b : _GEN_4294; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4296 = 7'h2e == r_count_41_io_out ? io_r_46_b : _GEN_4295; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4297 = 7'h2f == r_count_41_io_out ? io_r_47_b : _GEN_4296; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4298 = 7'h30 == r_count_41_io_out ? io_r_48_b : _GEN_4297; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4299 = 7'h31 == r_count_41_io_out ? io_r_49_b : _GEN_4298; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4300 = 7'h32 == r_count_41_io_out ? io_r_50_b : _GEN_4299; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4301 = 7'h33 == r_count_41_io_out ? io_r_51_b : _GEN_4300; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4302 = 7'h34 == r_count_41_io_out ? io_r_52_b : _GEN_4301; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4303 = 7'h35 == r_count_41_io_out ? io_r_53_b : _GEN_4302; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4304 = 7'h36 == r_count_41_io_out ? io_r_54_b : _GEN_4303; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4305 = 7'h37 == r_count_41_io_out ? io_r_55_b : _GEN_4304; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4306 = 7'h38 == r_count_41_io_out ? io_r_56_b : _GEN_4305; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4307 = 7'h39 == r_count_41_io_out ? io_r_57_b : _GEN_4306; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4308 = 7'h3a == r_count_41_io_out ? io_r_58_b : _GEN_4307; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4309 = 7'h3b == r_count_41_io_out ? io_r_59_b : _GEN_4308; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4310 = 7'h3c == r_count_41_io_out ? io_r_60_b : _GEN_4309; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4311 = 7'h3d == r_count_41_io_out ? io_r_61_b : _GEN_4310; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4312 = 7'h3e == r_count_41_io_out ? io_r_62_b : _GEN_4311; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4313 = 7'h3f == r_count_41_io_out ? io_r_63_b : _GEN_4312; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4314 = 7'h40 == r_count_41_io_out ? io_r_64_b : _GEN_4313; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4315 = 7'h41 == r_count_41_io_out ? io_r_65_b : _GEN_4314; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4316 = 7'h42 == r_count_41_io_out ? io_r_66_b : _GEN_4315; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4317 = 7'h43 == r_count_41_io_out ? io_r_67_b : _GEN_4316; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4318 = 7'h44 == r_count_41_io_out ? io_r_68_b : _GEN_4317; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4319 = 7'h45 == r_count_41_io_out ? io_r_69_b : _GEN_4318; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4320 = 7'h46 == r_count_41_io_out ? io_r_70_b : _GEN_4319; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4321 = 7'h47 == r_count_41_io_out ? io_r_71_b : _GEN_4320; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4322 = 7'h48 == r_count_41_io_out ? io_r_72_b : _GEN_4321; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4323 = 7'h49 == r_count_41_io_out ? io_r_73_b : _GEN_4322; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4324 = 7'h4a == r_count_41_io_out ? io_r_74_b : _GEN_4323; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4325 = 7'h4b == r_count_41_io_out ? io_r_75_b : _GEN_4324; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4326 = 7'h4c == r_count_41_io_out ? io_r_76_b : _GEN_4325; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4327 = 7'h4d == r_count_41_io_out ? io_r_77_b : _GEN_4326; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4328 = 7'h4e == r_count_41_io_out ? io_r_78_b : _GEN_4327; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4329 = 7'h4f == r_count_41_io_out ? io_r_79_b : _GEN_4328; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4330 = 7'h50 == r_count_41_io_out ? io_r_80_b : _GEN_4329; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4331 = 7'h51 == r_count_41_io_out ? io_r_81_b : _GEN_4330; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4332 = 7'h52 == r_count_41_io_out ? io_r_82_b : _GEN_4331; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4333 = 7'h53 == r_count_41_io_out ? io_r_83_b : _GEN_4332; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4334 = 7'h54 == r_count_41_io_out ? io_r_84_b : _GEN_4333; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4335 = 7'h55 == r_count_41_io_out ? io_r_85_b : _GEN_4334; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4336 = 7'h56 == r_count_41_io_out ? io_r_86_b : _GEN_4335; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4337 = 7'h57 == r_count_41_io_out ? io_r_87_b : _GEN_4336; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4338 = 7'h58 == r_count_41_io_out ? io_r_88_b : _GEN_4337; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4339 = 7'h59 == r_count_41_io_out ? io_r_89_b : _GEN_4338; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4340 = 7'h5a == r_count_41_io_out ? io_r_90_b : _GEN_4339; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4341 = 7'h5b == r_count_41_io_out ? io_r_91_b : _GEN_4340; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4342 = 7'h5c == r_count_41_io_out ? io_r_92_b : _GEN_4341; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4343 = 7'h5d == r_count_41_io_out ? io_r_93_b : _GEN_4342; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4344 = 7'h5e == r_count_41_io_out ? io_r_94_b : _GEN_4343; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4345 = 7'h5f == r_count_41_io_out ? io_r_95_b : _GEN_4344; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4346 = 7'h60 == r_count_41_io_out ? io_r_96_b : _GEN_4345; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4347 = 7'h61 == r_count_41_io_out ? io_r_97_b : _GEN_4346; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4348 = 7'h62 == r_count_41_io_out ? io_r_98_b : _GEN_4347; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4351 = 7'h1 == r_count_42_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4352 = 7'h2 == r_count_42_io_out ? io_r_2_b : _GEN_4351; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4353 = 7'h3 == r_count_42_io_out ? io_r_3_b : _GEN_4352; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4354 = 7'h4 == r_count_42_io_out ? io_r_4_b : _GEN_4353; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4355 = 7'h5 == r_count_42_io_out ? io_r_5_b : _GEN_4354; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4356 = 7'h6 == r_count_42_io_out ? io_r_6_b : _GEN_4355; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4357 = 7'h7 == r_count_42_io_out ? io_r_7_b : _GEN_4356; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4358 = 7'h8 == r_count_42_io_out ? io_r_8_b : _GEN_4357; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4359 = 7'h9 == r_count_42_io_out ? io_r_9_b : _GEN_4358; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4360 = 7'ha == r_count_42_io_out ? io_r_10_b : _GEN_4359; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4361 = 7'hb == r_count_42_io_out ? io_r_11_b : _GEN_4360; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4362 = 7'hc == r_count_42_io_out ? io_r_12_b : _GEN_4361; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4363 = 7'hd == r_count_42_io_out ? io_r_13_b : _GEN_4362; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4364 = 7'he == r_count_42_io_out ? io_r_14_b : _GEN_4363; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4365 = 7'hf == r_count_42_io_out ? io_r_15_b : _GEN_4364; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4366 = 7'h10 == r_count_42_io_out ? io_r_16_b : _GEN_4365; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4367 = 7'h11 == r_count_42_io_out ? io_r_17_b : _GEN_4366; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4368 = 7'h12 == r_count_42_io_out ? io_r_18_b : _GEN_4367; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4369 = 7'h13 == r_count_42_io_out ? io_r_19_b : _GEN_4368; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4370 = 7'h14 == r_count_42_io_out ? io_r_20_b : _GEN_4369; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4371 = 7'h15 == r_count_42_io_out ? io_r_21_b : _GEN_4370; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4372 = 7'h16 == r_count_42_io_out ? io_r_22_b : _GEN_4371; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4373 = 7'h17 == r_count_42_io_out ? io_r_23_b : _GEN_4372; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4374 = 7'h18 == r_count_42_io_out ? io_r_24_b : _GEN_4373; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4375 = 7'h19 == r_count_42_io_out ? io_r_25_b : _GEN_4374; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4376 = 7'h1a == r_count_42_io_out ? io_r_26_b : _GEN_4375; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4377 = 7'h1b == r_count_42_io_out ? io_r_27_b : _GEN_4376; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4378 = 7'h1c == r_count_42_io_out ? io_r_28_b : _GEN_4377; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4379 = 7'h1d == r_count_42_io_out ? io_r_29_b : _GEN_4378; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4380 = 7'h1e == r_count_42_io_out ? io_r_30_b : _GEN_4379; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4381 = 7'h1f == r_count_42_io_out ? io_r_31_b : _GEN_4380; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4382 = 7'h20 == r_count_42_io_out ? io_r_32_b : _GEN_4381; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4383 = 7'h21 == r_count_42_io_out ? io_r_33_b : _GEN_4382; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4384 = 7'h22 == r_count_42_io_out ? io_r_34_b : _GEN_4383; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4385 = 7'h23 == r_count_42_io_out ? io_r_35_b : _GEN_4384; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4386 = 7'h24 == r_count_42_io_out ? io_r_36_b : _GEN_4385; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4387 = 7'h25 == r_count_42_io_out ? io_r_37_b : _GEN_4386; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4388 = 7'h26 == r_count_42_io_out ? io_r_38_b : _GEN_4387; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4389 = 7'h27 == r_count_42_io_out ? io_r_39_b : _GEN_4388; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4390 = 7'h28 == r_count_42_io_out ? io_r_40_b : _GEN_4389; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4391 = 7'h29 == r_count_42_io_out ? io_r_41_b : _GEN_4390; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4392 = 7'h2a == r_count_42_io_out ? io_r_42_b : _GEN_4391; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4393 = 7'h2b == r_count_42_io_out ? io_r_43_b : _GEN_4392; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4394 = 7'h2c == r_count_42_io_out ? io_r_44_b : _GEN_4393; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4395 = 7'h2d == r_count_42_io_out ? io_r_45_b : _GEN_4394; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4396 = 7'h2e == r_count_42_io_out ? io_r_46_b : _GEN_4395; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4397 = 7'h2f == r_count_42_io_out ? io_r_47_b : _GEN_4396; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4398 = 7'h30 == r_count_42_io_out ? io_r_48_b : _GEN_4397; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4399 = 7'h31 == r_count_42_io_out ? io_r_49_b : _GEN_4398; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4400 = 7'h32 == r_count_42_io_out ? io_r_50_b : _GEN_4399; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4401 = 7'h33 == r_count_42_io_out ? io_r_51_b : _GEN_4400; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4402 = 7'h34 == r_count_42_io_out ? io_r_52_b : _GEN_4401; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4403 = 7'h35 == r_count_42_io_out ? io_r_53_b : _GEN_4402; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4404 = 7'h36 == r_count_42_io_out ? io_r_54_b : _GEN_4403; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4405 = 7'h37 == r_count_42_io_out ? io_r_55_b : _GEN_4404; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4406 = 7'h38 == r_count_42_io_out ? io_r_56_b : _GEN_4405; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4407 = 7'h39 == r_count_42_io_out ? io_r_57_b : _GEN_4406; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4408 = 7'h3a == r_count_42_io_out ? io_r_58_b : _GEN_4407; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4409 = 7'h3b == r_count_42_io_out ? io_r_59_b : _GEN_4408; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4410 = 7'h3c == r_count_42_io_out ? io_r_60_b : _GEN_4409; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4411 = 7'h3d == r_count_42_io_out ? io_r_61_b : _GEN_4410; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4412 = 7'h3e == r_count_42_io_out ? io_r_62_b : _GEN_4411; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4413 = 7'h3f == r_count_42_io_out ? io_r_63_b : _GEN_4412; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4414 = 7'h40 == r_count_42_io_out ? io_r_64_b : _GEN_4413; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4415 = 7'h41 == r_count_42_io_out ? io_r_65_b : _GEN_4414; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4416 = 7'h42 == r_count_42_io_out ? io_r_66_b : _GEN_4415; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4417 = 7'h43 == r_count_42_io_out ? io_r_67_b : _GEN_4416; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4418 = 7'h44 == r_count_42_io_out ? io_r_68_b : _GEN_4417; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4419 = 7'h45 == r_count_42_io_out ? io_r_69_b : _GEN_4418; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4420 = 7'h46 == r_count_42_io_out ? io_r_70_b : _GEN_4419; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4421 = 7'h47 == r_count_42_io_out ? io_r_71_b : _GEN_4420; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4422 = 7'h48 == r_count_42_io_out ? io_r_72_b : _GEN_4421; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4423 = 7'h49 == r_count_42_io_out ? io_r_73_b : _GEN_4422; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4424 = 7'h4a == r_count_42_io_out ? io_r_74_b : _GEN_4423; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4425 = 7'h4b == r_count_42_io_out ? io_r_75_b : _GEN_4424; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4426 = 7'h4c == r_count_42_io_out ? io_r_76_b : _GEN_4425; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4427 = 7'h4d == r_count_42_io_out ? io_r_77_b : _GEN_4426; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4428 = 7'h4e == r_count_42_io_out ? io_r_78_b : _GEN_4427; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4429 = 7'h4f == r_count_42_io_out ? io_r_79_b : _GEN_4428; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4430 = 7'h50 == r_count_42_io_out ? io_r_80_b : _GEN_4429; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4431 = 7'h51 == r_count_42_io_out ? io_r_81_b : _GEN_4430; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4432 = 7'h52 == r_count_42_io_out ? io_r_82_b : _GEN_4431; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4433 = 7'h53 == r_count_42_io_out ? io_r_83_b : _GEN_4432; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4434 = 7'h54 == r_count_42_io_out ? io_r_84_b : _GEN_4433; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4435 = 7'h55 == r_count_42_io_out ? io_r_85_b : _GEN_4434; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4436 = 7'h56 == r_count_42_io_out ? io_r_86_b : _GEN_4435; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4437 = 7'h57 == r_count_42_io_out ? io_r_87_b : _GEN_4436; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4438 = 7'h58 == r_count_42_io_out ? io_r_88_b : _GEN_4437; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4439 = 7'h59 == r_count_42_io_out ? io_r_89_b : _GEN_4438; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4440 = 7'h5a == r_count_42_io_out ? io_r_90_b : _GEN_4439; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4441 = 7'h5b == r_count_42_io_out ? io_r_91_b : _GEN_4440; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4442 = 7'h5c == r_count_42_io_out ? io_r_92_b : _GEN_4441; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4443 = 7'h5d == r_count_42_io_out ? io_r_93_b : _GEN_4442; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4444 = 7'h5e == r_count_42_io_out ? io_r_94_b : _GEN_4443; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4445 = 7'h5f == r_count_42_io_out ? io_r_95_b : _GEN_4444; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4446 = 7'h60 == r_count_42_io_out ? io_r_96_b : _GEN_4445; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4447 = 7'h61 == r_count_42_io_out ? io_r_97_b : _GEN_4446; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4448 = 7'h62 == r_count_42_io_out ? io_r_98_b : _GEN_4447; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4451 = 7'h1 == r_count_43_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4452 = 7'h2 == r_count_43_io_out ? io_r_2_b : _GEN_4451; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4453 = 7'h3 == r_count_43_io_out ? io_r_3_b : _GEN_4452; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4454 = 7'h4 == r_count_43_io_out ? io_r_4_b : _GEN_4453; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4455 = 7'h5 == r_count_43_io_out ? io_r_5_b : _GEN_4454; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4456 = 7'h6 == r_count_43_io_out ? io_r_6_b : _GEN_4455; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4457 = 7'h7 == r_count_43_io_out ? io_r_7_b : _GEN_4456; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4458 = 7'h8 == r_count_43_io_out ? io_r_8_b : _GEN_4457; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4459 = 7'h9 == r_count_43_io_out ? io_r_9_b : _GEN_4458; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4460 = 7'ha == r_count_43_io_out ? io_r_10_b : _GEN_4459; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4461 = 7'hb == r_count_43_io_out ? io_r_11_b : _GEN_4460; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4462 = 7'hc == r_count_43_io_out ? io_r_12_b : _GEN_4461; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4463 = 7'hd == r_count_43_io_out ? io_r_13_b : _GEN_4462; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4464 = 7'he == r_count_43_io_out ? io_r_14_b : _GEN_4463; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4465 = 7'hf == r_count_43_io_out ? io_r_15_b : _GEN_4464; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4466 = 7'h10 == r_count_43_io_out ? io_r_16_b : _GEN_4465; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4467 = 7'h11 == r_count_43_io_out ? io_r_17_b : _GEN_4466; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4468 = 7'h12 == r_count_43_io_out ? io_r_18_b : _GEN_4467; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4469 = 7'h13 == r_count_43_io_out ? io_r_19_b : _GEN_4468; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4470 = 7'h14 == r_count_43_io_out ? io_r_20_b : _GEN_4469; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4471 = 7'h15 == r_count_43_io_out ? io_r_21_b : _GEN_4470; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4472 = 7'h16 == r_count_43_io_out ? io_r_22_b : _GEN_4471; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4473 = 7'h17 == r_count_43_io_out ? io_r_23_b : _GEN_4472; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4474 = 7'h18 == r_count_43_io_out ? io_r_24_b : _GEN_4473; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4475 = 7'h19 == r_count_43_io_out ? io_r_25_b : _GEN_4474; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4476 = 7'h1a == r_count_43_io_out ? io_r_26_b : _GEN_4475; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4477 = 7'h1b == r_count_43_io_out ? io_r_27_b : _GEN_4476; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4478 = 7'h1c == r_count_43_io_out ? io_r_28_b : _GEN_4477; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4479 = 7'h1d == r_count_43_io_out ? io_r_29_b : _GEN_4478; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4480 = 7'h1e == r_count_43_io_out ? io_r_30_b : _GEN_4479; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4481 = 7'h1f == r_count_43_io_out ? io_r_31_b : _GEN_4480; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4482 = 7'h20 == r_count_43_io_out ? io_r_32_b : _GEN_4481; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4483 = 7'h21 == r_count_43_io_out ? io_r_33_b : _GEN_4482; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4484 = 7'h22 == r_count_43_io_out ? io_r_34_b : _GEN_4483; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4485 = 7'h23 == r_count_43_io_out ? io_r_35_b : _GEN_4484; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4486 = 7'h24 == r_count_43_io_out ? io_r_36_b : _GEN_4485; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4487 = 7'h25 == r_count_43_io_out ? io_r_37_b : _GEN_4486; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4488 = 7'h26 == r_count_43_io_out ? io_r_38_b : _GEN_4487; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4489 = 7'h27 == r_count_43_io_out ? io_r_39_b : _GEN_4488; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4490 = 7'h28 == r_count_43_io_out ? io_r_40_b : _GEN_4489; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4491 = 7'h29 == r_count_43_io_out ? io_r_41_b : _GEN_4490; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4492 = 7'h2a == r_count_43_io_out ? io_r_42_b : _GEN_4491; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4493 = 7'h2b == r_count_43_io_out ? io_r_43_b : _GEN_4492; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4494 = 7'h2c == r_count_43_io_out ? io_r_44_b : _GEN_4493; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4495 = 7'h2d == r_count_43_io_out ? io_r_45_b : _GEN_4494; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4496 = 7'h2e == r_count_43_io_out ? io_r_46_b : _GEN_4495; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4497 = 7'h2f == r_count_43_io_out ? io_r_47_b : _GEN_4496; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4498 = 7'h30 == r_count_43_io_out ? io_r_48_b : _GEN_4497; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4499 = 7'h31 == r_count_43_io_out ? io_r_49_b : _GEN_4498; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4500 = 7'h32 == r_count_43_io_out ? io_r_50_b : _GEN_4499; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4501 = 7'h33 == r_count_43_io_out ? io_r_51_b : _GEN_4500; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4502 = 7'h34 == r_count_43_io_out ? io_r_52_b : _GEN_4501; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4503 = 7'h35 == r_count_43_io_out ? io_r_53_b : _GEN_4502; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4504 = 7'h36 == r_count_43_io_out ? io_r_54_b : _GEN_4503; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4505 = 7'h37 == r_count_43_io_out ? io_r_55_b : _GEN_4504; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4506 = 7'h38 == r_count_43_io_out ? io_r_56_b : _GEN_4505; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4507 = 7'h39 == r_count_43_io_out ? io_r_57_b : _GEN_4506; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4508 = 7'h3a == r_count_43_io_out ? io_r_58_b : _GEN_4507; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4509 = 7'h3b == r_count_43_io_out ? io_r_59_b : _GEN_4508; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4510 = 7'h3c == r_count_43_io_out ? io_r_60_b : _GEN_4509; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4511 = 7'h3d == r_count_43_io_out ? io_r_61_b : _GEN_4510; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4512 = 7'h3e == r_count_43_io_out ? io_r_62_b : _GEN_4511; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4513 = 7'h3f == r_count_43_io_out ? io_r_63_b : _GEN_4512; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4514 = 7'h40 == r_count_43_io_out ? io_r_64_b : _GEN_4513; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4515 = 7'h41 == r_count_43_io_out ? io_r_65_b : _GEN_4514; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4516 = 7'h42 == r_count_43_io_out ? io_r_66_b : _GEN_4515; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4517 = 7'h43 == r_count_43_io_out ? io_r_67_b : _GEN_4516; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4518 = 7'h44 == r_count_43_io_out ? io_r_68_b : _GEN_4517; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4519 = 7'h45 == r_count_43_io_out ? io_r_69_b : _GEN_4518; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4520 = 7'h46 == r_count_43_io_out ? io_r_70_b : _GEN_4519; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4521 = 7'h47 == r_count_43_io_out ? io_r_71_b : _GEN_4520; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4522 = 7'h48 == r_count_43_io_out ? io_r_72_b : _GEN_4521; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4523 = 7'h49 == r_count_43_io_out ? io_r_73_b : _GEN_4522; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4524 = 7'h4a == r_count_43_io_out ? io_r_74_b : _GEN_4523; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4525 = 7'h4b == r_count_43_io_out ? io_r_75_b : _GEN_4524; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4526 = 7'h4c == r_count_43_io_out ? io_r_76_b : _GEN_4525; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4527 = 7'h4d == r_count_43_io_out ? io_r_77_b : _GEN_4526; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4528 = 7'h4e == r_count_43_io_out ? io_r_78_b : _GEN_4527; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4529 = 7'h4f == r_count_43_io_out ? io_r_79_b : _GEN_4528; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4530 = 7'h50 == r_count_43_io_out ? io_r_80_b : _GEN_4529; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4531 = 7'h51 == r_count_43_io_out ? io_r_81_b : _GEN_4530; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4532 = 7'h52 == r_count_43_io_out ? io_r_82_b : _GEN_4531; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4533 = 7'h53 == r_count_43_io_out ? io_r_83_b : _GEN_4532; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4534 = 7'h54 == r_count_43_io_out ? io_r_84_b : _GEN_4533; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4535 = 7'h55 == r_count_43_io_out ? io_r_85_b : _GEN_4534; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4536 = 7'h56 == r_count_43_io_out ? io_r_86_b : _GEN_4535; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4537 = 7'h57 == r_count_43_io_out ? io_r_87_b : _GEN_4536; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4538 = 7'h58 == r_count_43_io_out ? io_r_88_b : _GEN_4537; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4539 = 7'h59 == r_count_43_io_out ? io_r_89_b : _GEN_4538; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4540 = 7'h5a == r_count_43_io_out ? io_r_90_b : _GEN_4539; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4541 = 7'h5b == r_count_43_io_out ? io_r_91_b : _GEN_4540; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4542 = 7'h5c == r_count_43_io_out ? io_r_92_b : _GEN_4541; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4543 = 7'h5d == r_count_43_io_out ? io_r_93_b : _GEN_4542; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4544 = 7'h5e == r_count_43_io_out ? io_r_94_b : _GEN_4543; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4545 = 7'h5f == r_count_43_io_out ? io_r_95_b : _GEN_4544; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4546 = 7'h60 == r_count_43_io_out ? io_r_96_b : _GEN_4545; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4547 = 7'h61 == r_count_43_io_out ? io_r_97_b : _GEN_4546; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4548 = 7'h62 == r_count_43_io_out ? io_r_98_b : _GEN_4547; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4551 = 7'h1 == r_count_44_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4552 = 7'h2 == r_count_44_io_out ? io_r_2_b : _GEN_4551; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4553 = 7'h3 == r_count_44_io_out ? io_r_3_b : _GEN_4552; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4554 = 7'h4 == r_count_44_io_out ? io_r_4_b : _GEN_4553; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4555 = 7'h5 == r_count_44_io_out ? io_r_5_b : _GEN_4554; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4556 = 7'h6 == r_count_44_io_out ? io_r_6_b : _GEN_4555; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4557 = 7'h7 == r_count_44_io_out ? io_r_7_b : _GEN_4556; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4558 = 7'h8 == r_count_44_io_out ? io_r_8_b : _GEN_4557; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4559 = 7'h9 == r_count_44_io_out ? io_r_9_b : _GEN_4558; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4560 = 7'ha == r_count_44_io_out ? io_r_10_b : _GEN_4559; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4561 = 7'hb == r_count_44_io_out ? io_r_11_b : _GEN_4560; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4562 = 7'hc == r_count_44_io_out ? io_r_12_b : _GEN_4561; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4563 = 7'hd == r_count_44_io_out ? io_r_13_b : _GEN_4562; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4564 = 7'he == r_count_44_io_out ? io_r_14_b : _GEN_4563; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4565 = 7'hf == r_count_44_io_out ? io_r_15_b : _GEN_4564; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4566 = 7'h10 == r_count_44_io_out ? io_r_16_b : _GEN_4565; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4567 = 7'h11 == r_count_44_io_out ? io_r_17_b : _GEN_4566; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4568 = 7'h12 == r_count_44_io_out ? io_r_18_b : _GEN_4567; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4569 = 7'h13 == r_count_44_io_out ? io_r_19_b : _GEN_4568; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4570 = 7'h14 == r_count_44_io_out ? io_r_20_b : _GEN_4569; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4571 = 7'h15 == r_count_44_io_out ? io_r_21_b : _GEN_4570; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4572 = 7'h16 == r_count_44_io_out ? io_r_22_b : _GEN_4571; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4573 = 7'h17 == r_count_44_io_out ? io_r_23_b : _GEN_4572; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4574 = 7'h18 == r_count_44_io_out ? io_r_24_b : _GEN_4573; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4575 = 7'h19 == r_count_44_io_out ? io_r_25_b : _GEN_4574; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4576 = 7'h1a == r_count_44_io_out ? io_r_26_b : _GEN_4575; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4577 = 7'h1b == r_count_44_io_out ? io_r_27_b : _GEN_4576; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4578 = 7'h1c == r_count_44_io_out ? io_r_28_b : _GEN_4577; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4579 = 7'h1d == r_count_44_io_out ? io_r_29_b : _GEN_4578; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4580 = 7'h1e == r_count_44_io_out ? io_r_30_b : _GEN_4579; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4581 = 7'h1f == r_count_44_io_out ? io_r_31_b : _GEN_4580; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4582 = 7'h20 == r_count_44_io_out ? io_r_32_b : _GEN_4581; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4583 = 7'h21 == r_count_44_io_out ? io_r_33_b : _GEN_4582; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4584 = 7'h22 == r_count_44_io_out ? io_r_34_b : _GEN_4583; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4585 = 7'h23 == r_count_44_io_out ? io_r_35_b : _GEN_4584; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4586 = 7'h24 == r_count_44_io_out ? io_r_36_b : _GEN_4585; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4587 = 7'h25 == r_count_44_io_out ? io_r_37_b : _GEN_4586; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4588 = 7'h26 == r_count_44_io_out ? io_r_38_b : _GEN_4587; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4589 = 7'h27 == r_count_44_io_out ? io_r_39_b : _GEN_4588; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4590 = 7'h28 == r_count_44_io_out ? io_r_40_b : _GEN_4589; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4591 = 7'h29 == r_count_44_io_out ? io_r_41_b : _GEN_4590; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4592 = 7'h2a == r_count_44_io_out ? io_r_42_b : _GEN_4591; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4593 = 7'h2b == r_count_44_io_out ? io_r_43_b : _GEN_4592; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4594 = 7'h2c == r_count_44_io_out ? io_r_44_b : _GEN_4593; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4595 = 7'h2d == r_count_44_io_out ? io_r_45_b : _GEN_4594; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4596 = 7'h2e == r_count_44_io_out ? io_r_46_b : _GEN_4595; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4597 = 7'h2f == r_count_44_io_out ? io_r_47_b : _GEN_4596; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4598 = 7'h30 == r_count_44_io_out ? io_r_48_b : _GEN_4597; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4599 = 7'h31 == r_count_44_io_out ? io_r_49_b : _GEN_4598; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4600 = 7'h32 == r_count_44_io_out ? io_r_50_b : _GEN_4599; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4601 = 7'h33 == r_count_44_io_out ? io_r_51_b : _GEN_4600; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4602 = 7'h34 == r_count_44_io_out ? io_r_52_b : _GEN_4601; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4603 = 7'h35 == r_count_44_io_out ? io_r_53_b : _GEN_4602; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4604 = 7'h36 == r_count_44_io_out ? io_r_54_b : _GEN_4603; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4605 = 7'h37 == r_count_44_io_out ? io_r_55_b : _GEN_4604; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4606 = 7'h38 == r_count_44_io_out ? io_r_56_b : _GEN_4605; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4607 = 7'h39 == r_count_44_io_out ? io_r_57_b : _GEN_4606; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4608 = 7'h3a == r_count_44_io_out ? io_r_58_b : _GEN_4607; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4609 = 7'h3b == r_count_44_io_out ? io_r_59_b : _GEN_4608; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4610 = 7'h3c == r_count_44_io_out ? io_r_60_b : _GEN_4609; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4611 = 7'h3d == r_count_44_io_out ? io_r_61_b : _GEN_4610; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4612 = 7'h3e == r_count_44_io_out ? io_r_62_b : _GEN_4611; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4613 = 7'h3f == r_count_44_io_out ? io_r_63_b : _GEN_4612; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4614 = 7'h40 == r_count_44_io_out ? io_r_64_b : _GEN_4613; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4615 = 7'h41 == r_count_44_io_out ? io_r_65_b : _GEN_4614; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4616 = 7'h42 == r_count_44_io_out ? io_r_66_b : _GEN_4615; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4617 = 7'h43 == r_count_44_io_out ? io_r_67_b : _GEN_4616; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4618 = 7'h44 == r_count_44_io_out ? io_r_68_b : _GEN_4617; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4619 = 7'h45 == r_count_44_io_out ? io_r_69_b : _GEN_4618; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4620 = 7'h46 == r_count_44_io_out ? io_r_70_b : _GEN_4619; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4621 = 7'h47 == r_count_44_io_out ? io_r_71_b : _GEN_4620; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4622 = 7'h48 == r_count_44_io_out ? io_r_72_b : _GEN_4621; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4623 = 7'h49 == r_count_44_io_out ? io_r_73_b : _GEN_4622; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4624 = 7'h4a == r_count_44_io_out ? io_r_74_b : _GEN_4623; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4625 = 7'h4b == r_count_44_io_out ? io_r_75_b : _GEN_4624; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4626 = 7'h4c == r_count_44_io_out ? io_r_76_b : _GEN_4625; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4627 = 7'h4d == r_count_44_io_out ? io_r_77_b : _GEN_4626; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4628 = 7'h4e == r_count_44_io_out ? io_r_78_b : _GEN_4627; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4629 = 7'h4f == r_count_44_io_out ? io_r_79_b : _GEN_4628; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4630 = 7'h50 == r_count_44_io_out ? io_r_80_b : _GEN_4629; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4631 = 7'h51 == r_count_44_io_out ? io_r_81_b : _GEN_4630; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4632 = 7'h52 == r_count_44_io_out ? io_r_82_b : _GEN_4631; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4633 = 7'h53 == r_count_44_io_out ? io_r_83_b : _GEN_4632; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4634 = 7'h54 == r_count_44_io_out ? io_r_84_b : _GEN_4633; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4635 = 7'h55 == r_count_44_io_out ? io_r_85_b : _GEN_4634; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4636 = 7'h56 == r_count_44_io_out ? io_r_86_b : _GEN_4635; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4637 = 7'h57 == r_count_44_io_out ? io_r_87_b : _GEN_4636; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4638 = 7'h58 == r_count_44_io_out ? io_r_88_b : _GEN_4637; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4639 = 7'h59 == r_count_44_io_out ? io_r_89_b : _GEN_4638; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4640 = 7'h5a == r_count_44_io_out ? io_r_90_b : _GEN_4639; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4641 = 7'h5b == r_count_44_io_out ? io_r_91_b : _GEN_4640; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4642 = 7'h5c == r_count_44_io_out ? io_r_92_b : _GEN_4641; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4643 = 7'h5d == r_count_44_io_out ? io_r_93_b : _GEN_4642; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4644 = 7'h5e == r_count_44_io_out ? io_r_94_b : _GEN_4643; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4645 = 7'h5f == r_count_44_io_out ? io_r_95_b : _GEN_4644; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4646 = 7'h60 == r_count_44_io_out ? io_r_96_b : _GEN_4645; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4647 = 7'h61 == r_count_44_io_out ? io_r_97_b : _GEN_4646; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4648 = 7'h62 == r_count_44_io_out ? io_r_98_b : _GEN_4647; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4651 = 7'h1 == r_count_45_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4652 = 7'h2 == r_count_45_io_out ? io_r_2_b : _GEN_4651; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4653 = 7'h3 == r_count_45_io_out ? io_r_3_b : _GEN_4652; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4654 = 7'h4 == r_count_45_io_out ? io_r_4_b : _GEN_4653; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4655 = 7'h5 == r_count_45_io_out ? io_r_5_b : _GEN_4654; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4656 = 7'h6 == r_count_45_io_out ? io_r_6_b : _GEN_4655; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4657 = 7'h7 == r_count_45_io_out ? io_r_7_b : _GEN_4656; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4658 = 7'h8 == r_count_45_io_out ? io_r_8_b : _GEN_4657; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4659 = 7'h9 == r_count_45_io_out ? io_r_9_b : _GEN_4658; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4660 = 7'ha == r_count_45_io_out ? io_r_10_b : _GEN_4659; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4661 = 7'hb == r_count_45_io_out ? io_r_11_b : _GEN_4660; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4662 = 7'hc == r_count_45_io_out ? io_r_12_b : _GEN_4661; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4663 = 7'hd == r_count_45_io_out ? io_r_13_b : _GEN_4662; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4664 = 7'he == r_count_45_io_out ? io_r_14_b : _GEN_4663; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4665 = 7'hf == r_count_45_io_out ? io_r_15_b : _GEN_4664; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4666 = 7'h10 == r_count_45_io_out ? io_r_16_b : _GEN_4665; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4667 = 7'h11 == r_count_45_io_out ? io_r_17_b : _GEN_4666; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4668 = 7'h12 == r_count_45_io_out ? io_r_18_b : _GEN_4667; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4669 = 7'h13 == r_count_45_io_out ? io_r_19_b : _GEN_4668; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4670 = 7'h14 == r_count_45_io_out ? io_r_20_b : _GEN_4669; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4671 = 7'h15 == r_count_45_io_out ? io_r_21_b : _GEN_4670; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4672 = 7'h16 == r_count_45_io_out ? io_r_22_b : _GEN_4671; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4673 = 7'h17 == r_count_45_io_out ? io_r_23_b : _GEN_4672; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4674 = 7'h18 == r_count_45_io_out ? io_r_24_b : _GEN_4673; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4675 = 7'h19 == r_count_45_io_out ? io_r_25_b : _GEN_4674; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4676 = 7'h1a == r_count_45_io_out ? io_r_26_b : _GEN_4675; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4677 = 7'h1b == r_count_45_io_out ? io_r_27_b : _GEN_4676; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4678 = 7'h1c == r_count_45_io_out ? io_r_28_b : _GEN_4677; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4679 = 7'h1d == r_count_45_io_out ? io_r_29_b : _GEN_4678; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4680 = 7'h1e == r_count_45_io_out ? io_r_30_b : _GEN_4679; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4681 = 7'h1f == r_count_45_io_out ? io_r_31_b : _GEN_4680; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4682 = 7'h20 == r_count_45_io_out ? io_r_32_b : _GEN_4681; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4683 = 7'h21 == r_count_45_io_out ? io_r_33_b : _GEN_4682; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4684 = 7'h22 == r_count_45_io_out ? io_r_34_b : _GEN_4683; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4685 = 7'h23 == r_count_45_io_out ? io_r_35_b : _GEN_4684; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4686 = 7'h24 == r_count_45_io_out ? io_r_36_b : _GEN_4685; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4687 = 7'h25 == r_count_45_io_out ? io_r_37_b : _GEN_4686; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4688 = 7'h26 == r_count_45_io_out ? io_r_38_b : _GEN_4687; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4689 = 7'h27 == r_count_45_io_out ? io_r_39_b : _GEN_4688; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4690 = 7'h28 == r_count_45_io_out ? io_r_40_b : _GEN_4689; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4691 = 7'h29 == r_count_45_io_out ? io_r_41_b : _GEN_4690; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4692 = 7'h2a == r_count_45_io_out ? io_r_42_b : _GEN_4691; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4693 = 7'h2b == r_count_45_io_out ? io_r_43_b : _GEN_4692; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4694 = 7'h2c == r_count_45_io_out ? io_r_44_b : _GEN_4693; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4695 = 7'h2d == r_count_45_io_out ? io_r_45_b : _GEN_4694; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4696 = 7'h2e == r_count_45_io_out ? io_r_46_b : _GEN_4695; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4697 = 7'h2f == r_count_45_io_out ? io_r_47_b : _GEN_4696; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4698 = 7'h30 == r_count_45_io_out ? io_r_48_b : _GEN_4697; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4699 = 7'h31 == r_count_45_io_out ? io_r_49_b : _GEN_4698; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4700 = 7'h32 == r_count_45_io_out ? io_r_50_b : _GEN_4699; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4701 = 7'h33 == r_count_45_io_out ? io_r_51_b : _GEN_4700; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4702 = 7'h34 == r_count_45_io_out ? io_r_52_b : _GEN_4701; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4703 = 7'h35 == r_count_45_io_out ? io_r_53_b : _GEN_4702; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4704 = 7'h36 == r_count_45_io_out ? io_r_54_b : _GEN_4703; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4705 = 7'h37 == r_count_45_io_out ? io_r_55_b : _GEN_4704; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4706 = 7'h38 == r_count_45_io_out ? io_r_56_b : _GEN_4705; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4707 = 7'h39 == r_count_45_io_out ? io_r_57_b : _GEN_4706; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4708 = 7'h3a == r_count_45_io_out ? io_r_58_b : _GEN_4707; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4709 = 7'h3b == r_count_45_io_out ? io_r_59_b : _GEN_4708; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4710 = 7'h3c == r_count_45_io_out ? io_r_60_b : _GEN_4709; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4711 = 7'h3d == r_count_45_io_out ? io_r_61_b : _GEN_4710; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4712 = 7'h3e == r_count_45_io_out ? io_r_62_b : _GEN_4711; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4713 = 7'h3f == r_count_45_io_out ? io_r_63_b : _GEN_4712; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4714 = 7'h40 == r_count_45_io_out ? io_r_64_b : _GEN_4713; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4715 = 7'h41 == r_count_45_io_out ? io_r_65_b : _GEN_4714; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4716 = 7'h42 == r_count_45_io_out ? io_r_66_b : _GEN_4715; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4717 = 7'h43 == r_count_45_io_out ? io_r_67_b : _GEN_4716; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4718 = 7'h44 == r_count_45_io_out ? io_r_68_b : _GEN_4717; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4719 = 7'h45 == r_count_45_io_out ? io_r_69_b : _GEN_4718; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4720 = 7'h46 == r_count_45_io_out ? io_r_70_b : _GEN_4719; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4721 = 7'h47 == r_count_45_io_out ? io_r_71_b : _GEN_4720; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4722 = 7'h48 == r_count_45_io_out ? io_r_72_b : _GEN_4721; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4723 = 7'h49 == r_count_45_io_out ? io_r_73_b : _GEN_4722; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4724 = 7'h4a == r_count_45_io_out ? io_r_74_b : _GEN_4723; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4725 = 7'h4b == r_count_45_io_out ? io_r_75_b : _GEN_4724; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4726 = 7'h4c == r_count_45_io_out ? io_r_76_b : _GEN_4725; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4727 = 7'h4d == r_count_45_io_out ? io_r_77_b : _GEN_4726; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4728 = 7'h4e == r_count_45_io_out ? io_r_78_b : _GEN_4727; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4729 = 7'h4f == r_count_45_io_out ? io_r_79_b : _GEN_4728; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4730 = 7'h50 == r_count_45_io_out ? io_r_80_b : _GEN_4729; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4731 = 7'h51 == r_count_45_io_out ? io_r_81_b : _GEN_4730; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4732 = 7'h52 == r_count_45_io_out ? io_r_82_b : _GEN_4731; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4733 = 7'h53 == r_count_45_io_out ? io_r_83_b : _GEN_4732; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4734 = 7'h54 == r_count_45_io_out ? io_r_84_b : _GEN_4733; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4735 = 7'h55 == r_count_45_io_out ? io_r_85_b : _GEN_4734; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4736 = 7'h56 == r_count_45_io_out ? io_r_86_b : _GEN_4735; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4737 = 7'h57 == r_count_45_io_out ? io_r_87_b : _GEN_4736; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4738 = 7'h58 == r_count_45_io_out ? io_r_88_b : _GEN_4737; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4739 = 7'h59 == r_count_45_io_out ? io_r_89_b : _GEN_4738; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4740 = 7'h5a == r_count_45_io_out ? io_r_90_b : _GEN_4739; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4741 = 7'h5b == r_count_45_io_out ? io_r_91_b : _GEN_4740; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4742 = 7'h5c == r_count_45_io_out ? io_r_92_b : _GEN_4741; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4743 = 7'h5d == r_count_45_io_out ? io_r_93_b : _GEN_4742; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4744 = 7'h5e == r_count_45_io_out ? io_r_94_b : _GEN_4743; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4745 = 7'h5f == r_count_45_io_out ? io_r_95_b : _GEN_4744; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4746 = 7'h60 == r_count_45_io_out ? io_r_96_b : _GEN_4745; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4747 = 7'h61 == r_count_45_io_out ? io_r_97_b : _GEN_4746; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4748 = 7'h62 == r_count_45_io_out ? io_r_98_b : _GEN_4747; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4751 = 7'h1 == r_count_46_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4752 = 7'h2 == r_count_46_io_out ? io_r_2_b : _GEN_4751; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4753 = 7'h3 == r_count_46_io_out ? io_r_3_b : _GEN_4752; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4754 = 7'h4 == r_count_46_io_out ? io_r_4_b : _GEN_4753; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4755 = 7'h5 == r_count_46_io_out ? io_r_5_b : _GEN_4754; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4756 = 7'h6 == r_count_46_io_out ? io_r_6_b : _GEN_4755; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4757 = 7'h7 == r_count_46_io_out ? io_r_7_b : _GEN_4756; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4758 = 7'h8 == r_count_46_io_out ? io_r_8_b : _GEN_4757; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4759 = 7'h9 == r_count_46_io_out ? io_r_9_b : _GEN_4758; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4760 = 7'ha == r_count_46_io_out ? io_r_10_b : _GEN_4759; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4761 = 7'hb == r_count_46_io_out ? io_r_11_b : _GEN_4760; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4762 = 7'hc == r_count_46_io_out ? io_r_12_b : _GEN_4761; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4763 = 7'hd == r_count_46_io_out ? io_r_13_b : _GEN_4762; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4764 = 7'he == r_count_46_io_out ? io_r_14_b : _GEN_4763; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4765 = 7'hf == r_count_46_io_out ? io_r_15_b : _GEN_4764; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4766 = 7'h10 == r_count_46_io_out ? io_r_16_b : _GEN_4765; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4767 = 7'h11 == r_count_46_io_out ? io_r_17_b : _GEN_4766; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4768 = 7'h12 == r_count_46_io_out ? io_r_18_b : _GEN_4767; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4769 = 7'h13 == r_count_46_io_out ? io_r_19_b : _GEN_4768; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4770 = 7'h14 == r_count_46_io_out ? io_r_20_b : _GEN_4769; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4771 = 7'h15 == r_count_46_io_out ? io_r_21_b : _GEN_4770; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4772 = 7'h16 == r_count_46_io_out ? io_r_22_b : _GEN_4771; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4773 = 7'h17 == r_count_46_io_out ? io_r_23_b : _GEN_4772; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4774 = 7'h18 == r_count_46_io_out ? io_r_24_b : _GEN_4773; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4775 = 7'h19 == r_count_46_io_out ? io_r_25_b : _GEN_4774; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4776 = 7'h1a == r_count_46_io_out ? io_r_26_b : _GEN_4775; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4777 = 7'h1b == r_count_46_io_out ? io_r_27_b : _GEN_4776; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4778 = 7'h1c == r_count_46_io_out ? io_r_28_b : _GEN_4777; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4779 = 7'h1d == r_count_46_io_out ? io_r_29_b : _GEN_4778; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4780 = 7'h1e == r_count_46_io_out ? io_r_30_b : _GEN_4779; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4781 = 7'h1f == r_count_46_io_out ? io_r_31_b : _GEN_4780; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4782 = 7'h20 == r_count_46_io_out ? io_r_32_b : _GEN_4781; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4783 = 7'h21 == r_count_46_io_out ? io_r_33_b : _GEN_4782; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4784 = 7'h22 == r_count_46_io_out ? io_r_34_b : _GEN_4783; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4785 = 7'h23 == r_count_46_io_out ? io_r_35_b : _GEN_4784; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4786 = 7'h24 == r_count_46_io_out ? io_r_36_b : _GEN_4785; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4787 = 7'h25 == r_count_46_io_out ? io_r_37_b : _GEN_4786; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4788 = 7'h26 == r_count_46_io_out ? io_r_38_b : _GEN_4787; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4789 = 7'h27 == r_count_46_io_out ? io_r_39_b : _GEN_4788; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4790 = 7'h28 == r_count_46_io_out ? io_r_40_b : _GEN_4789; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4791 = 7'h29 == r_count_46_io_out ? io_r_41_b : _GEN_4790; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4792 = 7'h2a == r_count_46_io_out ? io_r_42_b : _GEN_4791; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4793 = 7'h2b == r_count_46_io_out ? io_r_43_b : _GEN_4792; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4794 = 7'h2c == r_count_46_io_out ? io_r_44_b : _GEN_4793; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4795 = 7'h2d == r_count_46_io_out ? io_r_45_b : _GEN_4794; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4796 = 7'h2e == r_count_46_io_out ? io_r_46_b : _GEN_4795; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4797 = 7'h2f == r_count_46_io_out ? io_r_47_b : _GEN_4796; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4798 = 7'h30 == r_count_46_io_out ? io_r_48_b : _GEN_4797; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4799 = 7'h31 == r_count_46_io_out ? io_r_49_b : _GEN_4798; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4800 = 7'h32 == r_count_46_io_out ? io_r_50_b : _GEN_4799; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4801 = 7'h33 == r_count_46_io_out ? io_r_51_b : _GEN_4800; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4802 = 7'h34 == r_count_46_io_out ? io_r_52_b : _GEN_4801; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4803 = 7'h35 == r_count_46_io_out ? io_r_53_b : _GEN_4802; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4804 = 7'h36 == r_count_46_io_out ? io_r_54_b : _GEN_4803; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4805 = 7'h37 == r_count_46_io_out ? io_r_55_b : _GEN_4804; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4806 = 7'h38 == r_count_46_io_out ? io_r_56_b : _GEN_4805; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4807 = 7'h39 == r_count_46_io_out ? io_r_57_b : _GEN_4806; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4808 = 7'h3a == r_count_46_io_out ? io_r_58_b : _GEN_4807; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4809 = 7'h3b == r_count_46_io_out ? io_r_59_b : _GEN_4808; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4810 = 7'h3c == r_count_46_io_out ? io_r_60_b : _GEN_4809; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4811 = 7'h3d == r_count_46_io_out ? io_r_61_b : _GEN_4810; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4812 = 7'h3e == r_count_46_io_out ? io_r_62_b : _GEN_4811; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4813 = 7'h3f == r_count_46_io_out ? io_r_63_b : _GEN_4812; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4814 = 7'h40 == r_count_46_io_out ? io_r_64_b : _GEN_4813; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4815 = 7'h41 == r_count_46_io_out ? io_r_65_b : _GEN_4814; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4816 = 7'h42 == r_count_46_io_out ? io_r_66_b : _GEN_4815; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4817 = 7'h43 == r_count_46_io_out ? io_r_67_b : _GEN_4816; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4818 = 7'h44 == r_count_46_io_out ? io_r_68_b : _GEN_4817; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4819 = 7'h45 == r_count_46_io_out ? io_r_69_b : _GEN_4818; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4820 = 7'h46 == r_count_46_io_out ? io_r_70_b : _GEN_4819; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4821 = 7'h47 == r_count_46_io_out ? io_r_71_b : _GEN_4820; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4822 = 7'h48 == r_count_46_io_out ? io_r_72_b : _GEN_4821; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4823 = 7'h49 == r_count_46_io_out ? io_r_73_b : _GEN_4822; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4824 = 7'h4a == r_count_46_io_out ? io_r_74_b : _GEN_4823; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4825 = 7'h4b == r_count_46_io_out ? io_r_75_b : _GEN_4824; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4826 = 7'h4c == r_count_46_io_out ? io_r_76_b : _GEN_4825; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4827 = 7'h4d == r_count_46_io_out ? io_r_77_b : _GEN_4826; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4828 = 7'h4e == r_count_46_io_out ? io_r_78_b : _GEN_4827; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4829 = 7'h4f == r_count_46_io_out ? io_r_79_b : _GEN_4828; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4830 = 7'h50 == r_count_46_io_out ? io_r_80_b : _GEN_4829; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4831 = 7'h51 == r_count_46_io_out ? io_r_81_b : _GEN_4830; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4832 = 7'h52 == r_count_46_io_out ? io_r_82_b : _GEN_4831; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4833 = 7'h53 == r_count_46_io_out ? io_r_83_b : _GEN_4832; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4834 = 7'h54 == r_count_46_io_out ? io_r_84_b : _GEN_4833; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4835 = 7'h55 == r_count_46_io_out ? io_r_85_b : _GEN_4834; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4836 = 7'h56 == r_count_46_io_out ? io_r_86_b : _GEN_4835; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4837 = 7'h57 == r_count_46_io_out ? io_r_87_b : _GEN_4836; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4838 = 7'h58 == r_count_46_io_out ? io_r_88_b : _GEN_4837; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4839 = 7'h59 == r_count_46_io_out ? io_r_89_b : _GEN_4838; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4840 = 7'h5a == r_count_46_io_out ? io_r_90_b : _GEN_4839; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4841 = 7'h5b == r_count_46_io_out ? io_r_91_b : _GEN_4840; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4842 = 7'h5c == r_count_46_io_out ? io_r_92_b : _GEN_4841; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4843 = 7'h5d == r_count_46_io_out ? io_r_93_b : _GEN_4842; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4844 = 7'h5e == r_count_46_io_out ? io_r_94_b : _GEN_4843; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4845 = 7'h5f == r_count_46_io_out ? io_r_95_b : _GEN_4844; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4846 = 7'h60 == r_count_46_io_out ? io_r_96_b : _GEN_4845; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4847 = 7'h61 == r_count_46_io_out ? io_r_97_b : _GEN_4846; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4848 = 7'h62 == r_count_46_io_out ? io_r_98_b : _GEN_4847; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4851 = 7'h1 == r_count_47_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4852 = 7'h2 == r_count_47_io_out ? io_r_2_b : _GEN_4851; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4853 = 7'h3 == r_count_47_io_out ? io_r_3_b : _GEN_4852; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4854 = 7'h4 == r_count_47_io_out ? io_r_4_b : _GEN_4853; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4855 = 7'h5 == r_count_47_io_out ? io_r_5_b : _GEN_4854; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4856 = 7'h6 == r_count_47_io_out ? io_r_6_b : _GEN_4855; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4857 = 7'h7 == r_count_47_io_out ? io_r_7_b : _GEN_4856; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4858 = 7'h8 == r_count_47_io_out ? io_r_8_b : _GEN_4857; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4859 = 7'h9 == r_count_47_io_out ? io_r_9_b : _GEN_4858; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4860 = 7'ha == r_count_47_io_out ? io_r_10_b : _GEN_4859; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4861 = 7'hb == r_count_47_io_out ? io_r_11_b : _GEN_4860; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4862 = 7'hc == r_count_47_io_out ? io_r_12_b : _GEN_4861; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4863 = 7'hd == r_count_47_io_out ? io_r_13_b : _GEN_4862; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4864 = 7'he == r_count_47_io_out ? io_r_14_b : _GEN_4863; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4865 = 7'hf == r_count_47_io_out ? io_r_15_b : _GEN_4864; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4866 = 7'h10 == r_count_47_io_out ? io_r_16_b : _GEN_4865; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4867 = 7'h11 == r_count_47_io_out ? io_r_17_b : _GEN_4866; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4868 = 7'h12 == r_count_47_io_out ? io_r_18_b : _GEN_4867; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4869 = 7'h13 == r_count_47_io_out ? io_r_19_b : _GEN_4868; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4870 = 7'h14 == r_count_47_io_out ? io_r_20_b : _GEN_4869; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4871 = 7'h15 == r_count_47_io_out ? io_r_21_b : _GEN_4870; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4872 = 7'h16 == r_count_47_io_out ? io_r_22_b : _GEN_4871; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4873 = 7'h17 == r_count_47_io_out ? io_r_23_b : _GEN_4872; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4874 = 7'h18 == r_count_47_io_out ? io_r_24_b : _GEN_4873; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4875 = 7'h19 == r_count_47_io_out ? io_r_25_b : _GEN_4874; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4876 = 7'h1a == r_count_47_io_out ? io_r_26_b : _GEN_4875; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4877 = 7'h1b == r_count_47_io_out ? io_r_27_b : _GEN_4876; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4878 = 7'h1c == r_count_47_io_out ? io_r_28_b : _GEN_4877; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4879 = 7'h1d == r_count_47_io_out ? io_r_29_b : _GEN_4878; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4880 = 7'h1e == r_count_47_io_out ? io_r_30_b : _GEN_4879; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4881 = 7'h1f == r_count_47_io_out ? io_r_31_b : _GEN_4880; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4882 = 7'h20 == r_count_47_io_out ? io_r_32_b : _GEN_4881; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4883 = 7'h21 == r_count_47_io_out ? io_r_33_b : _GEN_4882; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4884 = 7'h22 == r_count_47_io_out ? io_r_34_b : _GEN_4883; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4885 = 7'h23 == r_count_47_io_out ? io_r_35_b : _GEN_4884; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4886 = 7'h24 == r_count_47_io_out ? io_r_36_b : _GEN_4885; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4887 = 7'h25 == r_count_47_io_out ? io_r_37_b : _GEN_4886; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4888 = 7'h26 == r_count_47_io_out ? io_r_38_b : _GEN_4887; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4889 = 7'h27 == r_count_47_io_out ? io_r_39_b : _GEN_4888; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4890 = 7'h28 == r_count_47_io_out ? io_r_40_b : _GEN_4889; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4891 = 7'h29 == r_count_47_io_out ? io_r_41_b : _GEN_4890; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4892 = 7'h2a == r_count_47_io_out ? io_r_42_b : _GEN_4891; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4893 = 7'h2b == r_count_47_io_out ? io_r_43_b : _GEN_4892; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4894 = 7'h2c == r_count_47_io_out ? io_r_44_b : _GEN_4893; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4895 = 7'h2d == r_count_47_io_out ? io_r_45_b : _GEN_4894; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4896 = 7'h2e == r_count_47_io_out ? io_r_46_b : _GEN_4895; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4897 = 7'h2f == r_count_47_io_out ? io_r_47_b : _GEN_4896; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4898 = 7'h30 == r_count_47_io_out ? io_r_48_b : _GEN_4897; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4899 = 7'h31 == r_count_47_io_out ? io_r_49_b : _GEN_4898; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4900 = 7'h32 == r_count_47_io_out ? io_r_50_b : _GEN_4899; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4901 = 7'h33 == r_count_47_io_out ? io_r_51_b : _GEN_4900; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4902 = 7'h34 == r_count_47_io_out ? io_r_52_b : _GEN_4901; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4903 = 7'h35 == r_count_47_io_out ? io_r_53_b : _GEN_4902; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4904 = 7'h36 == r_count_47_io_out ? io_r_54_b : _GEN_4903; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4905 = 7'h37 == r_count_47_io_out ? io_r_55_b : _GEN_4904; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4906 = 7'h38 == r_count_47_io_out ? io_r_56_b : _GEN_4905; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4907 = 7'h39 == r_count_47_io_out ? io_r_57_b : _GEN_4906; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4908 = 7'h3a == r_count_47_io_out ? io_r_58_b : _GEN_4907; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4909 = 7'h3b == r_count_47_io_out ? io_r_59_b : _GEN_4908; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4910 = 7'h3c == r_count_47_io_out ? io_r_60_b : _GEN_4909; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4911 = 7'h3d == r_count_47_io_out ? io_r_61_b : _GEN_4910; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4912 = 7'h3e == r_count_47_io_out ? io_r_62_b : _GEN_4911; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4913 = 7'h3f == r_count_47_io_out ? io_r_63_b : _GEN_4912; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4914 = 7'h40 == r_count_47_io_out ? io_r_64_b : _GEN_4913; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4915 = 7'h41 == r_count_47_io_out ? io_r_65_b : _GEN_4914; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4916 = 7'h42 == r_count_47_io_out ? io_r_66_b : _GEN_4915; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4917 = 7'h43 == r_count_47_io_out ? io_r_67_b : _GEN_4916; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4918 = 7'h44 == r_count_47_io_out ? io_r_68_b : _GEN_4917; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4919 = 7'h45 == r_count_47_io_out ? io_r_69_b : _GEN_4918; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4920 = 7'h46 == r_count_47_io_out ? io_r_70_b : _GEN_4919; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4921 = 7'h47 == r_count_47_io_out ? io_r_71_b : _GEN_4920; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4922 = 7'h48 == r_count_47_io_out ? io_r_72_b : _GEN_4921; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4923 = 7'h49 == r_count_47_io_out ? io_r_73_b : _GEN_4922; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4924 = 7'h4a == r_count_47_io_out ? io_r_74_b : _GEN_4923; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4925 = 7'h4b == r_count_47_io_out ? io_r_75_b : _GEN_4924; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4926 = 7'h4c == r_count_47_io_out ? io_r_76_b : _GEN_4925; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4927 = 7'h4d == r_count_47_io_out ? io_r_77_b : _GEN_4926; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4928 = 7'h4e == r_count_47_io_out ? io_r_78_b : _GEN_4927; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4929 = 7'h4f == r_count_47_io_out ? io_r_79_b : _GEN_4928; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4930 = 7'h50 == r_count_47_io_out ? io_r_80_b : _GEN_4929; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4931 = 7'h51 == r_count_47_io_out ? io_r_81_b : _GEN_4930; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4932 = 7'h52 == r_count_47_io_out ? io_r_82_b : _GEN_4931; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4933 = 7'h53 == r_count_47_io_out ? io_r_83_b : _GEN_4932; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4934 = 7'h54 == r_count_47_io_out ? io_r_84_b : _GEN_4933; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4935 = 7'h55 == r_count_47_io_out ? io_r_85_b : _GEN_4934; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4936 = 7'h56 == r_count_47_io_out ? io_r_86_b : _GEN_4935; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4937 = 7'h57 == r_count_47_io_out ? io_r_87_b : _GEN_4936; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4938 = 7'h58 == r_count_47_io_out ? io_r_88_b : _GEN_4937; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4939 = 7'h59 == r_count_47_io_out ? io_r_89_b : _GEN_4938; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4940 = 7'h5a == r_count_47_io_out ? io_r_90_b : _GEN_4939; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4941 = 7'h5b == r_count_47_io_out ? io_r_91_b : _GEN_4940; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4942 = 7'h5c == r_count_47_io_out ? io_r_92_b : _GEN_4941; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4943 = 7'h5d == r_count_47_io_out ? io_r_93_b : _GEN_4942; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4944 = 7'h5e == r_count_47_io_out ? io_r_94_b : _GEN_4943; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4945 = 7'h5f == r_count_47_io_out ? io_r_95_b : _GEN_4944; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4946 = 7'h60 == r_count_47_io_out ? io_r_96_b : _GEN_4945; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4947 = 7'h61 == r_count_47_io_out ? io_r_97_b : _GEN_4946; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4948 = 7'h62 == r_count_47_io_out ? io_r_98_b : _GEN_4947; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4951 = 7'h1 == r_count_48_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4952 = 7'h2 == r_count_48_io_out ? io_r_2_b : _GEN_4951; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4953 = 7'h3 == r_count_48_io_out ? io_r_3_b : _GEN_4952; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4954 = 7'h4 == r_count_48_io_out ? io_r_4_b : _GEN_4953; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4955 = 7'h5 == r_count_48_io_out ? io_r_5_b : _GEN_4954; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4956 = 7'h6 == r_count_48_io_out ? io_r_6_b : _GEN_4955; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4957 = 7'h7 == r_count_48_io_out ? io_r_7_b : _GEN_4956; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4958 = 7'h8 == r_count_48_io_out ? io_r_8_b : _GEN_4957; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4959 = 7'h9 == r_count_48_io_out ? io_r_9_b : _GEN_4958; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4960 = 7'ha == r_count_48_io_out ? io_r_10_b : _GEN_4959; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4961 = 7'hb == r_count_48_io_out ? io_r_11_b : _GEN_4960; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4962 = 7'hc == r_count_48_io_out ? io_r_12_b : _GEN_4961; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4963 = 7'hd == r_count_48_io_out ? io_r_13_b : _GEN_4962; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4964 = 7'he == r_count_48_io_out ? io_r_14_b : _GEN_4963; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4965 = 7'hf == r_count_48_io_out ? io_r_15_b : _GEN_4964; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4966 = 7'h10 == r_count_48_io_out ? io_r_16_b : _GEN_4965; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4967 = 7'h11 == r_count_48_io_out ? io_r_17_b : _GEN_4966; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4968 = 7'h12 == r_count_48_io_out ? io_r_18_b : _GEN_4967; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4969 = 7'h13 == r_count_48_io_out ? io_r_19_b : _GEN_4968; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4970 = 7'h14 == r_count_48_io_out ? io_r_20_b : _GEN_4969; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4971 = 7'h15 == r_count_48_io_out ? io_r_21_b : _GEN_4970; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4972 = 7'h16 == r_count_48_io_out ? io_r_22_b : _GEN_4971; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4973 = 7'h17 == r_count_48_io_out ? io_r_23_b : _GEN_4972; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4974 = 7'h18 == r_count_48_io_out ? io_r_24_b : _GEN_4973; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4975 = 7'h19 == r_count_48_io_out ? io_r_25_b : _GEN_4974; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4976 = 7'h1a == r_count_48_io_out ? io_r_26_b : _GEN_4975; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4977 = 7'h1b == r_count_48_io_out ? io_r_27_b : _GEN_4976; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4978 = 7'h1c == r_count_48_io_out ? io_r_28_b : _GEN_4977; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4979 = 7'h1d == r_count_48_io_out ? io_r_29_b : _GEN_4978; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4980 = 7'h1e == r_count_48_io_out ? io_r_30_b : _GEN_4979; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4981 = 7'h1f == r_count_48_io_out ? io_r_31_b : _GEN_4980; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4982 = 7'h20 == r_count_48_io_out ? io_r_32_b : _GEN_4981; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4983 = 7'h21 == r_count_48_io_out ? io_r_33_b : _GEN_4982; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4984 = 7'h22 == r_count_48_io_out ? io_r_34_b : _GEN_4983; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4985 = 7'h23 == r_count_48_io_out ? io_r_35_b : _GEN_4984; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4986 = 7'h24 == r_count_48_io_out ? io_r_36_b : _GEN_4985; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4987 = 7'h25 == r_count_48_io_out ? io_r_37_b : _GEN_4986; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4988 = 7'h26 == r_count_48_io_out ? io_r_38_b : _GEN_4987; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4989 = 7'h27 == r_count_48_io_out ? io_r_39_b : _GEN_4988; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4990 = 7'h28 == r_count_48_io_out ? io_r_40_b : _GEN_4989; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4991 = 7'h29 == r_count_48_io_out ? io_r_41_b : _GEN_4990; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4992 = 7'h2a == r_count_48_io_out ? io_r_42_b : _GEN_4991; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4993 = 7'h2b == r_count_48_io_out ? io_r_43_b : _GEN_4992; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4994 = 7'h2c == r_count_48_io_out ? io_r_44_b : _GEN_4993; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4995 = 7'h2d == r_count_48_io_out ? io_r_45_b : _GEN_4994; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4996 = 7'h2e == r_count_48_io_out ? io_r_46_b : _GEN_4995; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4997 = 7'h2f == r_count_48_io_out ? io_r_47_b : _GEN_4996; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4998 = 7'h30 == r_count_48_io_out ? io_r_48_b : _GEN_4997; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_4999 = 7'h31 == r_count_48_io_out ? io_r_49_b : _GEN_4998; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5000 = 7'h32 == r_count_48_io_out ? io_r_50_b : _GEN_4999; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5001 = 7'h33 == r_count_48_io_out ? io_r_51_b : _GEN_5000; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5002 = 7'h34 == r_count_48_io_out ? io_r_52_b : _GEN_5001; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5003 = 7'h35 == r_count_48_io_out ? io_r_53_b : _GEN_5002; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5004 = 7'h36 == r_count_48_io_out ? io_r_54_b : _GEN_5003; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5005 = 7'h37 == r_count_48_io_out ? io_r_55_b : _GEN_5004; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5006 = 7'h38 == r_count_48_io_out ? io_r_56_b : _GEN_5005; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5007 = 7'h39 == r_count_48_io_out ? io_r_57_b : _GEN_5006; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5008 = 7'h3a == r_count_48_io_out ? io_r_58_b : _GEN_5007; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5009 = 7'h3b == r_count_48_io_out ? io_r_59_b : _GEN_5008; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5010 = 7'h3c == r_count_48_io_out ? io_r_60_b : _GEN_5009; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5011 = 7'h3d == r_count_48_io_out ? io_r_61_b : _GEN_5010; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5012 = 7'h3e == r_count_48_io_out ? io_r_62_b : _GEN_5011; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5013 = 7'h3f == r_count_48_io_out ? io_r_63_b : _GEN_5012; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5014 = 7'h40 == r_count_48_io_out ? io_r_64_b : _GEN_5013; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5015 = 7'h41 == r_count_48_io_out ? io_r_65_b : _GEN_5014; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5016 = 7'h42 == r_count_48_io_out ? io_r_66_b : _GEN_5015; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5017 = 7'h43 == r_count_48_io_out ? io_r_67_b : _GEN_5016; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5018 = 7'h44 == r_count_48_io_out ? io_r_68_b : _GEN_5017; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5019 = 7'h45 == r_count_48_io_out ? io_r_69_b : _GEN_5018; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5020 = 7'h46 == r_count_48_io_out ? io_r_70_b : _GEN_5019; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5021 = 7'h47 == r_count_48_io_out ? io_r_71_b : _GEN_5020; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5022 = 7'h48 == r_count_48_io_out ? io_r_72_b : _GEN_5021; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5023 = 7'h49 == r_count_48_io_out ? io_r_73_b : _GEN_5022; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5024 = 7'h4a == r_count_48_io_out ? io_r_74_b : _GEN_5023; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5025 = 7'h4b == r_count_48_io_out ? io_r_75_b : _GEN_5024; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5026 = 7'h4c == r_count_48_io_out ? io_r_76_b : _GEN_5025; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5027 = 7'h4d == r_count_48_io_out ? io_r_77_b : _GEN_5026; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5028 = 7'h4e == r_count_48_io_out ? io_r_78_b : _GEN_5027; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5029 = 7'h4f == r_count_48_io_out ? io_r_79_b : _GEN_5028; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5030 = 7'h50 == r_count_48_io_out ? io_r_80_b : _GEN_5029; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5031 = 7'h51 == r_count_48_io_out ? io_r_81_b : _GEN_5030; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5032 = 7'h52 == r_count_48_io_out ? io_r_82_b : _GEN_5031; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5033 = 7'h53 == r_count_48_io_out ? io_r_83_b : _GEN_5032; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5034 = 7'h54 == r_count_48_io_out ? io_r_84_b : _GEN_5033; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5035 = 7'h55 == r_count_48_io_out ? io_r_85_b : _GEN_5034; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5036 = 7'h56 == r_count_48_io_out ? io_r_86_b : _GEN_5035; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5037 = 7'h57 == r_count_48_io_out ? io_r_87_b : _GEN_5036; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5038 = 7'h58 == r_count_48_io_out ? io_r_88_b : _GEN_5037; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5039 = 7'h59 == r_count_48_io_out ? io_r_89_b : _GEN_5038; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5040 = 7'h5a == r_count_48_io_out ? io_r_90_b : _GEN_5039; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5041 = 7'h5b == r_count_48_io_out ? io_r_91_b : _GEN_5040; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5042 = 7'h5c == r_count_48_io_out ? io_r_92_b : _GEN_5041; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5043 = 7'h5d == r_count_48_io_out ? io_r_93_b : _GEN_5042; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5044 = 7'h5e == r_count_48_io_out ? io_r_94_b : _GEN_5043; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5045 = 7'h5f == r_count_48_io_out ? io_r_95_b : _GEN_5044; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5046 = 7'h60 == r_count_48_io_out ? io_r_96_b : _GEN_5045; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5047 = 7'h61 == r_count_48_io_out ? io_r_97_b : _GEN_5046; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5048 = 7'h62 == r_count_48_io_out ? io_r_98_b : _GEN_5047; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5051 = 7'h1 == r_count_49_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5052 = 7'h2 == r_count_49_io_out ? io_r_2_b : _GEN_5051; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5053 = 7'h3 == r_count_49_io_out ? io_r_3_b : _GEN_5052; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5054 = 7'h4 == r_count_49_io_out ? io_r_4_b : _GEN_5053; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5055 = 7'h5 == r_count_49_io_out ? io_r_5_b : _GEN_5054; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5056 = 7'h6 == r_count_49_io_out ? io_r_6_b : _GEN_5055; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5057 = 7'h7 == r_count_49_io_out ? io_r_7_b : _GEN_5056; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5058 = 7'h8 == r_count_49_io_out ? io_r_8_b : _GEN_5057; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5059 = 7'h9 == r_count_49_io_out ? io_r_9_b : _GEN_5058; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5060 = 7'ha == r_count_49_io_out ? io_r_10_b : _GEN_5059; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5061 = 7'hb == r_count_49_io_out ? io_r_11_b : _GEN_5060; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5062 = 7'hc == r_count_49_io_out ? io_r_12_b : _GEN_5061; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5063 = 7'hd == r_count_49_io_out ? io_r_13_b : _GEN_5062; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5064 = 7'he == r_count_49_io_out ? io_r_14_b : _GEN_5063; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5065 = 7'hf == r_count_49_io_out ? io_r_15_b : _GEN_5064; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5066 = 7'h10 == r_count_49_io_out ? io_r_16_b : _GEN_5065; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5067 = 7'h11 == r_count_49_io_out ? io_r_17_b : _GEN_5066; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5068 = 7'h12 == r_count_49_io_out ? io_r_18_b : _GEN_5067; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5069 = 7'h13 == r_count_49_io_out ? io_r_19_b : _GEN_5068; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5070 = 7'h14 == r_count_49_io_out ? io_r_20_b : _GEN_5069; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5071 = 7'h15 == r_count_49_io_out ? io_r_21_b : _GEN_5070; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5072 = 7'h16 == r_count_49_io_out ? io_r_22_b : _GEN_5071; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5073 = 7'h17 == r_count_49_io_out ? io_r_23_b : _GEN_5072; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5074 = 7'h18 == r_count_49_io_out ? io_r_24_b : _GEN_5073; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5075 = 7'h19 == r_count_49_io_out ? io_r_25_b : _GEN_5074; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5076 = 7'h1a == r_count_49_io_out ? io_r_26_b : _GEN_5075; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5077 = 7'h1b == r_count_49_io_out ? io_r_27_b : _GEN_5076; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5078 = 7'h1c == r_count_49_io_out ? io_r_28_b : _GEN_5077; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5079 = 7'h1d == r_count_49_io_out ? io_r_29_b : _GEN_5078; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5080 = 7'h1e == r_count_49_io_out ? io_r_30_b : _GEN_5079; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5081 = 7'h1f == r_count_49_io_out ? io_r_31_b : _GEN_5080; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5082 = 7'h20 == r_count_49_io_out ? io_r_32_b : _GEN_5081; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5083 = 7'h21 == r_count_49_io_out ? io_r_33_b : _GEN_5082; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5084 = 7'h22 == r_count_49_io_out ? io_r_34_b : _GEN_5083; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5085 = 7'h23 == r_count_49_io_out ? io_r_35_b : _GEN_5084; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5086 = 7'h24 == r_count_49_io_out ? io_r_36_b : _GEN_5085; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5087 = 7'h25 == r_count_49_io_out ? io_r_37_b : _GEN_5086; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5088 = 7'h26 == r_count_49_io_out ? io_r_38_b : _GEN_5087; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5089 = 7'h27 == r_count_49_io_out ? io_r_39_b : _GEN_5088; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5090 = 7'h28 == r_count_49_io_out ? io_r_40_b : _GEN_5089; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5091 = 7'h29 == r_count_49_io_out ? io_r_41_b : _GEN_5090; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5092 = 7'h2a == r_count_49_io_out ? io_r_42_b : _GEN_5091; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5093 = 7'h2b == r_count_49_io_out ? io_r_43_b : _GEN_5092; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5094 = 7'h2c == r_count_49_io_out ? io_r_44_b : _GEN_5093; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5095 = 7'h2d == r_count_49_io_out ? io_r_45_b : _GEN_5094; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5096 = 7'h2e == r_count_49_io_out ? io_r_46_b : _GEN_5095; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5097 = 7'h2f == r_count_49_io_out ? io_r_47_b : _GEN_5096; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5098 = 7'h30 == r_count_49_io_out ? io_r_48_b : _GEN_5097; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5099 = 7'h31 == r_count_49_io_out ? io_r_49_b : _GEN_5098; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5100 = 7'h32 == r_count_49_io_out ? io_r_50_b : _GEN_5099; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5101 = 7'h33 == r_count_49_io_out ? io_r_51_b : _GEN_5100; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5102 = 7'h34 == r_count_49_io_out ? io_r_52_b : _GEN_5101; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5103 = 7'h35 == r_count_49_io_out ? io_r_53_b : _GEN_5102; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5104 = 7'h36 == r_count_49_io_out ? io_r_54_b : _GEN_5103; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5105 = 7'h37 == r_count_49_io_out ? io_r_55_b : _GEN_5104; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5106 = 7'h38 == r_count_49_io_out ? io_r_56_b : _GEN_5105; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5107 = 7'h39 == r_count_49_io_out ? io_r_57_b : _GEN_5106; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5108 = 7'h3a == r_count_49_io_out ? io_r_58_b : _GEN_5107; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5109 = 7'h3b == r_count_49_io_out ? io_r_59_b : _GEN_5108; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5110 = 7'h3c == r_count_49_io_out ? io_r_60_b : _GEN_5109; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5111 = 7'h3d == r_count_49_io_out ? io_r_61_b : _GEN_5110; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5112 = 7'h3e == r_count_49_io_out ? io_r_62_b : _GEN_5111; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5113 = 7'h3f == r_count_49_io_out ? io_r_63_b : _GEN_5112; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5114 = 7'h40 == r_count_49_io_out ? io_r_64_b : _GEN_5113; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5115 = 7'h41 == r_count_49_io_out ? io_r_65_b : _GEN_5114; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5116 = 7'h42 == r_count_49_io_out ? io_r_66_b : _GEN_5115; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5117 = 7'h43 == r_count_49_io_out ? io_r_67_b : _GEN_5116; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5118 = 7'h44 == r_count_49_io_out ? io_r_68_b : _GEN_5117; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5119 = 7'h45 == r_count_49_io_out ? io_r_69_b : _GEN_5118; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5120 = 7'h46 == r_count_49_io_out ? io_r_70_b : _GEN_5119; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5121 = 7'h47 == r_count_49_io_out ? io_r_71_b : _GEN_5120; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5122 = 7'h48 == r_count_49_io_out ? io_r_72_b : _GEN_5121; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5123 = 7'h49 == r_count_49_io_out ? io_r_73_b : _GEN_5122; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5124 = 7'h4a == r_count_49_io_out ? io_r_74_b : _GEN_5123; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5125 = 7'h4b == r_count_49_io_out ? io_r_75_b : _GEN_5124; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5126 = 7'h4c == r_count_49_io_out ? io_r_76_b : _GEN_5125; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5127 = 7'h4d == r_count_49_io_out ? io_r_77_b : _GEN_5126; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5128 = 7'h4e == r_count_49_io_out ? io_r_78_b : _GEN_5127; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5129 = 7'h4f == r_count_49_io_out ? io_r_79_b : _GEN_5128; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5130 = 7'h50 == r_count_49_io_out ? io_r_80_b : _GEN_5129; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5131 = 7'h51 == r_count_49_io_out ? io_r_81_b : _GEN_5130; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5132 = 7'h52 == r_count_49_io_out ? io_r_82_b : _GEN_5131; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5133 = 7'h53 == r_count_49_io_out ? io_r_83_b : _GEN_5132; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5134 = 7'h54 == r_count_49_io_out ? io_r_84_b : _GEN_5133; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5135 = 7'h55 == r_count_49_io_out ? io_r_85_b : _GEN_5134; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5136 = 7'h56 == r_count_49_io_out ? io_r_86_b : _GEN_5135; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5137 = 7'h57 == r_count_49_io_out ? io_r_87_b : _GEN_5136; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5138 = 7'h58 == r_count_49_io_out ? io_r_88_b : _GEN_5137; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5139 = 7'h59 == r_count_49_io_out ? io_r_89_b : _GEN_5138; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5140 = 7'h5a == r_count_49_io_out ? io_r_90_b : _GEN_5139; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5141 = 7'h5b == r_count_49_io_out ? io_r_91_b : _GEN_5140; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5142 = 7'h5c == r_count_49_io_out ? io_r_92_b : _GEN_5141; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5143 = 7'h5d == r_count_49_io_out ? io_r_93_b : _GEN_5142; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5144 = 7'h5e == r_count_49_io_out ? io_r_94_b : _GEN_5143; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5145 = 7'h5f == r_count_49_io_out ? io_r_95_b : _GEN_5144; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5146 = 7'h60 == r_count_49_io_out ? io_r_96_b : _GEN_5145; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5147 = 7'h61 == r_count_49_io_out ? io_r_97_b : _GEN_5146; // @[SWChisel.scala 221:{19,19}]
  wire [1:0] _GEN_5148 = 7'h62 == r_count_49_io_out ? io_r_98_b : _GEN_5147; // @[SWChisel.scala 221:{19,19}]
  SWCell array_0 ( // @[SWChisel.scala 170:39]
    .io_q(array_0_io_q),
    .io_r(array_0_io_r),
    .io_e_i(array_0_io_e_i),
    .io_f_i(array_0_io_f_i),
    .io_ve_i(array_0_io_ve_i),
    .io_vf_i(array_0_io_vf_i),
    .io_vv_i(array_0_io_vv_i),
    .io_e_o(array_0_io_e_o),
    .io_f_o(array_0_io_f_o),
    .io_v_o(array_0_io_v_o)
  );
  SWCell array_1 ( // @[SWChisel.scala 170:39]
    .io_q(array_1_io_q),
    .io_r(array_1_io_r),
    .io_e_i(array_1_io_e_i),
    .io_f_i(array_1_io_f_i),
    .io_ve_i(array_1_io_ve_i),
    .io_vf_i(array_1_io_vf_i),
    .io_vv_i(array_1_io_vv_i),
    .io_e_o(array_1_io_e_o),
    .io_f_o(array_1_io_f_o),
    .io_v_o(array_1_io_v_o)
  );
  SWCell array_2 ( // @[SWChisel.scala 170:39]
    .io_q(array_2_io_q),
    .io_r(array_2_io_r),
    .io_e_i(array_2_io_e_i),
    .io_f_i(array_2_io_f_i),
    .io_ve_i(array_2_io_ve_i),
    .io_vf_i(array_2_io_vf_i),
    .io_vv_i(array_2_io_vv_i),
    .io_e_o(array_2_io_e_o),
    .io_f_o(array_2_io_f_o),
    .io_v_o(array_2_io_v_o)
  );
  SWCell array_3 ( // @[SWChisel.scala 170:39]
    .io_q(array_3_io_q),
    .io_r(array_3_io_r),
    .io_e_i(array_3_io_e_i),
    .io_f_i(array_3_io_f_i),
    .io_ve_i(array_3_io_ve_i),
    .io_vf_i(array_3_io_vf_i),
    .io_vv_i(array_3_io_vv_i),
    .io_e_o(array_3_io_e_o),
    .io_f_o(array_3_io_f_o),
    .io_v_o(array_3_io_v_o)
  );
  SWCell array_4 ( // @[SWChisel.scala 170:39]
    .io_q(array_4_io_q),
    .io_r(array_4_io_r),
    .io_e_i(array_4_io_e_i),
    .io_f_i(array_4_io_f_i),
    .io_ve_i(array_4_io_ve_i),
    .io_vf_i(array_4_io_vf_i),
    .io_vv_i(array_4_io_vv_i),
    .io_e_o(array_4_io_e_o),
    .io_f_o(array_4_io_f_o),
    .io_v_o(array_4_io_v_o)
  );
  SWCell array_5 ( // @[SWChisel.scala 170:39]
    .io_q(array_5_io_q),
    .io_r(array_5_io_r),
    .io_e_i(array_5_io_e_i),
    .io_f_i(array_5_io_f_i),
    .io_ve_i(array_5_io_ve_i),
    .io_vf_i(array_5_io_vf_i),
    .io_vv_i(array_5_io_vv_i),
    .io_e_o(array_5_io_e_o),
    .io_f_o(array_5_io_f_o),
    .io_v_o(array_5_io_v_o)
  );
  SWCell array_6 ( // @[SWChisel.scala 170:39]
    .io_q(array_6_io_q),
    .io_r(array_6_io_r),
    .io_e_i(array_6_io_e_i),
    .io_f_i(array_6_io_f_i),
    .io_ve_i(array_6_io_ve_i),
    .io_vf_i(array_6_io_vf_i),
    .io_vv_i(array_6_io_vv_i),
    .io_e_o(array_6_io_e_o),
    .io_f_o(array_6_io_f_o),
    .io_v_o(array_6_io_v_o)
  );
  SWCell array_7 ( // @[SWChisel.scala 170:39]
    .io_q(array_7_io_q),
    .io_r(array_7_io_r),
    .io_e_i(array_7_io_e_i),
    .io_f_i(array_7_io_f_i),
    .io_ve_i(array_7_io_ve_i),
    .io_vf_i(array_7_io_vf_i),
    .io_vv_i(array_7_io_vv_i),
    .io_e_o(array_7_io_e_o),
    .io_f_o(array_7_io_f_o),
    .io_v_o(array_7_io_v_o)
  );
  SWCell array_8 ( // @[SWChisel.scala 170:39]
    .io_q(array_8_io_q),
    .io_r(array_8_io_r),
    .io_e_i(array_8_io_e_i),
    .io_f_i(array_8_io_f_i),
    .io_ve_i(array_8_io_ve_i),
    .io_vf_i(array_8_io_vf_i),
    .io_vv_i(array_8_io_vv_i),
    .io_e_o(array_8_io_e_o),
    .io_f_o(array_8_io_f_o),
    .io_v_o(array_8_io_v_o)
  );
  SWCell array_9 ( // @[SWChisel.scala 170:39]
    .io_q(array_9_io_q),
    .io_r(array_9_io_r),
    .io_e_i(array_9_io_e_i),
    .io_f_i(array_9_io_f_i),
    .io_ve_i(array_9_io_ve_i),
    .io_vf_i(array_9_io_vf_i),
    .io_vv_i(array_9_io_vv_i),
    .io_e_o(array_9_io_e_o),
    .io_f_o(array_9_io_f_o),
    .io_v_o(array_9_io_v_o)
  );
  SWCell array_10 ( // @[SWChisel.scala 170:39]
    .io_q(array_10_io_q),
    .io_r(array_10_io_r),
    .io_e_i(array_10_io_e_i),
    .io_f_i(array_10_io_f_i),
    .io_ve_i(array_10_io_ve_i),
    .io_vf_i(array_10_io_vf_i),
    .io_vv_i(array_10_io_vv_i),
    .io_e_o(array_10_io_e_o),
    .io_f_o(array_10_io_f_o),
    .io_v_o(array_10_io_v_o)
  );
  SWCell array_11 ( // @[SWChisel.scala 170:39]
    .io_q(array_11_io_q),
    .io_r(array_11_io_r),
    .io_e_i(array_11_io_e_i),
    .io_f_i(array_11_io_f_i),
    .io_ve_i(array_11_io_ve_i),
    .io_vf_i(array_11_io_vf_i),
    .io_vv_i(array_11_io_vv_i),
    .io_e_o(array_11_io_e_o),
    .io_f_o(array_11_io_f_o),
    .io_v_o(array_11_io_v_o)
  );
  SWCell array_12 ( // @[SWChisel.scala 170:39]
    .io_q(array_12_io_q),
    .io_r(array_12_io_r),
    .io_e_i(array_12_io_e_i),
    .io_f_i(array_12_io_f_i),
    .io_ve_i(array_12_io_ve_i),
    .io_vf_i(array_12_io_vf_i),
    .io_vv_i(array_12_io_vv_i),
    .io_e_o(array_12_io_e_o),
    .io_f_o(array_12_io_f_o),
    .io_v_o(array_12_io_v_o)
  );
  SWCell array_13 ( // @[SWChisel.scala 170:39]
    .io_q(array_13_io_q),
    .io_r(array_13_io_r),
    .io_e_i(array_13_io_e_i),
    .io_f_i(array_13_io_f_i),
    .io_ve_i(array_13_io_ve_i),
    .io_vf_i(array_13_io_vf_i),
    .io_vv_i(array_13_io_vv_i),
    .io_e_o(array_13_io_e_o),
    .io_f_o(array_13_io_f_o),
    .io_v_o(array_13_io_v_o)
  );
  SWCell array_14 ( // @[SWChisel.scala 170:39]
    .io_q(array_14_io_q),
    .io_r(array_14_io_r),
    .io_e_i(array_14_io_e_i),
    .io_f_i(array_14_io_f_i),
    .io_ve_i(array_14_io_ve_i),
    .io_vf_i(array_14_io_vf_i),
    .io_vv_i(array_14_io_vv_i),
    .io_e_o(array_14_io_e_o),
    .io_f_o(array_14_io_f_o),
    .io_v_o(array_14_io_v_o)
  );
  SWCell array_15 ( // @[SWChisel.scala 170:39]
    .io_q(array_15_io_q),
    .io_r(array_15_io_r),
    .io_e_i(array_15_io_e_i),
    .io_f_i(array_15_io_f_i),
    .io_ve_i(array_15_io_ve_i),
    .io_vf_i(array_15_io_vf_i),
    .io_vv_i(array_15_io_vv_i),
    .io_e_o(array_15_io_e_o),
    .io_f_o(array_15_io_f_o),
    .io_v_o(array_15_io_v_o)
  );
  SWCell array_16 ( // @[SWChisel.scala 170:39]
    .io_q(array_16_io_q),
    .io_r(array_16_io_r),
    .io_e_i(array_16_io_e_i),
    .io_f_i(array_16_io_f_i),
    .io_ve_i(array_16_io_ve_i),
    .io_vf_i(array_16_io_vf_i),
    .io_vv_i(array_16_io_vv_i),
    .io_e_o(array_16_io_e_o),
    .io_f_o(array_16_io_f_o),
    .io_v_o(array_16_io_v_o)
  );
  SWCell array_17 ( // @[SWChisel.scala 170:39]
    .io_q(array_17_io_q),
    .io_r(array_17_io_r),
    .io_e_i(array_17_io_e_i),
    .io_f_i(array_17_io_f_i),
    .io_ve_i(array_17_io_ve_i),
    .io_vf_i(array_17_io_vf_i),
    .io_vv_i(array_17_io_vv_i),
    .io_e_o(array_17_io_e_o),
    .io_f_o(array_17_io_f_o),
    .io_v_o(array_17_io_v_o)
  );
  SWCell array_18 ( // @[SWChisel.scala 170:39]
    .io_q(array_18_io_q),
    .io_r(array_18_io_r),
    .io_e_i(array_18_io_e_i),
    .io_f_i(array_18_io_f_i),
    .io_ve_i(array_18_io_ve_i),
    .io_vf_i(array_18_io_vf_i),
    .io_vv_i(array_18_io_vv_i),
    .io_e_o(array_18_io_e_o),
    .io_f_o(array_18_io_f_o),
    .io_v_o(array_18_io_v_o)
  );
  SWCell array_19 ( // @[SWChisel.scala 170:39]
    .io_q(array_19_io_q),
    .io_r(array_19_io_r),
    .io_e_i(array_19_io_e_i),
    .io_f_i(array_19_io_f_i),
    .io_ve_i(array_19_io_ve_i),
    .io_vf_i(array_19_io_vf_i),
    .io_vv_i(array_19_io_vv_i),
    .io_e_o(array_19_io_e_o),
    .io_f_o(array_19_io_f_o),
    .io_v_o(array_19_io_v_o)
  );
  SWCell array_20 ( // @[SWChisel.scala 170:39]
    .io_q(array_20_io_q),
    .io_r(array_20_io_r),
    .io_e_i(array_20_io_e_i),
    .io_f_i(array_20_io_f_i),
    .io_ve_i(array_20_io_ve_i),
    .io_vf_i(array_20_io_vf_i),
    .io_vv_i(array_20_io_vv_i),
    .io_e_o(array_20_io_e_o),
    .io_f_o(array_20_io_f_o),
    .io_v_o(array_20_io_v_o)
  );
  SWCell array_21 ( // @[SWChisel.scala 170:39]
    .io_q(array_21_io_q),
    .io_r(array_21_io_r),
    .io_e_i(array_21_io_e_i),
    .io_f_i(array_21_io_f_i),
    .io_ve_i(array_21_io_ve_i),
    .io_vf_i(array_21_io_vf_i),
    .io_vv_i(array_21_io_vv_i),
    .io_e_o(array_21_io_e_o),
    .io_f_o(array_21_io_f_o),
    .io_v_o(array_21_io_v_o)
  );
  SWCell array_22 ( // @[SWChisel.scala 170:39]
    .io_q(array_22_io_q),
    .io_r(array_22_io_r),
    .io_e_i(array_22_io_e_i),
    .io_f_i(array_22_io_f_i),
    .io_ve_i(array_22_io_ve_i),
    .io_vf_i(array_22_io_vf_i),
    .io_vv_i(array_22_io_vv_i),
    .io_e_o(array_22_io_e_o),
    .io_f_o(array_22_io_f_o),
    .io_v_o(array_22_io_v_o)
  );
  SWCell array_23 ( // @[SWChisel.scala 170:39]
    .io_q(array_23_io_q),
    .io_r(array_23_io_r),
    .io_e_i(array_23_io_e_i),
    .io_f_i(array_23_io_f_i),
    .io_ve_i(array_23_io_ve_i),
    .io_vf_i(array_23_io_vf_i),
    .io_vv_i(array_23_io_vv_i),
    .io_e_o(array_23_io_e_o),
    .io_f_o(array_23_io_f_o),
    .io_v_o(array_23_io_v_o)
  );
  SWCell array_24 ( // @[SWChisel.scala 170:39]
    .io_q(array_24_io_q),
    .io_r(array_24_io_r),
    .io_e_i(array_24_io_e_i),
    .io_f_i(array_24_io_f_i),
    .io_ve_i(array_24_io_ve_i),
    .io_vf_i(array_24_io_vf_i),
    .io_vv_i(array_24_io_vv_i),
    .io_e_o(array_24_io_e_o),
    .io_f_o(array_24_io_f_o),
    .io_v_o(array_24_io_v_o)
  );
  SWCell array_25 ( // @[SWChisel.scala 170:39]
    .io_q(array_25_io_q),
    .io_r(array_25_io_r),
    .io_e_i(array_25_io_e_i),
    .io_f_i(array_25_io_f_i),
    .io_ve_i(array_25_io_ve_i),
    .io_vf_i(array_25_io_vf_i),
    .io_vv_i(array_25_io_vv_i),
    .io_e_o(array_25_io_e_o),
    .io_f_o(array_25_io_f_o),
    .io_v_o(array_25_io_v_o)
  );
  SWCell array_26 ( // @[SWChisel.scala 170:39]
    .io_q(array_26_io_q),
    .io_r(array_26_io_r),
    .io_e_i(array_26_io_e_i),
    .io_f_i(array_26_io_f_i),
    .io_ve_i(array_26_io_ve_i),
    .io_vf_i(array_26_io_vf_i),
    .io_vv_i(array_26_io_vv_i),
    .io_e_o(array_26_io_e_o),
    .io_f_o(array_26_io_f_o),
    .io_v_o(array_26_io_v_o)
  );
  SWCell array_27 ( // @[SWChisel.scala 170:39]
    .io_q(array_27_io_q),
    .io_r(array_27_io_r),
    .io_e_i(array_27_io_e_i),
    .io_f_i(array_27_io_f_i),
    .io_ve_i(array_27_io_ve_i),
    .io_vf_i(array_27_io_vf_i),
    .io_vv_i(array_27_io_vv_i),
    .io_e_o(array_27_io_e_o),
    .io_f_o(array_27_io_f_o),
    .io_v_o(array_27_io_v_o)
  );
  SWCell array_28 ( // @[SWChisel.scala 170:39]
    .io_q(array_28_io_q),
    .io_r(array_28_io_r),
    .io_e_i(array_28_io_e_i),
    .io_f_i(array_28_io_f_i),
    .io_ve_i(array_28_io_ve_i),
    .io_vf_i(array_28_io_vf_i),
    .io_vv_i(array_28_io_vv_i),
    .io_e_o(array_28_io_e_o),
    .io_f_o(array_28_io_f_o),
    .io_v_o(array_28_io_v_o)
  );
  SWCell array_29 ( // @[SWChisel.scala 170:39]
    .io_q(array_29_io_q),
    .io_r(array_29_io_r),
    .io_e_i(array_29_io_e_i),
    .io_f_i(array_29_io_f_i),
    .io_ve_i(array_29_io_ve_i),
    .io_vf_i(array_29_io_vf_i),
    .io_vv_i(array_29_io_vv_i),
    .io_e_o(array_29_io_e_o),
    .io_f_o(array_29_io_f_o),
    .io_v_o(array_29_io_v_o)
  );
  SWCell array_30 ( // @[SWChisel.scala 170:39]
    .io_q(array_30_io_q),
    .io_r(array_30_io_r),
    .io_e_i(array_30_io_e_i),
    .io_f_i(array_30_io_f_i),
    .io_ve_i(array_30_io_ve_i),
    .io_vf_i(array_30_io_vf_i),
    .io_vv_i(array_30_io_vv_i),
    .io_e_o(array_30_io_e_o),
    .io_f_o(array_30_io_f_o),
    .io_v_o(array_30_io_v_o)
  );
  SWCell array_31 ( // @[SWChisel.scala 170:39]
    .io_q(array_31_io_q),
    .io_r(array_31_io_r),
    .io_e_i(array_31_io_e_i),
    .io_f_i(array_31_io_f_i),
    .io_ve_i(array_31_io_ve_i),
    .io_vf_i(array_31_io_vf_i),
    .io_vv_i(array_31_io_vv_i),
    .io_e_o(array_31_io_e_o),
    .io_f_o(array_31_io_f_o),
    .io_v_o(array_31_io_v_o)
  );
  SWCell array_32 ( // @[SWChisel.scala 170:39]
    .io_q(array_32_io_q),
    .io_r(array_32_io_r),
    .io_e_i(array_32_io_e_i),
    .io_f_i(array_32_io_f_i),
    .io_ve_i(array_32_io_ve_i),
    .io_vf_i(array_32_io_vf_i),
    .io_vv_i(array_32_io_vv_i),
    .io_e_o(array_32_io_e_o),
    .io_f_o(array_32_io_f_o),
    .io_v_o(array_32_io_v_o)
  );
  SWCell array_33 ( // @[SWChisel.scala 170:39]
    .io_q(array_33_io_q),
    .io_r(array_33_io_r),
    .io_e_i(array_33_io_e_i),
    .io_f_i(array_33_io_f_i),
    .io_ve_i(array_33_io_ve_i),
    .io_vf_i(array_33_io_vf_i),
    .io_vv_i(array_33_io_vv_i),
    .io_e_o(array_33_io_e_o),
    .io_f_o(array_33_io_f_o),
    .io_v_o(array_33_io_v_o)
  );
  SWCell array_34 ( // @[SWChisel.scala 170:39]
    .io_q(array_34_io_q),
    .io_r(array_34_io_r),
    .io_e_i(array_34_io_e_i),
    .io_f_i(array_34_io_f_i),
    .io_ve_i(array_34_io_ve_i),
    .io_vf_i(array_34_io_vf_i),
    .io_vv_i(array_34_io_vv_i),
    .io_e_o(array_34_io_e_o),
    .io_f_o(array_34_io_f_o),
    .io_v_o(array_34_io_v_o)
  );
  SWCell array_35 ( // @[SWChisel.scala 170:39]
    .io_q(array_35_io_q),
    .io_r(array_35_io_r),
    .io_e_i(array_35_io_e_i),
    .io_f_i(array_35_io_f_i),
    .io_ve_i(array_35_io_ve_i),
    .io_vf_i(array_35_io_vf_i),
    .io_vv_i(array_35_io_vv_i),
    .io_e_o(array_35_io_e_o),
    .io_f_o(array_35_io_f_o),
    .io_v_o(array_35_io_v_o)
  );
  SWCell array_36 ( // @[SWChisel.scala 170:39]
    .io_q(array_36_io_q),
    .io_r(array_36_io_r),
    .io_e_i(array_36_io_e_i),
    .io_f_i(array_36_io_f_i),
    .io_ve_i(array_36_io_ve_i),
    .io_vf_i(array_36_io_vf_i),
    .io_vv_i(array_36_io_vv_i),
    .io_e_o(array_36_io_e_o),
    .io_f_o(array_36_io_f_o),
    .io_v_o(array_36_io_v_o)
  );
  SWCell array_37 ( // @[SWChisel.scala 170:39]
    .io_q(array_37_io_q),
    .io_r(array_37_io_r),
    .io_e_i(array_37_io_e_i),
    .io_f_i(array_37_io_f_i),
    .io_ve_i(array_37_io_ve_i),
    .io_vf_i(array_37_io_vf_i),
    .io_vv_i(array_37_io_vv_i),
    .io_e_o(array_37_io_e_o),
    .io_f_o(array_37_io_f_o),
    .io_v_o(array_37_io_v_o)
  );
  SWCell array_38 ( // @[SWChisel.scala 170:39]
    .io_q(array_38_io_q),
    .io_r(array_38_io_r),
    .io_e_i(array_38_io_e_i),
    .io_f_i(array_38_io_f_i),
    .io_ve_i(array_38_io_ve_i),
    .io_vf_i(array_38_io_vf_i),
    .io_vv_i(array_38_io_vv_i),
    .io_e_o(array_38_io_e_o),
    .io_f_o(array_38_io_f_o),
    .io_v_o(array_38_io_v_o)
  );
  SWCell array_39 ( // @[SWChisel.scala 170:39]
    .io_q(array_39_io_q),
    .io_r(array_39_io_r),
    .io_e_i(array_39_io_e_i),
    .io_f_i(array_39_io_f_i),
    .io_ve_i(array_39_io_ve_i),
    .io_vf_i(array_39_io_vf_i),
    .io_vv_i(array_39_io_vv_i),
    .io_e_o(array_39_io_e_o),
    .io_f_o(array_39_io_f_o),
    .io_v_o(array_39_io_v_o)
  );
  SWCell array_40 ( // @[SWChisel.scala 170:39]
    .io_q(array_40_io_q),
    .io_r(array_40_io_r),
    .io_e_i(array_40_io_e_i),
    .io_f_i(array_40_io_f_i),
    .io_ve_i(array_40_io_ve_i),
    .io_vf_i(array_40_io_vf_i),
    .io_vv_i(array_40_io_vv_i),
    .io_e_o(array_40_io_e_o),
    .io_f_o(array_40_io_f_o),
    .io_v_o(array_40_io_v_o)
  );
  SWCell array_41 ( // @[SWChisel.scala 170:39]
    .io_q(array_41_io_q),
    .io_r(array_41_io_r),
    .io_e_i(array_41_io_e_i),
    .io_f_i(array_41_io_f_i),
    .io_ve_i(array_41_io_ve_i),
    .io_vf_i(array_41_io_vf_i),
    .io_vv_i(array_41_io_vv_i),
    .io_e_o(array_41_io_e_o),
    .io_f_o(array_41_io_f_o),
    .io_v_o(array_41_io_v_o)
  );
  SWCell array_42 ( // @[SWChisel.scala 170:39]
    .io_q(array_42_io_q),
    .io_r(array_42_io_r),
    .io_e_i(array_42_io_e_i),
    .io_f_i(array_42_io_f_i),
    .io_ve_i(array_42_io_ve_i),
    .io_vf_i(array_42_io_vf_i),
    .io_vv_i(array_42_io_vv_i),
    .io_e_o(array_42_io_e_o),
    .io_f_o(array_42_io_f_o),
    .io_v_o(array_42_io_v_o)
  );
  SWCell array_43 ( // @[SWChisel.scala 170:39]
    .io_q(array_43_io_q),
    .io_r(array_43_io_r),
    .io_e_i(array_43_io_e_i),
    .io_f_i(array_43_io_f_i),
    .io_ve_i(array_43_io_ve_i),
    .io_vf_i(array_43_io_vf_i),
    .io_vv_i(array_43_io_vv_i),
    .io_e_o(array_43_io_e_o),
    .io_f_o(array_43_io_f_o),
    .io_v_o(array_43_io_v_o)
  );
  SWCell array_44 ( // @[SWChisel.scala 170:39]
    .io_q(array_44_io_q),
    .io_r(array_44_io_r),
    .io_e_i(array_44_io_e_i),
    .io_f_i(array_44_io_f_i),
    .io_ve_i(array_44_io_ve_i),
    .io_vf_i(array_44_io_vf_i),
    .io_vv_i(array_44_io_vv_i),
    .io_e_o(array_44_io_e_o),
    .io_f_o(array_44_io_f_o),
    .io_v_o(array_44_io_v_o)
  );
  SWCell array_45 ( // @[SWChisel.scala 170:39]
    .io_q(array_45_io_q),
    .io_r(array_45_io_r),
    .io_e_i(array_45_io_e_i),
    .io_f_i(array_45_io_f_i),
    .io_ve_i(array_45_io_ve_i),
    .io_vf_i(array_45_io_vf_i),
    .io_vv_i(array_45_io_vv_i),
    .io_e_o(array_45_io_e_o),
    .io_f_o(array_45_io_f_o),
    .io_v_o(array_45_io_v_o)
  );
  SWCell array_46 ( // @[SWChisel.scala 170:39]
    .io_q(array_46_io_q),
    .io_r(array_46_io_r),
    .io_e_i(array_46_io_e_i),
    .io_f_i(array_46_io_f_i),
    .io_ve_i(array_46_io_ve_i),
    .io_vf_i(array_46_io_vf_i),
    .io_vv_i(array_46_io_vv_i),
    .io_e_o(array_46_io_e_o),
    .io_f_o(array_46_io_f_o),
    .io_v_o(array_46_io_v_o)
  );
  SWCell array_47 ( // @[SWChisel.scala 170:39]
    .io_q(array_47_io_q),
    .io_r(array_47_io_r),
    .io_e_i(array_47_io_e_i),
    .io_f_i(array_47_io_f_i),
    .io_ve_i(array_47_io_ve_i),
    .io_vf_i(array_47_io_vf_i),
    .io_vv_i(array_47_io_vv_i),
    .io_e_o(array_47_io_e_o),
    .io_f_o(array_47_io_f_o),
    .io_v_o(array_47_io_v_o)
  );
  SWCell array_48 ( // @[SWChisel.scala 170:39]
    .io_q(array_48_io_q),
    .io_r(array_48_io_r),
    .io_e_i(array_48_io_e_i),
    .io_f_i(array_48_io_f_i),
    .io_ve_i(array_48_io_ve_i),
    .io_vf_i(array_48_io_vf_i),
    .io_vv_i(array_48_io_vv_i),
    .io_e_o(array_48_io_e_o),
    .io_f_o(array_48_io_f_o),
    .io_v_o(array_48_io_v_o)
  );
  SWCell array_49 ( // @[SWChisel.scala 170:39]
    .io_q(array_49_io_q),
    .io_r(array_49_io_r),
    .io_e_i(array_49_io_e_i),
    .io_f_i(array_49_io_f_i),
    .io_ve_i(array_49_io_ve_i),
    .io_vf_i(array_49_io_vf_i),
    .io_vv_i(array_49_io_vv_i),
    .io_e_o(array_49_io_e_o),
    .io_f_o(array_49_io_f_o),
    .io_v_o(array_49_io_v_o)
  );
  MyCounter r_count_0 ( // @[SWChisel.scala 171:41]
    .clock(r_count_0_clock),
    .reset(r_count_0_reset),
    .io_en(r_count_0_io_en),
    .io_out(r_count_0_io_out)
  );
  MyCounter r_count_1 ( // @[SWChisel.scala 171:41]
    .clock(r_count_1_clock),
    .reset(r_count_1_reset),
    .io_en(r_count_1_io_en),
    .io_out(r_count_1_io_out)
  );
  MyCounter r_count_2 ( // @[SWChisel.scala 171:41]
    .clock(r_count_2_clock),
    .reset(r_count_2_reset),
    .io_en(r_count_2_io_en),
    .io_out(r_count_2_io_out)
  );
  MyCounter r_count_3 ( // @[SWChisel.scala 171:41]
    .clock(r_count_3_clock),
    .reset(r_count_3_reset),
    .io_en(r_count_3_io_en),
    .io_out(r_count_3_io_out)
  );
  MyCounter r_count_4 ( // @[SWChisel.scala 171:41]
    .clock(r_count_4_clock),
    .reset(r_count_4_reset),
    .io_en(r_count_4_io_en),
    .io_out(r_count_4_io_out)
  );
  MyCounter r_count_5 ( // @[SWChisel.scala 171:41]
    .clock(r_count_5_clock),
    .reset(r_count_5_reset),
    .io_en(r_count_5_io_en),
    .io_out(r_count_5_io_out)
  );
  MyCounter r_count_6 ( // @[SWChisel.scala 171:41]
    .clock(r_count_6_clock),
    .reset(r_count_6_reset),
    .io_en(r_count_6_io_en),
    .io_out(r_count_6_io_out)
  );
  MyCounter r_count_7 ( // @[SWChisel.scala 171:41]
    .clock(r_count_7_clock),
    .reset(r_count_7_reset),
    .io_en(r_count_7_io_en),
    .io_out(r_count_7_io_out)
  );
  MyCounter r_count_8 ( // @[SWChisel.scala 171:41]
    .clock(r_count_8_clock),
    .reset(r_count_8_reset),
    .io_en(r_count_8_io_en),
    .io_out(r_count_8_io_out)
  );
  MyCounter r_count_9 ( // @[SWChisel.scala 171:41]
    .clock(r_count_9_clock),
    .reset(r_count_9_reset),
    .io_en(r_count_9_io_en),
    .io_out(r_count_9_io_out)
  );
  MyCounter r_count_10 ( // @[SWChisel.scala 171:41]
    .clock(r_count_10_clock),
    .reset(r_count_10_reset),
    .io_en(r_count_10_io_en),
    .io_out(r_count_10_io_out)
  );
  MyCounter r_count_11 ( // @[SWChisel.scala 171:41]
    .clock(r_count_11_clock),
    .reset(r_count_11_reset),
    .io_en(r_count_11_io_en),
    .io_out(r_count_11_io_out)
  );
  MyCounter r_count_12 ( // @[SWChisel.scala 171:41]
    .clock(r_count_12_clock),
    .reset(r_count_12_reset),
    .io_en(r_count_12_io_en),
    .io_out(r_count_12_io_out)
  );
  MyCounter r_count_13 ( // @[SWChisel.scala 171:41]
    .clock(r_count_13_clock),
    .reset(r_count_13_reset),
    .io_en(r_count_13_io_en),
    .io_out(r_count_13_io_out)
  );
  MyCounter r_count_14 ( // @[SWChisel.scala 171:41]
    .clock(r_count_14_clock),
    .reset(r_count_14_reset),
    .io_en(r_count_14_io_en),
    .io_out(r_count_14_io_out)
  );
  MyCounter r_count_15 ( // @[SWChisel.scala 171:41]
    .clock(r_count_15_clock),
    .reset(r_count_15_reset),
    .io_en(r_count_15_io_en),
    .io_out(r_count_15_io_out)
  );
  MyCounter r_count_16 ( // @[SWChisel.scala 171:41]
    .clock(r_count_16_clock),
    .reset(r_count_16_reset),
    .io_en(r_count_16_io_en),
    .io_out(r_count_16_io_out)
  );
  MyCounter r_count_17 ( // @[SWChisel.scala 171:41]
    .clock(r_count_17_clock),
    .reset(r_count_17_reset),
    .io_en(r_count_17_io_en),
    .io_out(r_count_17_io_out)
  );
  MyCounter r_count_18 ( // @[SWChisel.scala 171:41]
    .clock(r_count_18_clock),
    .reset(r_count_18_reset),
    .io_en(r_count_18_io_en),
    .io_out(r_count_18_io_out)
  );
  MyCounter r_count_19 ( // @[SWChisel.scala 171:41]
    .clock(r_count_19_clock),
    .reset(r_count_19_reset),
    .io_en(r_count_19_io_en),
    .io_out(r_count_19_io_out)
  );
  MyCounter r_count_20 ( // @[SWChisel.scala 171:41]
    .clock(r_count_20_clock),
    .reset(r_count_20_reset),
    .io_en(r_count_20_io_en),
    .io_out(r_count_20_io_out)
  );
  MyCounter r_count_21 ( // @[SWChisel.scala 171:41]
    .clock(r_count_21_clock),
    .reset(r_count_21_reset),
    .io_en(r_count_21_io_en),
    .io_out(r_count_21_io_out)
  );
  MyCounter r_count_22 ( // @[SWChisel.scala 171:41]
    .clock(r_count_22_clock),
    .reset(r_count_22_reset),
    .io_en(r_count_22_io_en),
    .io_out(r_count_22_io_out)
  );
  MyCounter r_count_23 ( // @[SWChisel.scala 171:41]
    .clock(r_count_23_clock),
    .reset(r_count_23_reset),
    .io_en(r_count_23_io_en),
    .io_out(r_count_23_io_out)
  );
  MyCounter r_count_24 ( // @[SWChisel.scala 171:41]
    .clock(r_count_24_clock),
    .reset(r_count_24_reset),
    .io_en(r_count_24_io_en),
    .io_out(r_count_24_io_out)
  );
  MyCounter r_count_25 ( // @[SWChisel.scala 171:41]
    .clock(r_count_25_clock),
    .reset(r_count_25_reset),
    .io_en(r_count_25_io_en),
    .io_out(r_count_25_io_out)
  );
  MyCounter r_count_26 ( // @[SWChisel.scala 171:41]
    .clock(r_count_26_clock),
    .reset(r_count_26_reset),
    .io_en(r_count_26_io_en),
    .io_out(r_count_26_io_out)
  );
  MyCounter r_count_27 ( // @[SWChisel.scala 171:41]
    .clock(r_count_27_clock),
    .reset(r_count_27_reset),
    .io_en(r_count_27_io_en),
    .io_out(r_count_27_io_out)
  );
  MyCounter r_count_28 ( // @[SWChisel.scala 171:41]
    .clock(r_count_28_clock),
    .reset(r_count_28_reset),
    .io_en(r_count_28_io_en),
    .io_out(r_count_28_io_out)
  );
  MyCounter r_count_29 ( // @[SWChisel.scala 171:41]
    .clock(r_count_29_clock),
    .reset(r_count_29_reset),
    .io_en(r_count_29_io_en),
    .io_out(r_count_29_io_out)
  );
  MyCounter r_count_30 ( // @[SWChisel.scala 171:41]
    .clock(r_count_30_clock),
    .reset(r_count_30_reset),
    .io_en(r_count_30_io_en),
    .io_out(r_count_30_io_out)
  );
  MyCounter r_count_31 ( // @[SWChisel.scala 171:41]
    .clock(r_count_31_clock),
    .reset(r_count_31_reset),
    .io_en(r_count_31_io_en),
    .io_out(r_count_31_io_out)
  );
  MyCounter r_count_32 ( // @[SWChisel.scala 171:41]
    .clock(r_count_32_clock),
    .reset(r_count_32_reset),
    .io_en(r_count_32_io_en),
    .io_out(r_count_32_io_out)
  );
  MyCounter r_count_33 ( // @[SWChisel.scala 171:41]
    .clock(r_count_33_clock),
    .reset(r_count_33_reset),
    .io_en(r_count_33_io_en),
    .io_out(r_count_33_io_out)
  );
  MyCounter r_count_34 ( // @[SWChisel.scala 171:41]
    .clock(r_count_34_clock),
    .reset(r_count_34_reset),
    .io_en(r_count_34_io_en),
    .io_out(r_count_34_io_out)
  );
  MyCounter r_count_35 ( // @[SWChisel.scala 171:41]
    .clock(r_count_35_clock),
    .reset(r_count_35_reset),
    .io_en(r_count_35_io_en),
    .io_out(r_count_35_io_out)
  );
  MyCounter r_count_36 ( // @[SWChisel.scala 171:41]
    .clock(r_count_36_clock),
    .reset(r_count_36_reset),
    .io_en(r_count_36_io_en),
    .io_out(r_count_36_io_out)
  );
  MyCounter r_count_37 ( // @[SWChisel.scala 171:41]
    .clock(r_count_37_clock),
    .reset(r_count_37_reset),
    .io_en(r_count_37_io_en),
    .io_out(r_count_37_io_out)
  );
  MyCounter r_count_38 ( // @[SWChisel.scala 171:41]
    .clock(r_count_38_clock),
    .reset(r_count_38_reset),
    .io_en(r_count_38_io_en),
    .io_out(r_count_38_io_out)
  );
  MyCounter r_count_39 ( // @[SWChisel.scala 171:41]
    .clock(r_count_39_clock),
    .reset(r_count_39_reset),
    .io_en(r_count_39_io_en),
    .io_out(r_count_39_io_out)
  );
  MyCounter r_count_40 ( // @[SWChisel.scala 171:41]
    .clock(r_count_40_clock),
    .reset(r_count_40_reset),
    .io_en(r_count_40_io_en),
    .io_out(r_count_40_io_out)
  );
  MyCounter r_count_41 ( // @[SWChisel.scala 171:41]
    .clock(r_count_41_clock),
    .reset(r_count_41_reset),
    .io_en(r_count_41_io_en),
    .io_out(r_count_41_io_out)
  );
  MyCounter r_count_42 ( // @[SWChisel.scala 171:41]
    .clock(r_count_42_clock),
    .reset(r_count_42_reset),
    .io_en(r_count_42_io_en),
    .io_out(r_count_42_io_out)
  );
  MyCounter r_count_43 ( // @[SWChisel.scala 171:41]
    .clock(r_count_43_clock),
    .reset(r_count_43_reset),
    .io_en(r_count_43_io_en),
    .io_out(r_count_43_io_out)
  );
  MyCounter r_count_44 ( // @[SWChisel.scala 171:41]
    .clock(r_count_44_clock),
    .reset(r_count_44_reset),
    .io_en(r_count_44_io_en),
    .io_out(r_count_44_io_out)
  );
  MyCounter r_count_45 ( // @[SWChisel.scala 171:41]
    .clock(r_count_45_clock),
    .reset(r_count_45_reset),
    .io_en(r_count_45_io_en),
    .io_out(r_count_45_io_out)
  );
  MyCounter r_count_46 ( // @[SWChisel.scala 171:41]
    .clock(r_count_46_clock),
    .reset(r_count_46_reset),
    .io_en(r_count_46_io_en),
    .io_out(r_count_46_io_out)
  );
  MyCounter r_count_47 ( // @[SWChisel.scala 171:41]
    .clock(r_count_47_clock),
    .reset(r_count_47_reset),
    .io_en(r_count_47_io_en),
    .io_out(r_count_47_io_out)
  );
  MyCounter r_count_48 ( // @[SWChisel.scala 171:41]
    .clock(r_count_48_clock),
    .reset(r_count_48_reset),
    .io_en(r_count_48_io_en),
    .io_out(r_count_48_io_out)
  );
  MyCounter r_count_49 ( // @[SWChisel.scala 171:41]
    .clock(r_count_49_clock),
    .reset(r_count_49_reset),
    .io_en(r_count_49_io_en),
    .io_out(r_count_49_io_out)
  );
  MAX max ( // @[SWChisel.scala 174:19]
    .clock(max_clock),
    .reset(max_reset),
    .io_start(max_io_start),
    .io_in(max_io_in),
    .io_done(max_io_done),
    .io_out(max_io_out)
  );
  assign io_result = max_io_out; // @[SWChisel.scala 181:13]
  assign io_done = max_io_done; // @[SWChisel.scala 182:11]
  assign array_0_io_q = io_q_0_b; // @[SWChisel.scala 220:19]
  assign array_0_io_r = 7'h63 == r_count_0_io_out ? io_r_99_b : _GEN_248; // @[SWChisel.scala 221:{19,19}]
  assign array_0_io_e_i = E_0; // @[SWChisel.scala 196:21]
  assign array_0_io_f_i = 16'sh0; // @[SWChisel.scala 198:21]
  assign array_0_io_ve_i = V1_1; // @[SWChisel.scala 197:22]
  assign array_0_io_vf_i = V1_0; // @[SWChisel.scala 199:22]
  assign array_0_io_vv_i = V2_0; // @[SWChisel.scala 200:22]
  assign array_1_io_q = io_q_1_b; // @[SWChisel.scala 220:19]
  assign array_1_io_r = 7'h63 == r_count_1_io_out ? io_r_99_b : _GEN_348; // @[SWChisel.scala 221:{19,19}]
  assign array_1_io_e_i = E_1; // @[SWChisel.scala 196:21]
  assign array_1_io_f_i = F_1; // @[SWChisel.scala 198:21]
  assign array_1_io_ve_i = V1_2; // @[SWChisel.scala 197:22]
  assign array_1_io_vf_i = V1_1; // @[SWChisel.scala 199:22]
  assign array_1_io_vv_i = V2_1; // @[SWChisel.scala 200:22]
  assign array_2_io_q = io_q_2_b; // @[SWChisel.scala 220:19]
  assign array_2_io_r = 7'h63 == r_count_2_io_out ? io_r_99_b : _GEN_448; // @[SWChisel.scala 221:{19,19}]
  assign array_2_io_e_i = E_2; // @[SWChisel.scala 196:21]
  assign array_2_io_f_i = F_2; // @[SWChisel.scala 198:21]
  assign array_2_io_ve_i = V1_3; // @[SWChisel.scala 197:22]
  assign array_2_io_vf_i = V1_2; // @[SWChisel.scala 199:22]
  assign array_2_io_vv_i = V2_2; // @[SWChisel.scala 200:22]
  assign array_3_io_q = io_q_3_b; // @[SWChisel.scala 220:19]
  assign array_3_io_r = 7'h63 == r_count_3_io_out ? io_r_99_b : _GEN_548; // @[SWChisel.scala 221:{19,19}]
  assign array_3_io_e_i = E_3; // @[SWChisel.scala 196:21]
  assign array_3_io_f_i = F_3; // @[SWChisel.scala 198:21]
  assign array_3_io_ve_i = V1_4; // @[SWChisel.scala 197:22]
  assign array_3_io_vf_i = V1_3; // @[SWChisel.scala 199:22]
  assign array_3_io_vv_i = V2_3; // @[SWChisel.scala 200:22]
  assign array_4_io_q = io_q_4_b; // @[SWChisel.scala 220:19]
  assign array_4_io_r = 7'h63 == r_count_4_io_out ? io_r_99_b : _GEN_648; // @[SWChisel.scala 221:{19,19}]
  assign array_4_io_e_i = E_4; // @[SWChisel.scala 196:21]
  assign array_4_io_f_i = F_4; // @[SWChisel.scala 198:21]
  assign array_4_io_ve_i = V1_5; // @[SWChisel.scala 197:22]
  assign array_4_io_vf_i = V1_4; // @[SWChisel.scala 199:22]
  assign array_4_io_vv_i = V2_4; // @[SWChisel.scala 200:22]
  assign array_5_io_q = io_q_5_b; // @[SWChisel.scala 220:19]
  assign array_5_io_r = 7'h63 == r_count_5_io_out ? io_r_99_b : _GEN_748; // @[SWChisel.scala 221:{19,19}]
  assign array_5_io_e_i = E_5; // @[SWChisel.scala 196:21]
  assign array_5_io_f_i = F_5; // @[SWChisel.scala 198:21]
  assign array_5_io_ve_i = V1_6; // @[SWChisel.scala 197:22]
  assign array_5_io_vf_i = V1_5; // @[SWChisel.scala 199:22]
  assign array_5_io_vv_i = V2_5; // @[SWChisel.scala 200:22]
  assign array_6_io_q = io_q_6_b; // @[SWChisel.scala 220:19]
  assign array_6_io_r = 7'h63 == r_count_6_io_out ? io_r_99_b : _GEN_848; // @[SWChisel.scala 221:{19,19}]
  assign array_6_io_e_i = E_6; // @[SWChisel.scala 196:21]
  assign array_6_io_f_i = F_6; // @[SWChisel.scala 198:21]
  assign array_6_io_ve_i = V1_7; // @[SWChisel.scala 197:22]
  assign array_6_io_vf_i = V1_6; // @[SWChisel.scala 199:22]
  assign array_6_io_vv_i = V2_6; // @[SWChisel.scala 200:22]
  assign array_7_io_q = io_q_7_b; // @[SWChisel.scala 220:19]
  assign array_7_io_r = 7'h63 == r_count_7_io_out ? io_r_99_b : _GEN_948; // @[SWChisel.scala 221:{19,19}]
  assign array_7_io_e_i = E_7; // @[SWChisel.scala 196:21]
  assign array_7_io_f_i = F_7; // @[SWChisel.scala 198:21]
  assign array_7_io_ve_i = V1_8; // @[SWChisel.scala 197:22]
  assign array_7_io_vf_i = V1_7; // @[SWChisel.scala 199:22]
  assign array_7_io_vv_i = V2_7; // @[SWChisel.scala 200:22]
  assign array_8_io_q = io_q_8_b; // @[SWChisel.scala 220:19]
  assign array_8_io_r = 7'h63 == r_count_8_io_out ? io_r_99_b : _GEN_1048; // @[SWChisel.scala 221:{19,19}]
  assign array_8_io_e_i = E_8; // @[SWChisel.scala 196:21]
  assign array_8_io_f_i = F_8; // @[SWChisel.scala 198:21]
  assign array_8_io_ve_i = V1_9; // @[SWChisel.scala 197:22]
  assign array_8_io_vf_i = V1_8; // @[SWChisel.scala 199:22]
  assign array_8_io_vv_i = V2_8; // @[SWChisel.scala 200:22]
  assign array_9_io_q = io_q_9_b; // @[SWChisel.scala 220:19]
  assign array_9_io_r = 7'h63 == r_count_9_io_out ? io_r_99_b : _GEN_1148; // @[SWChisel.scala 221:{19,19}]
  assign array_9_io_e_i = E_9; // @[SWChisel.scala 196:21]
  assign array_9_io_f_i = F_9; // @[SWChisel.scala 198:21]
  assign array_9_io_ve_i = V1_10; // @[SWChisel.scala 197:22]
  assign array_9_io_vf_i = V1_9; // @[SWChisel.scala 199:22]
  assign array_9_io_vv_i = V2_9; // @[SWChisel.scala 200:22]
  assign array_10_io_q = io_q_10_b; // @[SWChisel.scala 220:19]
  assign array_10_io_r = 7'h63 == r_count_10_io_out ? io_r_99_b : _GEN_1248; // @[SWChisel.scala 221:{19,19}]
  assign array_10_io_e_i = E_10; // @[SWChisel.scala 196:21]
  assign array_10_io_f_i = F_10; // @[SWChisel.scala 198:21]
  assign array_10_io_ve_i = V1_11; // @[SWChisel.scala 197:22]
  assign array_10_io_vf_i = V1_10; // @[SWChisel.scala 199:22]
  assign array_10_io_vv_i = V2_10; // @[SWChisel.scala 200:22]
  assign array_11_io_q = io_q_11_b; // @[SWChisel.scala 220:19]
  assign array_11_io_r = 7'h63 == r_count_11_io_out ? io_r_99_b : _GEN_1348; // @[SWChisel.scala 221:{19,19}]
  assign array_11_io_e_i = E_11; // @[SWChisel.scala 196:21]
  assign array_11_io_f_i = F_11; // @[SWChisel.scala 198:21]
  assign array_11_io_ve_i = V1_12; // @[SWChisel.scala 197:22]
  assign array_11_io_vf_i = V1_11; // @[SWChisel.scala 199:22]
  assign array_11_io_vv_i = V2_11; // @[SWChisel.scala 200:22]
  assign array_12_io_q = io_q_12_b; // @[SWChisel.scala 220:19]
  assign array_12_io_r = 7'h63 == r_count_12_io_out ? io_r_99_b : _GEN_1448; // @[SWChisel.scala 221:{19,19}]
  assign array_12_io_e_i = E_12; // @[SWChisel.scala 196:21]
  assign array_12_io_f_i = F_12; // @[SWChisel.scala 198:21]
  assign array_12_io_ve_i = V1_13; // @[SWChisel.scala 197:22]
  assign array_12_io_vf_i = V1_12; // @[SWChisel.scala 199:22]
  assign array_12_io_vv_i = V2_12; // @[SWChisel.scala 200:22]
  assign array_13_io_q = io_q_13_b; // @[SWChisel.scala 220:19]
  assign array_13_io_r = 7'h63 == r_count_13_io_out ? io_r_99_b : _GEN_1548; // @[SWChisel.scala 221:{19,19}]
  assign array_13_io_e_i = E_13; // @[SWChisel.scala 196:21]
  assign array_13_io_f_i = F_13; // @[SWChisel.scala 198:21]
  assign array_13_io_ve_i = V1_14; // @[SWChisel.scala 197:22]
  assign array_13_io_vf_i = V1_13; // @[SWChisel.scala 199:22]
  assign array_13_io_vv_i = V2_13; // @[SWChisel.scala 200:22]
  assign array_14_io_q = io_q_14_b; // @[SWChisel.scala 220:19]
  assign array_14_io_r = 7'h63 == r_count_14_io_out ? io_r_99_b : _GEN_1648; // @[SWChisel.scala 221:{19,19}]
  assign array_14_io_e_i = E_14; // @[SWChisel.scala 196:21]
  assign array_14_io_f_i = F_14; // @[SWChisel.scala 198:21]
  assign array_14_io_ve_i = V1_15; // @[SWChisel.scala 197:22]
  assign array_14_io_vf_i = V1_14; // @[SWChisel.scala 199:22]
  assign array_14_io_vv_i = V2_14; // @[SWChisel.scala 200:22]
  assign array_15_io_q = io_q_15_b; // @[SWChisel.scala 220:19]
  assign array_15_io_r = 7'h63 == r_count_15_io_out ? io_r_99_b : _GEN_1748; // @[SWChisel.scala 221:{19,19}]
  assign array_15_io_e_i = E_15; // @[SWChisel.scala 196:21]
  assign array_15_io_f_i = F_15; // @[SWChisel.scala 198:21]
  assign array_15_io_ve_i = V1_16; // @[SWChisel.scala 197:22]
  assign array_15_io_vf_i = V1_15; // @[SWChisel.scala 199:22]
  assign array_15_io_vv_i = V2_15; // @[SWChisel.scala 200:22]
  assign array_16_io_q = io_q_16_b; // @[SWChisel.scala 220:19]
  assign array_16_io_r = 7'h63 == r_count_16_io_out ? io_r_99_b : _GEN_1848; // @[SWChisel.scala 221:{19,19}]
  assign array_16_io_e_i = E_16; // @[SWChisel.scala 196:21]
  assign array_16_io_f_i = F_16; // @[SWChisel.scala 198:21]
  assign array_16_io_ve_i = V1_17; // @[SWChisel.scala 197:22]
  assign array_16_io_vf_i = V1_16; // @[SWChisel.scala 199:22]
  assign array_16_io_vv_i = V2_16; // @[SWChisel.scala 200:22]
  assign array_17_io_q = io_q_17_b; // @[SWChisel.scala 220:19]
  assign array_17_io_r = 7'h63 == r_count_17_io_out ? io_r_99_b : _GEN_1948; // @[SWChisel.scala 221:{19,19}]
  assign array_17_io_e_i = E_17; // @[SWChisel.scala 196:21]
  assign array_17_io_f_i = F_17; // @[SWChisel.scala 198:21]
  assign array_17_io_ve_i = V1_18; // @[SWChisel.scala 197:22]
  assign array_17_io_vf_i = V1_17; // @[SWChisel.scala 199:22]
  assign array_17_io_vv_i = V2_17; // @[SWChisel.scala 200:22]
  assign array_18_io_q = io_q_18_b; // @[SWChisel.scala 220:19]
  assign array_18_io_r = 7'h63 == r_count_18_io_out ? io_r_99_b : _GEN_2048; // @[SWChisel.scala 221:{19,19}]
  assign array_18_io_e_i = E_18; // @[SWChisel.scala 196:21]
  assign array_18_io_f_i = F_18; // @[SWChisel.scala 198:21]
  assign array_18_io_ve_i = V1_19; // @[SWChisel.scala 197:22]
  assign array_18_io_vf_i = V1_18; // @[SWChisel.scala 199:22]
  assign array_18_io_vv_i = V2_18; // @[SWChisel.scala 200:22]
  assign array_19_io_q = io_q_19_b; // @[SWChisel.scala 220:19]
  assign array_19_io_r = 7'h63 == r_count_19_io_out ? io_r_99_b : _GEN_2148; // @[SWChisel.scala 221:{19,19}]
  assign array_19_io_e_i = E_19; // @[SWChisel.scala 196:21]
  assign array_19_io_f_i = F_19; // @[SWChisel.scala 198:21]
  assign array_19_io_ve_i = V1_20; // @[SWChisel.scala 197:22]
  assign array_19_io_vf_i = V1_19; // @[SWChisel.scala 199:22]
  assign array_19_io_vv_i = V2_19; // @[SWChisel.scala 200:22]
  assign array_20_io_q = io_q_20_b; // @[SWChisel.scala 220:19]
  assign array_20_io_r = 7'h63 == r_count_20_io_out ? io_r_99_b : _GEN_2248; // @[SWChisel.scala 221:{19,19}]
  assign array_20_io_e_i = E_20; // @[SWChisel.scala 196:21]
  assign array_20_io_f_i = F_20; // @[SWChisel.scala 198:21]
  assign array_20_io_ve_i = V1_21; // @[SWChisel.scala 197:22]
  assign array_20_io_vf_i = V1_20; // @[SWChisel.scala 199:22]
  assign array_20_io_vv_i = V2_20; // @[SWChisel.scala 200:22]
  assign array_21_io_q = io_q_21_b; // @[SWChisel.scala 220:19]
  assign array_21_io_r = 7'h63 == r_count_21_io_out ? io_r_99_b : _GEN_2348; // @[SWChisel.scala 221:{19,19}]
  assign array_21_io_e_i = E_21; // @[SWChisel.scala 196:21]
  assign array_21_io_f_i = F_21; // @[SWChisel.scala 198:21]
  assign array_21_io_ve_i = V1_22; // @[SWChisel.scala 197:22]
  assign array_21_io_vf_i = V1_21; // @[SWChisel.scala 199:22]
  assign array_21_io_vv_i = V2_21; // @[SWChisel.scala 200:22]
  assign array_22_io_q = io_q_22_b; // @[SWChisel.scala 220:19]
  assign array_22_io_r = 7'h63 == r_count_22_io_out ? io_r_99_b : _GEN_2448; // @[SWChisel.scala 221:{19,19}]
  assign array_22_io_e_i = E_22; // @[SWChisel.scala 196:21]
  assign array_22_io_f_i = F_22; // @[SWChisel.scala 198:21]
  assign array_22_io_ve_i = V1_23; // @[SWChisel.scala 197:22]
  assign array_22_io_vf_i = V1_22; // @[SWChisel.scala 199:22]
  assign array_22_io_vv_i = V2_22; // @[SWChisel.scala 200:22]
  assign array_23_io_q = io_q_23_b; // @[SWChisel.scala 220:19]
  assign array_23_io_r = 7'h63 == r_count_23_io_out ? io_r_99_b : _GEN_2548; // @[SWChisel.scala 221:{19,19}]
  assign array_23_io_e_i = E_23; // @[SWChisel.scala 196:21]
  assign array_23_io_f_i = F_23; // @[SWChisel.scala 198:21]
  assign array_23_io_ve_i = V1_24; // @[SWChisel.scala 197:22]
  assign array_23_io_vf_i = V1_23; // @[SWChisel.scala 199:22]
  assign array_23_io_vv_i = V2_23; // @[SWChisel.scala 200:22]
  assign array_24_io_q = io_q_24_b; // @[SWChisel.scala 220:19]
  assign array_24_io_r = 7'h63 == r_count_24_io_out ? io_r_99_b : _GEN_2648; // @[SWChisel.scala 221:{19,19}]
  assign array_24_io_e_i = E_24; // @[SWChisel.scala 196:21]
  assign array_24_io_f_i = F_24; // @[SWChisel.scala 198:21]
  assign array_24_io_ve_i = V1_25; // @[SWChisel.scala 197:22]
  assign array_24_io_vf_i = V1_24; // @[SWChisel.scala 199:22]
  assign array_24_io_vv_i = V2_24; // @[SWChisel.scala 200:22]
  assign array_25_io_q = io_q_25_b; // @[SWChisel.scala 220:19]
  assign array_25_io_r = 7'h63 == r_count_25_io_out ? io_r_99_b : _GEN_2748; // @[SWChisel.scala 221:{19,19}]
  assign array_25_io_e_i = E_25; // @[SWChisel.scala 196:21]
  assign array_25_io_f_i = F_25; // @[SWChisel.scala 198:21]
  assign array_25_io_ve_i = V1_26; // @[SWChisel.scala 197:22]
  assign array_25_io_vf_i = V1_25; // @[SWChisel.scala 199:22]
  assign array_25_io_vv_i = V2_25; // @[SWChisel.scala 200:22]
  assign array_26_io_q = io_q_26_b; // @[SWChisel.scala 220:19]
  assign array_26_io_r = 7'h63 == r_count_26_io_out ? io_r_99_b : _GEN_2848; // @[SWChisel.scala 221:{19,19}]
  assign array_26_io_e_i = E_26; // @[SWChisel.scala 196:21]
  assign array_26_io_f_i = F_26; // @[SWChisel.scala 198:21]
  assign array_26_io_ve_i = V1_27; // @[SWChisel.scala 197:22]
  assign array_26_io_vf_i = V1_26; // @[SWChisel.scala 199:22]
  assign array_26_io_vv_i = V2_26; // @[SWChisel.scala 200:22]
  assign array_27_io_q = io_q_27_b; // @[SWChisel.scala 220:19]
  assign array_27_io_r = 7'h63 == r_count_27_io_out ? io_r_99_b : _GEN_2948; // @[SWChisel.scala 221:{19,19}]
  assign array_27_io_e_i = E_27; // @[SWChisel.scala 196:21]
  assign array_27_io_f_i = F_27; // @[SWChisel.scala 198:21]
  assign array_27_io_ve_i = V1_28; // @[SWChisel.scala 197:22]
  assign array_27_io_vf_i = V1_27; // @[SWChisel.scala 199:22]
  assign array_27_io_vv_i = V2_27; // @[SWChisel.scala 200:22]
  assign array_28_io_q = io_q_28_b; // @[SWChisel.scala 220:19]
  assign array_28_io_r = 7'h63 == r_count_28_io_out ? io_r_99_b : _GEN_3048; // @[SWChisel.scala 221:{19,19}]
  assign array_28_io_e_i = E_28; // @[SWChisel.scala 196:21]
  assign array_28_io_f_i = F_28; // @[SWChisel.scala 198:21]
  assign array_28_io_ve_i = V1_29; // @[SWChisel.scala 197:22]
  assign array_28_io_vf_i = V1_28; // @[SWChisel.scala 199:22]
  assign array_28_io_vv_i = V2_28; // @[SWChisel.scala 200:22]
  assign array_29_io_q = io_q_29_b; // @[SWChisel.scala 220:19]
  assign array_29_io_r = 7'h63 == r_count_29_io_out ? io_r_99_b : _GEN_3148; // @[SWChisel.scala 221:{19,19}]
  assign array_29_io_e_i = E_29; // @[SWChisel.scala 196:21]
  assign array_29_io_f_i = F_29; // @[SWChisel.scala 198:21]
  assign array_29_io_ve_i = V1_30; // @[SWChisel.scala 197:22]
  assign array_29_io_vf_i = V1_29; // @[SWChisel.scala 199:22]
  assign array_29_io_vv_i = V2_29; // @[SWChisel.scala 200:22]
  assign array_30_io_q = io_q_30_b; // @[SWChisel.scala 220:19]
  assign array_30_io_r = 7'h63 == r_count_30_io_out ? io_r_99_b : _GEN_3248; // @[SWChisel.scala 221:{19,19}]
  assign array_30_io_e_i = E_30; // @[SWChisel.scala 196:21]
  assign array_30_io_f_i = F_30; // @[SWChisel.scala 198:21]
  assign array_30_io_ve_i = V1_31; // @[SWChisel.scala 197:22]
  assign array_30_io_vf_i = V1_30; // @[SWChisel.scala 199:22]
  assign array_30_io_vv_i = V2_30; // @[SWChisel.scala 200:22]
  assign array_31_io_q = io_q_31_b; // @[SWChisel.scala 220:19]
  assign array_31_io_r = 7'h63 == r_count_31_io_out ? io_r_99_b : _GEN_3348; // @[SWChisel.scala 221:{19,19}]
  assign array_31_io_e_i = E_31; // @[SWChisel.scala 196:21]
  assign array_31_io_f_i = F_31; // @[SWChisel.scala 198:21]
  assign array_31_io_ve_i = V1_32; // @[SWChisel.scala 197:22]
  assign array_31_io_vf_i = V1_31; // @[SWChisel.scala 199:22]
  assign array_31_io_vv_i = V2_31; // @[SWChisel.scala 200:22]
  assign array_32_io_q = io_q_32_b; // @[SWChisel.scala 220:19]
  assign array_32_io_r = 7'h63 == r_count_32_io_out ? io_r_99_b : _GEN_3448; // @[SWChisel.scala 221:{19,19}]
  assign array_32_io_e_i = E_32; // @[SWChisel.scala 196:21]
  assign array_32_io_f_i = F_32; // @[SWChisel.scala 198:21]
  assign array_32_io_ve_i = V1_33; // @[SWChisel.scala 197:22]
  assign array_32_io_vf_i = V1_32; // @[SWChisel.scala 199:22]
  assign array_32_io_vv_i = V2_32; // @[SWChisel.scala 200:22]
  assign array_33_io_q = io_q_33_b; // @[SWChisel.scala 220:19]
  assign array_33_io_r = 7'h63 == r_count_33_io_out ? io_r_99_b : _GEN_3548; // @[SWChisel.scala 221:{19,19}]
  assign array_33_io_e_i = E_33; // @[SWChisel.scala 196:21]
  assign array_33_io_f_i = F_33; // @[SWChisel.scala 198:21]
  assign array_33_io_ve_i = V1_34; // @[SWChisel.scala 197:22]
  assign array_33_io_vf_i = V1_33; // @[SWChisel.scala 199:22]
  assign array_33_io_vv_i = V2_33; // @[SWChisel.scala 200:22]
  assign array_34_io_q = io_q_34_b; // @[SWChisel.scala 220:19]
  assign array_34_io_r = 7'h63 == r_count_34_io_out ? io_r_99_b : _GEN_3648; // @[SWChisel.scala 221:{19,19}]
  assign array_34_io_e_i = E_34; // @[SWChisel.scala 196:21]
  assign array_34_io_f_i = F_34; // @[SWChisel.scala 198:21]
  assign array_34_io_ve_i = V1_35; // @[SWChisel.scala 197:22]
  assign array_34_io_vf_i = V1_34; // @[SWChisel.scala 199:22]
  assign array_34_io_vv_i = V2_34; // @[SWChisel.scala 200:22]
  assign array_35_io_q = io_q_35_b; // @[SWChisel.scala 220:19]
  assign array_35_io_r = 7'h63 == r_count_35_io_out ? io_r_99_b : _GEN_3748; // @[SWChisel.scala 221:{19,19}]
  assign array_35_io_e_i = E_35; // @[SWChisel.scala 196:21]
  assign array_35_io_f_i = F_35; // @[SWChisel.scala 198:21]
  assign array_35_io_ve_i = V1_36; // @[SWChisel.scala 197:22]
  assign array_35_io_vf_i = V1_35; // @[SWChisel.scala 199:22]
  assign array_35_io_vv_i = V2_35; // @[SWChisel.scala 200:22]
  assign array_36_io_q = io_q_36_b; // @[SWChisel.scala 220:19]
  assign array_36_io_r = 7'h63 == r_count_36_io_out ? io_r_99_b : _GEN_3848; // @[SWChisel.scala 221:{19,19}]
  assign array_36_io_e_i = E_36; // @[SWChisel.scala 196:21]
  assign array_36_io_f_i = F_36; // @[SWChisel.scala 198:21]
  assign array_36_io_ve_i = V1_37; // @[SWChisel.scala 197:22]
  assign array_36_io_vf_i = V1_36; // @[SWChisel.scala 199:22]
  assign array_36_io_vv_i = V2_36; // @[SWChisel.scala 200:22]
  assign array_37_io_q = io_q_37_b; // @[SWChisel.scala 220:19]
  assign array_37_io_r = 7'h63 == r_count_37_io_out ? io_r_99_b : _GEN_3948; // @[SWChisel.scala 221:{19,19}]
  assign array_37_io_e_i = E_37; // @[SWChisel.scala 196:21]
  assign array_37_io_f_i = F_37; // @[SWChisel.scala 198:21]
  assign array_37_io_ve_i = V1_38; // @[SWChisel.scala 197:22]
  assign array_37_io_vf_i = V1_37; // @[SWChisel.scala 199:22]
  assign array_37_io_vv_i = V2_37; // @[SWChisel.scala 200:22]
  assign array_38_io_q = io_q_38_b; // @[SWChisel.scala 220:19]
  assign array_38_io_r = 7'h63 == r_count_38_io_out ? io_r_99_b : _GEN_4048; // @[SWChisel.scala 221:{19,19}]
  assign array_38_io_e_i = E_38; // @[SWChisel.scala 196:21]
  assign array_38_io_f_i = F_38; // @[SWChisel.scala 198:21]
  assign array_38_io_ve_i = V1_39; // @[SWChisel.scala 197:22]
  assign array_38_io_vf_i = V1_38; // @[SWChisel.scala 199:22]
  assign array_38_io_vv_i = V2_38; // @[SWChisel.scala 200:22]
  assign array_39_io_q = io_q_39_b; // @[SWChisel.scala 220:19]
  assign array_39_io_r = 7'h63 == r_count_39_io_out ? io_r_99_b : _GEN_4148; // @[SWChisel.scala 221:{19,19}]
  assign array_39_io_e_i = E_39; // @[SWChisel.scala 196:21]
  assign array_39_io_f_i = F_39; // @[SWChisel.scala 198:21]
  assign array_39_io_ve_i = V1_40; // @[SWChisel.scala 197:22]
  assign array_39_io_vf_i = V1_39; // @[SWChisel.scala 199:22]
  assign array_39_io_vv_i = V2_39; // @[SWChisel.scala 200:22]
  assign array_40_io_q = io_q_40_b; // @[SWChisel.scala 220:19]
  assign array_40_io_r = 7'h63 == r_count_40_io_out ? io_r_99_b : _GEN_4248; // @[SWChisel.scala 221:{19,19}]
  assign array_40_io_e_i = E_40; // @[SWChisel.scala 196:21]
  assign array_40_io_f_i = F_40; // @[SWChisel.scala 198:21]
  assign array_40_io_ve_i = V1_41; // @[SWChisel.scala 197:22]
  assign array_40_io_vf_i = V1_40; // @[SWChisel.scala 199:22]
  assign array_40_io_vv_i = V2_40; // @[SWChisel.scala 200:22]
  assign array_41_io_q = io_q_41_b; // @[SWChisel.scala 220:19]
  assign array_41_io_r = 7'h63 == r_count_41_io_out ? io_r_99_b : _GEN_4348; // @[SWChisel.scala 221:{19,19}]
  assign array_41_io_e_i = E_41; // @[SWChisel.scala 196:21]
  assign array_41_io_f_i = F_41; // @[SWChisel.scala 198:21]
  assign array_41_io_ve_i = V1_42; // @[SWChisel.scala 197:22]
  assign array_41_io_vf_i = V1_41; // @[SWChisel.scala 199:22]
  assign array_41_io_vv_i = V2_41; // @[SWChisel.scala 200:22]
  assign array_42_io_q = io_q_42_b; // @[SWChisel.scala 220:19]
  assign array_42_io_r = 7'h63 == r_count_42_io_out ? io_r_99_b : _GEN_4448; // @[SWChisel.scala 221:{19,19}]
  assign array_42_io_e_i = E_42; // @[SWChisel.scala 196:21]
  assign array_42_io_f_i = F_42; // @[SWChisel.scala 198:21]
  assign array_42_io_ve_i = V1_43; // @[SWChisel.scala 197:22]
  assign array_42_io_vf_i = V1_42; // @[SWChisel.scala 199:22]
  assign array_42_io_vv_i = V2_42; // @[SWChisel.scala 200:22]
  assign array_43_io_q = io_q_43_b; // @[SWChisel.scala 220:19]
  assign array_43_io_r = 7'h63 == r_count_43_io_out ? io_r_99_b : _GEN_4548; // @[SWChisel.scala 221:{19,19}]
  assign array_43_io_e_i = E_43; // @[SWChisel.scala 196:21]
  assign array_43_io_f_i = F_43; // @[SWChisel.scala 198:21]
  assign array_43_io_ve_i = V1_44; // @[SWChisel.scala 197:22]
  assign array_43_io_vf_i = V1_43; // @[SWChisel.scala 199:22]
  assign array_43_io_vv_i = V2_43; // @[SWChisel.scala 200:22]
  assign array_44_io_q = io_q_44_b; // @[SWChisel.scala 220:19]
  assign array_44_io_r = 7'h63 == r_count_44_io_out ? io_r_99_b : _GEN_4648; // @[SWChisel.scala 221:{19,19}]
  assign array_44_io_e_i = E_44; // @[SWChisel.scala 196:21]
  assign array_44_io_f_i = F_44; // @[SWChisel.scala 198:21]
  assign array_44_io_ve_i = V1_45; // @[SWChisel.scala 197:22]
  assign array_44_io_vf_i = V1_44; // @[SWChisel.scala 199:22]
  assign array_44_io_vv_i = V2_44; // @[SWChisel.scala 200:22]
  assign array_45_io_q = io_q_45_b; // @[SWChisel.scala 220:19]
  assign array_45_io_r = 7'h63 == r_count_45_io_out ? io_r_99_b : _GEN_4748; // @[SWChisel.scala 221:{19,19}]
  assign array_45_io_e_i = E_45; // @[SWChisel.scala 196:21]
  assign array_45_io_f_i = F_45; // @[SWChisel.scala 198:21]
  assign array_45_io_ve_i = V1_46; // @[SWChisel.scala 197:22]
  assign array_45_io_vf_i = V1_45; // @[SWChisel.scala 199:22]
  assign array_45_io_vv_i = V2_45; // @[SWChisel.scala 200:22]
  assign array_46_io_q = io_q_46_b; // @[SWChisel.scala 220:19]
  assign array_46_io_r = 7'h63 == r_count_46_io_out ? io_r_99_b : _GEN_4848; // @[SWChisel.scala 221:{19,19}]
  assign array_46_io_e_i = E_46; // @[SWChisel.scala 196:21]
  assign array_46_io_f_i = F_46; // @[SWChisel.scala 198:21]
  assign array_46_io_ve_i = V1_47; // @[SWChisel.scala 197:22]
  assign array_46_io_vf_i = V1_46; // @[SWChisel.scala 199:22]
  assign array_46_io_vv_i = V2_46; // @[SWChisel.scala 200:22]
  assign array_47_io_q = io_q_47_b; // @[SWChisel.scala 220:19]
  assign array_47_io_r = 7'h63 == r_count_47_io_out ? io_r_99_b : _GEN_4948; // @[SWChisel.scala 221:{19,19}]
  assign array_47_io_e_i = E_47; // @[SWChisel.scala 196:21]
  assign array_47_io_f_i = F_47; // @[SWChisel.scala 198:21]
  assign array_47_io_ve_i = V1_48; // @[SWChisel.scala 197:22]
  assign array_47_io_vf_i = V1_47; // @[SWChisel.scala 199:22]
  assign array_47_io_vv_i = V2_47; // @[SWChisel.scala 200:22]
  assign array_48_io_q = io_q_48_b; // @[SWChisel.scala 220:19]
  assign array_48_io_r = 7'h63 == r_count_48_io_out ? io_r_99_b : _GEN_5048; // @[SWChisel.scala 221:{19,19}]
  assign array_48_io_e_i = E_48; // @[SWChisel.scala 196:21]
  assign array_48_io_f_i = F_48; // @[SWChisel.scala 198:21]
  assign array_48_io_ve_i = V1_49; // @[SWChisel.scala 197:22]
  assign array_48_io_vf_i = V1_48; // @[SWChisel.scala 199:22]
  assign array_48_io_vv_i = V2_48; // @[SWChisel.scala 200:22]
  assign array_49_io_q = io_q_49_b; // @[SWChisel.scala 220:19]
  assign array_49_io_r = 7'h63 == r_count_49_io_out ? io_r_99_b : _GEN_5148; // @[SWChisel.scala 221:{19,19}]
  assign array_49_io_e_i = E_49; // @[SWChisel.scala 196:21]
  assign array_49_io_f_i = F_49; // @[SWChisel.scala 198:21]
  assign array_49_io_ve_i = V1_50; // @[SWChisel.scala 197:22]
  assign array_49_io_vf_i = V1_49; // @[SWChisel.scala 199:22]
  assign array_49_io_vv_i = V2_49; // @[SWChisel.scala 200:22]
  assign r_count_0_clock = clock;
  assign r_count_0_reset = reset;
  assign r_count_0_io_en = start_reg_0; // @[SWChisel.scala 192:22]
  assign r_count_1_clock = clock;
  assign r_count_1_reset = reset;
  assign r_count_1_io_en = start_reg_1; // @[SWChisel.scala 192:22]
  assign r_count_2_clock = clock;
  assign r_count_2_reset = reset;
  assign r_count_2_io_en = start_reg_2; // @[SWChisel.scala 192:22]
  assign r_count_3_clock = clock;
  assign r_count_3_reset = reset;
  assign r_count_3_io_en = start_reg_3; // @[SWChisel.scala 192:22]
  assign r_count_4_clock = clock;
  assign r_count_4_reset = reset;
  assign r_count_4_io_en = start_reg_4; // @[SWChisel.scala 192:22]
  assign r_count_5_clock = clock;
  assign r_count_5_reset = reset;
  assign r_count_5_io_en = start_reg_5; // @[SWChisel.scala 192:22]
  assign r_count_6_clock = clock;
  assign r_count_6_reset = reset;
  assign r_count_6_io_en = start_reg_6; // @[SWChisel.scala 192:22]
  assign r_count_7_clock = clock;
  assign r_count_7_reset = reset;
  assign r_count_7_io_en = start_reg_7; // @[SWChisel.scala 192:22]
  assign r_count_8_clock = clock;
  assign r_count_8_reset = reset;
  assign r_count_8_io_en = start_reg_8; // @[SWChisel.scala 192:22]
  assign r_count_9_clock = clock;
  assign r_count_9_reset = reset;
  assign r_count_9_io_en = start_reg_9; // @[SWChisel.scala 192:22]
  assign r_count_10_clock = clock;
  assign r_count_10_reset = reset;
  assign r_count_10_io_en = start_reg_10; // @[SWChisel.scala 192:22]
  assign r_count_11_clock = clock;
  assign r_count_11_reset = reset;
  assign r_count_11_io_en = start_reg_11; // @[SWChisel.scala 192:22]
  assign r_count_12_clock = clock;
  assign r_count_12_reset = reset;
  assign r_count_12_io_en = start_reg_12; // @[SWChisel.scala 192:22]
  assign r_count_13_clock = clock;
  assign r_count_13_reset = reset;
  assign r_count_13_io_en = start_reg_13; // @[SWChisel.scala 192:22]
  assign r_count_14_clock = clock;
  assign r_count_14_reset = reset;
  assign r_count_14_io_en = start_reg_14; // @[SWChisel.scala 192:22]
  assign r_count_15_clock = clock;
  assign r_count_15_reset = reset;
  assign r_count_15_io_en = start_reg_15; // @[SWChisel.scala 192:22]
  assign r_count_16_clock = clock;
  assign r_count_16_reset = reset;
  assign r_count_16_io_en = start_reg_16; // @[SWChisel.scala 192:22]
  assign r_count_17_clock = clock;
  assign r_count_17_reset = reset;
  assign r_count_17_io_en = start_reg_17; // @[SWChisel.scala 192:22]
  assign r_count_18_clock = clock;
  assign r_count_18_reset = reset;
  assign r_count_18_io_en = start_reg_18; // @[SWChisel.scala 192:22]
  assign r_count_19_clock = clock;
  assign r_count_19_reset = reset;
  assign r_count_19_io_en = start_reg_19; // @[SWChisel.scala 192:22]
  assign r_count_20_clock = clock;
  assign r_count_20_reset = reset;
  assign r_count_20_io_en = start_reg_20; // @[SWChisel.scala 192:22]
  assign r_count_21_clock = clock;
  assign r_count_21_reset = reset;
  assign r_count_21_io_en = start_reg_21; // @[SWChisel.scala 192:22]
  assign r_count_22_clock = clock;
  assign r_count_22_reset = reset;
  assign r_count_22_io_en = start_reg_22; // @[SWChisel.scala 192:22]
  assign r_count_23_clock = clock;
  assign r_count_23_reset = reset;
  assign r_count_23_io_en = start_reg_23; // @[SWChisel.scala 192:22]
  assign r_count_24_clock = clock;
  assign r_count_24_reset = reset;
  assign r_count_24_io_en = start_reg_24; // @[SWChisel.scala 192:22]
  assign r_count_25_clock = clock;
  assign r_count_25_reset = reset;
  assign r_count_25_io_en = start_reg_25; // @[SWChisel.scala 192:22]
  assign r_count_26_clock = clock;
  assign r_count_26_reset = reset;
  assign r_count_26_io_en = start_reg_26; // @[SWChisel.scala 192:22]
  assign r_count_27_clock = clock;
  assign r_count_27_reset = reset;
  assign r_count_27_io_en = start_reg_27; // @[SWChisel.scala 192:22]
  assign r_count_28_clock = clock;
  assign r_count_28_reset = reset;
  assign r_count_28_io_en = start_reg_28; // @[SWChisel.scala 192:22]
  assign r_count_29_clock = clock;
  assign r_count_29_reset = reset;
  assign r_count_29_io_en = start_reg_29; // @[SWChisel.scala 192:22]
  assign r_count_30_clock = clock;
  assign r_count_30_reset = reset;
  assign r_count_30_io_en = start_reg_30; // @[SWChisel.scala 192:22]
  assign r_count_31_clock = clock;
  assign r_count_31_reset = reset;
  assign r_count_31_io_en = start_reg_31; // @[SWChisel.scala 192:22]
  assign r_count_32_clock = clock;
  assign r_count_32_reset = reset;
  assign r_count_32_io_en = start_reg_32; // @[SWChisel.scala 192:22]
  assign r_count_33_clock = clock;
  assign r_count_33_reset = reset;
  assign r_count_33_io_en = start_reg_33; // @[SWChisel.scala 192:22]
  assign r_count_34_clock = clock;
  assign r_count_34_reset = reset;
  assign r_count_34_io_en = start_reg_34; // @[SWChisel.scala 192:22]
  assign r_count_35_clock = clock;
  assign r_count_35_reset = reset;
  assign r_count_35_io_en = start_reg_35; // @[SWChisel.scala 192:22]
  assign r_count_36_clock = clock;
  assign r_count_36_reset = reset;
  assign r_count_36_io_en = start_reg_36; // @[SWChisel.scala 192:22]
  assign r_count_37_clock = clock;
  assign r_count_37_reset = reset;
  assign r_count_37_io_en = start_reg_37; // @[SWChisel.scala 192:22]
  assign r_count_38_clock = clock;
  assign r_count_38_reset = reset;
  assign r_count_38_io_en = start_reg_38; // @[SWChisel.scala 192:22]
  assign r_count_39_clock = clock;
  assign r_count_39_reset = reset;
  assign r_count_39_io_en = start_reg_39; // @[SWChisel.scala 192:22]
  assign r_count_40_clock = clock;
  assign r_count_40_reset = reset;
  assign r_count_40_io_en = start_reg_40; // @[SWChisel.scala 192:22]
  assign r_count_41_clock = clock;
  assign r_count_41_reset = reset;
  assign r_count_41_io_en = start_reg_41; // @[SWChisel.scala 192:22]
  assign r_count_42_clock = clock;
  assign r_count_42_reset = reset;
  assign r_count_42_io_en = start_reg_42; // @[SWChisel.scala 192:22]
  assign r_count_43_clock = clock;
  assign r_count_43_reset = reset;
  assign r_count_43_io_en = start_reg_43; // @[SWChisel.scala 192:22]
  assign r_count_44_clock = clock;
  assign r_count_44_reset = reset;
  assign r_count_44_io_en = start_reg_44; // @[SWChisel.scala 192:22]
  assign r_count_45_clock = clock;
  assign r_count_45_reset = reset;
  assign r_count_45_io_en = start_reg_45; // @[SWChisel.scala 192:22]
  assign r_count_46_clock = clock;
  assign r_count_46_reset = reset;
  assign r_count_46_io_en = start_reg_46; // @[SWChisel.scala 192:22]
  assign r_count_47_clock = clock;
  assign r_count_47_reset = reset;
  assign r_count_47_io_en = start_reg_47; // @[SWChisel.scala 192:22]
  assign r_count_48_clock = clock;
  assign r_count_48_reset = reset;
  assign r_count_48_io_en = start_reg_48; // @[SWChisel.scala 192:22]
  assign r_count_49_clock = clock;
  assign r_count_49_reset = reset;
  assign r_count_49_io_en = start_reg_49; // @[SWChisel.scala 192:22]
  assign max_clock = clock;
  assign max_reset = reset;
  assign max_io_start = start_reg_49; // @[SWChisel.scala 178:16]
  assign max_io_in = V1_50; // @[SWChisel.scala 177:13]
  always @(posedge clock) begin
    if (reset) begin // @[SWChisel.scala 162:18]
      E_0 <= -16'sh2; // @[SWChisel.scala 162:18]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      E_0 <= array_0_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_1 <= -16'sh3; // @[SWChisel.scala 162:18]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      E_1 <= array_1_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_2 <= -16'sh4; // @[SWChisel.scala 162:18]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      E_2 <= array_2_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_3 <= -16'sh5; // @[SWChisel.scala 162:18]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      E_3 <= array_3_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_4 <= -16'sh6; // @[SWChisel.scala 162:18]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      E_4 <= array_4_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_5 <= -16'sh7; // @[SWChisel.scala 162:18]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      E_5 <= array_5_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_6 <= -16'sh8; // @[SWChisel.scala 162:18]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      E_6 <= array_6_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_7 <= -16'sh9; // @[SWChisel.scala 162:18]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      E_7 <= array_7_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_8 <= -16'sha; // @[SWChisel.scala 162:18]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      E_8 <= array_8_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_9 <= -16'shb; // @[SWChisel.scala 162:18]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      E_9 <= array_9_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_10 <= -16'shc; // @[SWChisel.scala 162:18]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      E_10 <= array_10_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_11 <= -16'shd; // @[SWChisel.scala 162:18]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      E_11 <= array_11_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_12 <= -16'she; // @[SWChisel.scala 162:18]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      E_12 <= array_12_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_13 <= -16'shf; // @[SWChisel.scala 162:18]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      E_13 <= array_13_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_14 <= -16'sh10; // @[SWChisel.scala 162:18]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      E_14 <= array_14_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_15 <= -16'sh11; // @[SWChisel.scala 162:18]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      E_15 <= array_15_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_16 <= -16'sh12; // @[SWChisel.scala 162:18]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      E_16 <= array_16_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_17 <= -16'sh13; // @[SWChisel.scala 162:18]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      E_17 <= array_17_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_18 <= -16'sh14; // @[SWChisel.scala 162:18]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      E_18 <= array_18_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_19 <= -16'sh15; // @[SWChisel.scala 162:18]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      E_19 <= array_19_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_20 <= -16'sh16; // @[SWChisel.scala 162:18]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      E_20 <= array_20_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_21 <= -16'sh17; // @[SWChisel.scala 162:18]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      E_21 <= array_21_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_22 <= -16'sh18; // @[SWChisel.scala 162:18]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      E_22 <= array_22_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_23 <= -16'sh19; // @[SWChisel.scala 162:18]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      E_23 <= array_23_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_24 <= -16'sh1a; // @[SWChisel.scala 162:18]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      E_24 <= array_24_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_25 <= -16'sh1b; // @[SWChisel.scala 162:18]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      E_25 <= array_25_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_26 <= -16'sh1c; // @[SWChisel.scala 162:18]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      E_26 <= array_26_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_27 <= -16'sh1d; // @[SWChisel.scala 162:18]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      E_27 <= array_27_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_28 <= -16'sh1e; // @[SWChisel.scala 162:18]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      E_28 <= array_28_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_29 <= -16'sh1f; // @[SWChisel.scala 162:18]
    end else if (start_reg_29) begin // @[SWChisel.scala 207:25]
      E_29 <= array_29_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_30 <= -16'sh20; // @[SWChisel.scala 162:18]
    end else if (start_reg_30) begin // @[SWChisel.scala 207:25]
      E_30 <= array_30_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_31 <= -16'sh21; // @[SWChisel.scala 162:18]
    end else if (start_reg_31) begin // @[SWChisel.scala 207:25]
      E_31 <= array_31_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_32 <= -16'sh22; // @[SWChisel.scala 162:18]
    end else if (start_reg_32) begin // @[SWChisel.scala 207:25]
      E_32 <= array_32_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_33 <= -16'sh23; // @[SWChisel.scala 162:18]
    end else if (start_reg_33) begin // @[SWChisel.scala 207:25]
      E_33 <= array_33_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_34 <= -16'sh24; // @[SWChisel.scala 162:18]
    end else if (start_reg_34) begin // @[SWChisel.scala 207:25]
      E_34 <= array_34_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_35 <= -16'sh25; // @[SWChisel.scala 162:18]
    end else if (start_reg_35) begin // @[SWChisel.scala 207:25]
      E_35 <= array_35_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_36 <= -16'sh26; // @[SWChisel.scala 162:18]
    end else if (start_reg_36) begin // @[SWChisel.scala 207:25]
      E_36 <= array_36_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_37 <= -16'sh27; // @[SWChisel.scala 162:18]
    end else if (start_reg_37) begin // @[SWChisel.scala 207:25]
      E_37 <= array_37_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_38 <= -16'sh28; // @[SWChisel.scala 162:18]
    end else if (start_reg_38) begin // @[SWChisel.scala 207:25]
      E_38 <= array_38_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_39 <= -16'sh29; // @[SWChisel.scala 162:18]
    end else if (start_reg_39) begin // @[SWChisel.scala 207:25]
      E_39 <= array_39_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_40 <= -16'sh2a; // @[SWChisel.scala 162:18]
    end else if (start_reg_40) begin // @[SWChisel.scala 207:25]
      E_40 <= array_40_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_41 <= -16'sh2b; // @[SWChisel.scala 162:18]
    end else if (start_reg_41) begin // @[SWChisel.scala 207:25]
      E_41 <= array_41_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_42 <= -16'sh2c; // @[SWChisel.scala 162:18]
    end else if (start_reg_42) begin // @[SWChisel.scala 207:25]
      E_42 <= array_42_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_43 <= -16'sh2d; // @[SWChisel.scala 162:18]
    end else if (start_reg_43) begin // @[SWChisel.scala 207:25]
      E_43 <= array_43_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_44 <= -16'sh2e; // @[SWChisel.scala 162:18]
    end else if (start_reg_44) begin // @[SWChisel.scala 207:25]
      E_44 <= array_44_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_45 <= -16'sh2f; // @[SWChisel.scala 162:18]
    end else if (start_reg_45) begin // @[SWChisel.scala 207:25]
      E_45 <= array_45_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_46 <= -16'sh30; // @[SWChisel.scala 162:18]
    end else if (start_reg_46) begin // @[SWChisel.scala 207:25]
      E_46 <= array_46_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_47 <= -16'sh31; // @[SWChisel.scala 162:18]
    end else if (start_reg_47) begin // @[SWChisel.scala 207:25]
      E_47 <= array_47_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_48 <= -16'sh32; // @[SWChisel.scala 162:18]
    end else if (start_reg_48) begin // @[SWChisel.scala 207:25]
      E_48 <= array_48_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_49 <= -16'sh33; // @[SWChisel.scala 162:18]
    end else if (start_reg_49) begin // @[SWChisel.scala 207:25]
      E_49 <= array_49_io_e_o; // @[SWChisel.scala 208:12]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_1 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      F_1 <= array_0_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_2 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      F_2 <= array_1_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_3 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      F_3 <= array_2_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_4 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      F_4 <= array_3_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_5 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      F_5 <= array_4_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_6 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      F_6 <= array_5_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_7 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      F_7 <= array_6_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_8 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      F_8 <= array_7_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_9 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      F_9 <= array_8_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_10 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      F_10 <= array_9_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_11 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      F_11 <= array_10_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_12 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      F_12 <= array_11_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_13 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      F_13 <= array_12_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_14 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      F_14 <= array_13_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_15 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      F_15 <= array_14_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_16 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      F_16 <= array_15_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_17 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      F_17 <= array_16_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_18 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      F_18 <= array_17_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_19 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      F_19 <= array_18_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_20 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      F_20 <= array_19_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_21 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      F_21 <= array_20_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_22 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      F_22 <= array_21_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_23 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      F_23 <= array_22_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_24 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      F_24 <= array_23_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_25 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      F_25 <= array_24_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_26 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      F_26 <= array_25_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_27 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      F_27 <= array_26_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_28 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      F_28 <= array_27_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_29 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      F_29 <= array_28_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_30 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_29) begin // @[SWChisel.scala 207:25]
      F_30 <= array_29_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_31 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_30) begin // @[SWChisel.scala 207:25]
      F_31 <= array_30_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_32 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_31) begin // @[SWChisel.scala 207:25]
      F_32 <= array_31_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_33 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_32) begin // @[SWChisel.scala 207:25]
      F_33 <= array_32_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_34 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_33) begin // @[SWChisel.scala 207:25]
      F_34 <= array_33_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_35 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_34) begin // @[SWChisel.scala 207:25]
      F_35 <= array_34_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_36 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_35) begin // @[SWChisel.scala 207:25]
      F_36 <= array_35_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_37 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_36) begin // @[SWChisel.scala 207:25]
      F_37 <= array_36_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_38 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_37) begin // @[SWChisel.scala 207:25]
      F_38 <= array_37_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_39 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_38) begin // @[SWChisel.scala 207:25]
      F_39 <= array_38_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_40 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_39) begin // @[SWChisel.scala 207:25]
      F_40 <= array_39_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_41 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_40) begin // @[SWChisel.scala 207:25]
      F_41 <= array_40_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_42 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_41) begin // @[SWChisel.scala 207:25]
      F_42 <= array_41_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_43 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_42) begin // @[SWChisel.scala 207:25]
      F_43 <= array_42_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_44 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_43) begin // @[SWChisel.scala 207:25]
      F_44 <= array_43_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_45 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_44) begin // @[SWChisel.scala 207:25]
      F_45 <= array_44_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_46 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_45) begin // @[SWChisel.scala 207:25]
      F_46 <= array_45_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_47 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_46) begin // @[SWChisel.scala 207:25]
      F_47 <= array_46_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_48 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_47) begin // @[SWChisel.scala 207:25]
      F_48 <= array_47_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_49 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_48) begin // @[SWChisel.scala 207:25]
      F_49 <= array_48_io_f_o; // @[SWChisel.scala 209:14]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_0 <= -16'sh1; // @[SWChisel.scala 164:19]
    end else begin
      V1_0 <= 16'sh0; // @[SWChisel.scala 165:9]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_1 <= -16'sh2; // @[SWChisel.scala 164:19]
    end else if (start_reg_0) begin // @[SWChisel.scala 207:25]
      V1_1 <= array_0_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_2 <= -16'sh3; // @[SWChisel.scala 164:19]
    end else if (start_reg_1) begin // @[SWChisel.scala 207:25]
      V1_2 <= array_1_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_3 <= -16'sh4; // @[SWChisel.scala 164:19]
    end else if (start_reg_2) begin // @[SWChisel.scala 207:25]
      V1_3 <= array_2_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_4 <= -16'sh5; // @[SWChisel.scala 164:19]
    end else if (start_reg_3) begin // @[SWChisel.scala 207:25]
      V1_4 <= array_3_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_5 <= -16'sh6; // @[SWChisel.scala 164:19]
    end else if (start_reg_4) begin // @[SWChisel.scala 207:25]
      V1_5 <= array_4_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_6 <= -16'sh7; // @[SWChisel.scala 164:19]
    end else if (start_reg_5) begin // @[SWChisel.scala 207:25]
      V1_6 <= array_5_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_7 <= -16'sh8; // @[SWChisel.scala 164:19]
    end else if (start_reg_6) begin // @[SWChisel.scala 207:25]
      V1_7 <= array_6_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_8 <= -16'sh9; // @[SWChisel.scala 164:19]
    end else if (start_reg_7) begin // @[SWChisel.scala 207:25]
      V1_8 <= array_7_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_9 <= -16'sha; // @[SWChisel.scala 164:19]
    end else if (start_reg_8) begin // @[SWChisel.scala 207:25]
      V1_9 <= array_8_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_10 <= -16'shb; // @[SWChisel.scala 164:19]
    end else if (start_reg_9) begin // @[SWChisel.scala 207:25]
      V1_10 <= array_9_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_11 <= -16'shc; // @[SWChisel.scala 164:19]
    end else if (start_reg_10) begin // @[SWChisel.scala 207:25]
      V1_11 <= array_10_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_12 <= -16'shd; // @[SWChisel.scala 164:19]
    end else if (start_reg_11) begin // @[SWChisel.scala 207:25]
      V1_12 <= array_11_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_13 <= -16'she; // @[SWChisel.scala 164:19]
    end else if (start_reg_12) begin // @[SWChisel.scala 207:25]
      V1_13 <= array_12_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_14 <= -16'shf; // @[SWChisel.scala 164:19]
    end else if (start_reg_13) begin // @[SWChisel.scala 207:25]
      V1_14 <= array_13_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_15 <= -16'sh10; // @[SWChisel.scala 164:19]
    end else if (start_reg_14) begin // @[SWChisel.scala 207:25]
      V1_15 <= array_14_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_16 <= -16'sh11; // @[SWChisel.scala 164:19]
    end else if (start_reg_15) begin // @[SWChisel.scala 207:25]
      V1_16 <= array_15_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_17 <= -16'sh12; // @[SWChisel.scala 164:19]
    end else if (start_reg_16) begin // @[SWChisel.scala 207:25]
      V1_17 <= array_16_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_18 <= -16'sh13; // @[SWChisel.scala 164:19]
    end else if (start_reg_17) begin // @[SWChisel.scala 207:25]
      V1_18 <= array_17_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_19 <= -16'sh14; // @[SWChisel.scala 164:19]
    end else if (start_reg_18) begin // @[SWChisel.scala 207:25]
      V1_19 <= array_18_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_20 <= -16'sh15; // @[SWChisel.scala 164:19]
    end else if (start_reg_19) begin // @[SWChisel.scala 207:25]
      V1_20 <= array_19_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_21 <= -16'sh16; // @[SWChisel.scala 164:19]
    end else if (start_reg_20) begin // @[SWChisel.scala 207:25]
      V1_21 <= array_20_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_22 <= -16'sh17; // @[SWChisel.scala 164:19]
    end else if (start_reg_21) begin // @[SWChisel.scala 207:25]
      V1_22 <= array_21_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_23 <= -16'sh18; // @[SWChisel.scala 164:19]
    end else if (start_reg_22) begin // @[SWChisel.scala 207:25]
      V1_23 <= array_22_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_24 <= -16'sh19; // @[SWChisel.scala 164:19]
    end else if (start_reg_23) begin // @[SWChisel.scala 207:25]
      V1_24 <= array_23_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_25 <= -16'sh1a; // @[SWChisel.scala 164:19]
    end else if (start_reg_24) begin // @[SWChisel.scala 207:25]
      V1_25 <= array_24_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_26 <= -16'sh1b; // @[SWChisel.scala 164:19]
    end else if (start_reg_25) begin // @[SWChisel.scala 207:25]
      V1_26 <= array_25_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_27 <= -16'sh1c; // @[SWChisel.scala 164:19]
    end else if (start_reg_26) begin // @[SWChisel.scala 207:25]
      V1_27 <= array_26_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_28 <= -16'sh1d; // @[SWChisel.scala 164:19]
    end else if (start_reg_27) begin // @[SWChisel.scala 207:25]
      V1_28 <= array_27_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_29 <= -16'sh1e; // @[SWChisel.scala 164:19]
    end else if (start_reg_28) begin // @[SWChisel.scala 207:25]
      V1_29 <= array_28_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_30 <= -16'sh1f; // @[SWChisel.scala 164:19]
    end else if (start_reg_29) begin // @[SWChisel.scala 207:25]
      V1_30 <= array_29_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_31 <= -16'sh20; // @[SWChisel.scala 164:19]
    end else if (start_reg_30) begin // @[SWChisel.scala 207:25]
      V1_31 <= array_30_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_32 <= -16'sh21; // @[SWChisel.scala 164:19]
    end else if (start_reg_31) begin // @[SWChisel.scala 207:25]
      V1_32 <= array_31_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_33 <= -16'sh22; // @[SWChisel.scala 164:19]
    end else if (start_reg_32) begin // @[SWChisel.scala 207:25]
      V1_33 <= array_32_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_34 <= -16'sh23; // @[SWChisel.scala 164:19]
    end else if (start_reg_33) begin // @[SWChisel.scala 207:25]
      V1_34 <= array_33_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_35 <= -16'sh24; // @[SWChisel.scala 164:19]
    end else if (start_reg_34) begin // @[SWChisel.scala 207:25]
      V1_35 <= array_34_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_36 <= -16'sh25; // @[SWChisel.scala 164:19]
    end else if (start_reg_35) begin // @[SWChisel.scala 207:25]
      V1_36 <= array_35_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_37 <= -16'sh26; // @[SWChisel.scala 164:19]
    end else if (start_reg_36) begin // @[SWChisel.scala 207:25]
      V1_37 <= array_36_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_38 <= -16'sh27; // @[SWChisel.scala 164:19]
    end else if (start_reg_37) begin // @[SWChisel.scala 207:25]
      V1_38 <= array_37_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_39 <= -16'sh28; // @[SWChisel.scala 164:19]
    end else if (start_reg_38) begin // @[SWChisel.scala 207:25]
      V1_39 <= array_38_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_40 <= -16'sh29; // @[SWChisel.scala 164:19]
    end else if (start_reg_39) begin // @[SWChisel.scala 207:25]
      V1_40 <= array_39_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_41 <= -16'sh2a; // @[SWChisel.scala 164:19]
    end else if (start_reg_40) begin // @[SWChisel.scala 207:25]
      V1_41 <= array_40_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_42 <= -16'sh2b; // @[SWChisel.scala 164:19]
    end else if (start_reg_41) begin // @[SWChisel.scala 207:25]
      V1_42 <= array_41_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_43 <= -16'sh2c; // @[SWChisel.scala 164:19]
    end else if (start_reg_42) begin // @[SWChisel.scala 207:25]
      V1_43 <= array_42_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_44 <= -16'sh2d; // @[SWChisel.scala 164:19]
    end else if (start_reg_43) begin // @[SWChisel.scala 207:25]
      V1_44 <= array_43_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_45 <= -16'sh2e; // @[SWChisel.scala 164:19]
    end else if (start_reg_44) begin // @[SWChisel.scala 207:25]
      V1_45 <= array_44_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_46 <= -16'sh2f; // @[SWChisel.scala 164:19]
    end else if (start_reg_45) begin // @[SWChisel.scala 207:25]
      V1_46 <= array_45_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_47 <= -16'sh30; // @[SWChisel.scala 164:19]
    end else if (start_reg_46) begin // @[SWChisel.scala 207:25]
      V1_47 <= array_46_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_48 <= -16'sh31; // @[SWChisel.scala 164:19]
    end else if (start_reg_47) begin // @[SWChisel.scala 207:25]
      V1_48 <= array_47_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_49 <= -16'sh32; // @[SWChisel.scala 164:19]
    end else if (start_reg_48) begin // @[SWChisel.scala 207:25]
      V1_49 <= array_48_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_50 <= -16'sh33; // @[SWChisel.scala 164:19]
    end else if (start_reg_49) begin // @[SWChisel.scala 207:25]
      V1_50 <= array_49_io_v_o; // @[SWChisel.scala 210:15]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_0 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_0 <= V1_0; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_1 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_1 <= V1_1; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_2 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_2 <= V1_2; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_3 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_3 <= V1_3; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_4 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_4 <= V1_4; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_5 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_5 <= V1_5; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_6 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_6 <= V1_6; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_7 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_7 <= V1_7; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_8 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_8 <= V1_8; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_9 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_9 <= V1_9; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_10 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_10 <= V1_10; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_11 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_11 <= V1_11; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_12 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_12 <= V1_12; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_13 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_13 <= V1_13; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_14 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_14 <= V1_14; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_15 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_15 <= V1_15; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_16 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_16 <= V1_16; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_17 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_17 <= V1_17; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_18 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_18 <= V1_18; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_19 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_19 <= V1_19; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_20 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_20 <= V1_20; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_21 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_21 <= V1_21; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_22 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_22 <= V1_22; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_23 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_23 <= V1_23; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_24 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_24 <= V1_24; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_25 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_25 <= V1_25; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_26 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_26 <= V1_26; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_27 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_27 <= V1_27; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_28 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_28 <= V1_28; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_29 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_29 <= V1_29; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_30 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_30 <= V1_30; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_31 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_31 <= V1_31; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_32 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_32 <= V1_32; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_33 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_33 <= V1_33; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_34 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_34 <= V1_34; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_35 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_35 <= V1_35; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_36 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_36 <= V1_36; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_37 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_37 <= V1_37; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_38 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_38 <= V1_38; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_39 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_39 <= V1_39; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_40 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_40 <= V1_40; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_41 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_41 <= V1_41; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_42 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_42 <= V1_42; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_43 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_43 <= V1_43; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_44 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_44 <= V1_44; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_45 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_45 <= V1_45; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_46 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_46 <= V1_46; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_47 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_47 <= V1_47; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_48 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_48 <= V1_48; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 166:19]
      V2_49 <= 16'sh0; // @[SWChisel.scala 166:19]
    end else begin
      V2_49 <= V1_49; // @[SWChisel.scala 226:11]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_0 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_0 <= io_start; // @[SWChisel.scala 185:16]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_1 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_1 <= start_reg_0; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_2 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_2 <= start_reg_1; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_3 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_3 <= start_reg_2; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_4 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_4 <= start_reg_3; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_5 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_5 <= start_reg_4; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_6 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_6 <= start_reg_5; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_7 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_7 <= start_reg_6; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_8 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_8 <= start_reg_7; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_9 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_9 <= start_reg_8; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_10 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_10 <= start_reg_9; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_11 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_11 <= start_reg_10; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_12 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_12 <= start_reg_11; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_13 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_13 <= start_reg_12; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_14 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_14 <= start_reg_13; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_15 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_15 <= start_reg_14; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_16 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_16 <= start_reg_15; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_17 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_17 <= start_reg_16; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_18 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_18 <= start_reg_17; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_19 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_19 <= start_reg_18; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_20 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_20 <= start_reg_19; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_21 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_21 <= start_reg_20; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_22 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_22 <= start_reg_21; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_23 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_23 <= start_reg_22; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_24 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_24 <= start_reg_23; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_25 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_25 <= start_reg_24; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_26 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_26 <= start_reg_25; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_27 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_27 <= start_reg_26; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_28 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_28 <= start_reg_27; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_29 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_29 <= start_reg_28; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_30 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_30 <= start_reg_29; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_31 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_31 <= start_reg_30; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_32 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_32 <= start_reg_31; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_33 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_33 <= start_reg_32; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_34 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_34 <= start_reg_33; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_35 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_35 <= start_reg_34; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_36 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_36 <= start_reg_35; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_37 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_37 <= start_reg_36; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_38 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_38 <= start_reg_37; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_39 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_39 <= start_reg_38; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_40 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_40 <= start_reg_39; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_41 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_41 <= start_reg_40; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_42 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_42 <= start_reg_41; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_43 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_43 <= start_reg_42; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_44 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_44 <= start_reg_43; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_45 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_45 <= start_reg_44; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_46 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_46 <= start_reg_45; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_47 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_47 <= start_reg_46; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_48 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_48 <= start_reg_47; // @[SWChisel.scala 187:18]
    end
    if (reset) begin // @[SWChisel.scala 167:26]
      start_reg_49 <= 1'h0; // @[SWChisel.scala 167:26]
    end else begin
      start_reg_49 <= start_reg_48; // @[SWChisel.scala 187:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  E_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  E_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  E_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  E_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  E_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  E_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  E_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  E_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  E_8 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  E_9 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  E_10 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  E_11 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  E_12 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  E_13 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  E_14 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  E_15 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  E_16 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  E_17 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  E_18 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  E_19 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  E_20 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  E_21 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  E_22 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  E_23 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  E_24 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  E_25 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  E_26 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  E_27 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  E_28 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  E_29 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  E_30 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  E_31 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  E_32 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  E_33 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  E_34 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  E_35 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  E_36 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  E_37 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  E_38 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  E_39 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  E_40 = _RAND_40[15:0];
  _RAND_41 = {1{`RANDOM}};
  E_41 = _RAND_41[15:0];
  _RAND_42 = {1{`RANDOM}};
  E_42 = _RAND_42[15:0];
  _RAND_43 = {1{`RANDOM}};
  E_43 = _RAND_43[15:0];
  _RAND_44 = {1{`RANDOM}};
  E_44 = _RAND_44[15:0];
  _RAND_45 = {1{`RANDOM}};
  E_45 = _RAND_45[15:0];
  _RAND_46 = {1{`RANDOM}};
  E_46 = _RAND_46[15:0];
  _RAND_47 = {1{`RANDOM}};
  E_47 = _RAND_47[15:0];
  _RAND_48 = {1{`RANDOM}};
  E_48 = _RAND_48[15:0];
  _RAND_49 = {1{`RANDOM}};
  E_49 = _RAND_49[15:0];
  _RAND_50 = {1{`RANDOM}};
  F_1 = _RAND_50[15:0];
  _RAND_51 = {1{`RANDOM}};
  F_2 = _RAND_51[15:0];
  _RAND_52 = {1{`RANDOM}};
  F_3 = _RAND_52[15:0];
  _RAND_53 = {1{`RANDOM}};
  F_4 = _RAND_53[15:0];
  _RAND_54 = {1{`RANDOM}};
  F_5 = _RAND_54[15:0];
  _RAND_55 = {1{`RANDOM}};
  F_6 = _RAND_55[15:0];
  _RAND_56 = {1{`RANDOM}};
  F_7 = _RAND_56[15:0];
  _RAND_57 = {1{`RANDOM}};
  F_8 = _RAND_57[15:0];
  _RAND_58 = {1{`RANDOM}};
  F_9 = _RAND_58[15:0];
  _RAND_59 = {1{`RANDOM}};
  F_10 = _RAND_59[15:0];
  _RAND_60 = {1{`RANDOM}};
  F_11 = _RAND_60[15:0];
  _RAND_61 = {1{`RANDOM}};
  F_12 = _RAND_61[15:0];
  _RAND_62 = {1{`RANDOM}};
  F_13 = _RAND_62[15:0];
  _RAND_63 = {1{`RANDOM}};
  F_14 = _RAND_63[15:0];
  _RAND_64 = {1{`RANDOM}};
  F_15 = _RAND_64[15:0];
  _RAND_65 = {1{`RANDOM}};
  F_16 = _RAND_65[15:0];
  _RAND_66 = {1{`RANDOM}};
  F_17 = _RAND_66[15:0];
  _RAND_67 = {1{`RANDOM}};
  F_18 = _RAND_67[15:0];
  _RAND_68 = {1{`RANDOM}};
  F_19 = _RAND_68[15:0];
  _RAND_69 = {1{`RANDOM}};
  F_20 = _RAND_69[15:0];
  _RAND_70 = {1{`RANDOM}};
  F_21 = _RAND_70[15:0];
  _RAND_71 = {1{`RANDOM}};
  F_22 = _RAND_71[15:0];
  _RAND_72 = {1{`RANDOM}};
  F_23 = _RAND_72[15:0];
  _RAND_73 = {1{`RANDOM}};
  F_24 = _RAND_73[15:0];
  _RAND_74 = {1{`RANDOM}};
  F_25 = _RAND_74[15:0];
  _RAND_75 = {1{`RANDOM}};
  F_26 = _RAND_75[15:0];
  _RAND_76 = {1{`RANDOM}};
  F_27 = _RAND_76[15:0];
  _RAND_77 = {1{`RANDOM}};
  F_28 = _RAND_77[15:0];
  _RAND_78 = {1{`RANDOM}};
  F_29 = _RAND_78[15:0];
  _RAND_79 = {1{`RANDOM}};
  F_30 = _RAND_79[15:0];
  _RAND_80 = {1{`RANDOM}};
  F_31 = _RAND_80[15:0];
  _RAND_81 = {1{`RANDOM}};
  F_32 = _RAND_81[15:0];
  _RAND_82 = {1{`RANDOM}};
  F_33 = _RAND_82[15:0];
  _RAND_83 = {1{`RANDOM}};
  F_34 = _RAND_83[15:0];
  _RAND_84 = {1{`RANDOM}};
  F_35 = _RAND_84[15:0];
  _RAND_85 = {1{`RANDOM}};
  F_36 = _RAND_85[15:0];
  _RAND_86 = {1{`RANDOM}};
  F_37 = _RAND_86[15:0];
  _RAND_87 = {1{`RANDOM}};
  F_38 = _RAND_87[15:0];
  _RAND_88 = {1{`RANDOM}};
  F_39 = _RAND_88[15:0];
  _RAND_89 = {1{`RANDOM}};
  F_40 = _RAND_89[15:0];
  _RAND_90 = {1{`RANDOM}};
  F_41 = _RAND_90[15:0];
  _RAND_91 = {1{`RANDOM}};
  F_42 = _RAND_91[15:0];
  _RAND_92 = {1{`RANDOM}};
  F_43 = _RAND_92[15:0];
  _RAND_93 = {1{`RANDOM}};
  F_44 = _RAND_93[15:0];
  _RAND_94 = {1{`RANDOM}};
  F_45 = _RAND_94[15:0];
  _RAND_95 = {1{`RANDOM}};
  F_46 = _RAND_95[15:0];
  _RAND_96 = {1{`RANDOM}};
  F_47 = _RAND_96[15:0];
  _RAND_97 = {1{`RANDOM}};
  F_48 = _RAND_97[15:0];
  _RAND_98 = {1{`RANDOM}};
  F_49 = _RAND_98[15:0];
  _RAND_99 = {1{`RANDOM}};
  V1_0 = _RAND_99[15:0];
  _RAND_100 = {1{`RANDOM}};
  V1_1 = _RAND_100[15:0];
  _RAND_101 = {1{`RANDOM}};
  V1_2 = _RAND_101[15:0];
  _RAND_102 = {1{`RANDOM}};
  V1_3 = _RAND_102[15:0];
  _RAND_103 = {1{`RANDOM}};
  V1_4 = _RAND_103[15:0];
  _RAND_104 = {1{`RANDOM}};
  V1_5 = _RAND_104[15:0];
  _RAND_105 = {1{`RANDOM}};
  V1_6 = _RAND_105[15:0];
  _RAND_106 = {1{`RANDOM}};
  V1_7 = _RAND_106[15:0];
  _RAND_107 = {1{`RANDOM}};
  V1_8 = _RAND_107[15:0];
  _RAND_108 = {1{`RANDOM}};
  V1_9 = _RAND_108[15:0];
  _RAND_109 = {1{`RANDOM}};
  V1_10 = _RAND_109[15:0];
  _RAND_110 = {1{`RANDOM}};
  V1_11 = _RAND_110[15:0];
  _RAND_111 = {1{`RANDOM}};
  V1_12 = _RAND_111[15:0];
  _RAND_112 = {1{`RANDOM}};
  V1_13 = _RAND_112[15:0];
  _RAND_113 = {1{`RANDOM}};
  V1_14 = _RAND_113[15:0];
  _RAND_114 = {1{`RANDOM}};
  V1_15 = _RAND_114[15:0];
  _RAND_115 = {1{`RANDOM}};
  V1_16 = _RAND_115[15:0];
  _RAND_116 = {1{`RANDOM}};
  V1_17 = _RAND_116[15:0];
  _RAND_117 = {1{`RANDOM}};
  V1_18 = _RAND_117[15:0];
  _RAND_118 = {1{`RANDOM}};
  V1_19 = _RAND_118[15:0];
  _RAND_119 = {1{`RANDOM}};
  V1_20 = _RAND_119[15:0];
  _RAND_120 = {1{`RANDOM}};
  V1_21 = _RAND_120[15:0];
  _RAND_121 = {1{`RANDOM}};
  V1_22 = _RAND_121[15:0];
  _RAND_122 = {1{`RANDOM}};
  V1_23 = _RAND_122[15:0];
  _RAND_123 = {1{`RANDOM}};
  V1_24 = _RAND_123[15:0];
  _RAND_124 = {1{`RANDOM}};
  V1_25 = _RAND_124[15:0];
  _RAND_125 = {1{`RANDOM}};
  V1_26 = _RAND_125[15:0];
  _RAND_126 = {1{`RANDOM}};
  V1_27 = _RAND_126[15:0];
  _RAND_127 = {1{`RANDOM}};
  V1_28 = _RAND_127[15:0];
  _RAND_128 = {1{`RANDOM}};
  V1_29 = _RAND_128[15:0];
  _RAND_129 = {1{`RANDOM}};
  V1_30 = _RAND_129[15:0];
  _RAND_130 = {1{`RANDOM}};
  V1_31 = _RAND_130[15:0];
  _RAND_131 = {1{`RANDOM}};
  V1_32 = _RAND_131[15:0];
  _RAND_132 = {1{`RANDOM}};
  V1_33 = _RAND_132[15:0];
  _RAND_133 = {1{`RANDOM}};
  V1_34 = _RAND_133[15:0];
  _RAND_134 = {1{`RANDOM}};
  V1_35 = _RAND_134[15:0];
  _RAND_135 = {1{`RANDOM}};
  V1_36 = _RAND_135[15:0];
  _RAND_136 = {1{`RANDOM}};
  V1_37 = _RAND_136[15:0];
  _RAND_137 = {1{`RANDOM}};
  V1_38 = _RAND_137[15:0];
  _RAND_138 = {1{`RANDOM}};
  V1_39 = _RAND_138[15:0];
  _RAND_139 = {1{`RANDOM}};
  V1_40 = _RAND_139[15:0];
  _RAND_140 = {1{`RANDOM}};
  V1_41 = _RAND_140[15:0];
  _RAND_141 = {1{`RANDOM}};
  V1_42 = _RAND_141[15:0];
  _RAND_142 = {1{`RANDOM}};
  V1_43 = _RAND_142[15:0];
  _RAND_143 = {1{`RANDOM}};
  V1_44 = _RAND_143[15:0];
  _RAND_144 = {1{`RANDOM}};
  V1_45 = _RAND_144[15:0];
  _RAND_145 = {1{`RANDOM}};
  V1_46 = _RAND_145[15:0];
  _RAND_146 = {1{`RANDOM}};
  V1_47 = _RAND_146[15:0];
  _RAND_147 = {1{`RANDOM}};
  V1_48 = _RAND_147[15:0];
  _RAND_148 = {1{`RANDOM}};
  V1_49 = _RAND_148[15:0];
  _RAND_149 = {1{`RANDOM}};
  V1_50 = _RAND_149[15:0];
  _RAND_150 = {1{`RANDOM}};
  V2_0 = _RAND_150[15:0];
  _RAND_151 = {1{`RANDOM}};
  V2_1 = _RAND_151[15:0];
  _RAND_152 = {1{`RANDOM}};
  V2_2 = _RAND_152[15:0];
  _RAND_153 = {1{`RANDOM}};
  V2_3 = _RAND_153[15:0];
  _RAND_154 = {1{`RANDOM}};
  V2_4 = _RAND_154[15:0];
  _RAND_155 = {1{`RANDOM}};
  V2_5 = _RAND_155[15:0];
  _RAND_156 = {1{`RANDOM}};
  V2_6 = _RAND_156[15:0];
  _RAND_157 = {1{`RANDOM}};
  V2_7 = _RAND_157[15:0];
  _RAND_158 = {1{`RANDOM}};
  V2_8 = _RAND_158[15:0];
  _RAND_159 = {1{`RANDOM}};
  V2_9 = _RAND_159[15:0];
  _RAND_160 = {1{`RANDOM}};
  V2_10 = _RAND_160[15:0];
  _RAND_161 = {1{`RANDOM}};
  V2_11 = _RAND_161[15:0];
  _RAND_162 = {1{`RANDOM}};
  V2_12 = _RAND_162[15:0];
  _RAND_163 = {1{`RANDOM}};
  V2_13 = _RAND_163[15:0];
  _RAND_164 = {1{`RANDOM}};
  V2_14 = _RAND_164[15:0];
  _RAND_165 = {1{`RANDOM}};
  V2_15 = _RAND_165[15:0];
  _RAND_166 = {1{`RANDOM}};
  V2_16 = _RAND_166[15:0];
  _RAND_167 = {1{`RANDOM}};
  V2_17 = _RAND_167[15:0];
  _RAND_168 = {1{`RANDOM}};
  V2_18 = _RAND_168[15:0];
  _RAND_169 = {1{`RANDOM}};
  V2_19 = _RAND_169[15:0];
  _RAND_170 = {1{`RANDOM}};
  V2_20 = _RAND_170[15:0];
  _RAND_171 = {1{`RANDOM}};
  V2_21 = _RAND_171[15:0];
  _RAND_172 = {1{`RANDOM}};
  V2_22 = _RAND_172[15:0];
  _RAND_173 = {1{`RANDOM}};
  V2_23 = _RAND_173[15:0];
  _RAND_174 = {1{`RANDOM}};
  V2_24 = _RAND_174[15:0];
  _RAND_175 = {1{`RANDOM}};
  V2_25 = _RAND_175[15:0];
  _RAND_176 = {1{`RANDOM}};
  V2_26 = _RAND_176[15:0];
  _RAND_177 = {1{`RANDOM}};
  V2_27 = _RAND_177[15:0];
  _RAND_178 = {1{`RANDOM}};
  V2_28 = _RAND_178[15:0];
  _RAND_179 = {1{`RANDOM}};
  V2_29 = _RAND_179[15:0];
  _RAND_180 = {1{`RANDOM}};
  V2_30 = _RAND_180[15:0];
  _RAND_181 = {1{`RANDOM}};
  V2_31 = _RAND_181[15:0];
  _RAND_182 = {1{`RANDOM}};
  V2_32 = _RAND_182[15:0];
  _RAND_183 = {1{`RANDOM}};
  V2_33 = _RAND_183[15:0];
  _RAND_184 = {1{`RANDOM}};
  V2_34 = _RAND_184[15:0];
  _RAND_185 = {1{`RANDOM}};
  V2_35 = _RAND_185[15:0];
  _RAND_186 = {1{`RANDOM}};
  V2_36 = _RAND_186[15:0];
  _RAND_187 = {1{`RANDOM}};
  V2_37 = _RAND_187[15:0];
  _RAND_188 = {1{`RANDOM}};
  V2_38 = _RAND_188[15:0];
  _RAND_189 = {1{`RANDOM}};
  V2_39 = _RAND_189[15:0];
  _RAND_190 = {1{`RANDOM}};
  V2_40 = _RAND_190[15:0];
  _RAND_191 = {1{`RANDOM}};
  V2_41 = _RAND_191[15:0];
  _RAND_192 = {1{`RANDOM}};
  V2_42 = _RAND_192[15:0];
  _RAND_193 = {1{`RANDOM}};
  V2_43 = _RAND_193[15:0];
  _RAND_194 = {1{`RANDOM}};
  V2_44 = _RAND_194[15:0];
  _RAND_195 = {1{`RANDOM}};
  V2_45 = _RAND_195[15:0];
  _RAND_196 = {1{`RANDOM}};
  V2_46 = _RAND_196[15:0];
  _RAND_197 = {1{`RANDOM}};
  V2_47 = _RAND_197[15:0];
  _RAND_198 = {1{`RANDOM}};
  V2_48 = _RAND_198[15:0];
  _RAND_199 = {1{`RANDOM}};
  V2_49 = _RAND_199[15:0];
  _RAND_200 = {1{`RANDOM}};
  start_reg_0 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  start_reg_1 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  start_reg_2 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  start_reg_3 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  start_reg_4 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  start_reg_5 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  start_reg_6 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  start_reg_7 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  start_reg_8 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  start_reg_9 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  start_reg_10 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  start_reg_11 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  start_reg_12 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  start_reg_13 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  start_reg_14 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  start_reg_15 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  start_reg_16 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  start_reg_17 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  start_reg_18 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  start_reg_19 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  start_reg_20 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  start_reg_21 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  start_reg_22 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  start_reg_23 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  start_reg_24 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  start_reg_25 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  start_reg_26 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  start_reg_27 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  start_reg_28 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  start_reg_29 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  start_reg_30 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  start_reg_31 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  start_reg_32 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  start_reg_33 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  start_reg_34 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  start_reg_35 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  start_reg_36 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  start_reg_37 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  start_reg_38 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  start_reg_39 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  start_reg_40 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  start_reg_41 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  start_reg_42 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  start_reg_43 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  start_reg_44 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  start_reg_45 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  start_reg_46 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  start_reg_47 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  start_reg_48 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  start_reg_49 = _RAND_249[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
