/* verilator lint_off DECLFILENAME */
/* verilator lint_off UNUSEDSIGNAL */

module SW(
  input         clock,
  input         reset,
  input  [1:0]  io_q_0_b,
  input  [1:0]  io_q_1_b,
  input  [1:0]  io_q_2_b,
  input  [1:0]  io_q_3_b,
  input  [1:0]  io_q_4_b,
  input  [1:0]  io_q_5_b,
  input  [1:0]  io_q_6_b,
  input  [1:0]  io_q_7_b,
  input  [1:0]  io_q_8_b,
  input  [1:0]  io_q_9_b,
  input  [1:0]  io_r_0_b,
  input  [1:0]  io_r_1_b,
  input  [1:0]  io_r_2_b,
  input  [1:0]  io_r_3_b,
  input  [1:0]  io_r_4_b,
  input  [1:0]  io_r_5_b,
  input  [1:0]  io_r_6_b,
  input  [1:0]  io_r_7_b,
  input  [1:0]  io_r_8_b,
  input  [1:0]  io_r_9_b,
  input  [1:0]  io_r_10_b,
  input  [1:0]  io_r_11_b,
  input  [1:0]  io_r_12_b,
  input  [1:0]  io_r_13_b,
  input  [1:0]  io_r_14_b,
  input  [1:0]  io_r_15_b,
  input  [1:0]  io_r_16_b,
  input         io_start,
  output [15:0] io_result,
  output        io_done,
  output [15:0] io_v1_out_0,
  output [15:0] io_v1_out_1,
  output [15:0] io_v1_out_2,
  output [15:0] io_v1_out_3,
  output [15:0] io_v1_out_4,
  output [15:0] io_v1_out_5,
  output [15:0] io_v1_out_6,
  output [15:0] io_v1_out_7,
  output [15:0] io_v1_out_8,
  output [15:0] io_v1_out_9,
  output [15:0] io_v1_out_10,
  output [15:0] io_v2_out_0,
  output [15:0] io_v2_out_1,
  output [15:0] io_v2_out_2,
  output [15:0] io_v2_out_3,
  output [15:0] io_v2_out_4,
  output [15:0] io_v2_out_5,
  output [15:0] io_v2_out_6,
  output [15:0] io_v2_out_7,
  output [15:0] io_v2_out_8,
  output [15:0] io_v2_out_9,
  output [15:0] io_v2_out_10,
  output [15:0] io_e_out_0,
  output [15:0] io_e_out_1,
  output [15:0] io_e_out_2,
  output [15:0] io_e_out_3,
  output [15:0] io_e_out_4,
  output [15:0] io_e_out_5,
  output [15:0] io_e_out_6,
  output [15:0] io_e_out_7,
  output [15:0] io_e_out_8,
  output [15:0] io_e_out_9,
  output [15:0] io_f_out_0,
  output [15:0] io_f_out_1,
  output [15:0] io_f_out_2,
  output [15:0] io_f_out_3,
  output [15:0] io_f_out_4,
  output [15:0] io_f_out_5,
  output [15:0] io_f_out_6,
  output [15:0] io_f_out_7,
  output [15:0] io_f_out_8,
  output [15:0] io_f_out_9,
  output [15:0] io_f_out_10
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
`endif // RANDOMIZE_REG_INIT
  wire [1:0] array_0_io_q; // @[SWChisel.scala 171:39]
  wire [1:0] array_0_io_r; // @[SWChisel.scala 171:39]
  wire [15:0] array_0_io_e_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_0_io_f_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_0_io_ve_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_0_io_vf_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_0_io_vv_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_0_io_e_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_0_io_f_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_0_io_v_o; // @[SWChisel.scala 171:39]
  wire [1:0] array_1_io_q; // @[SWChisel.scala 171:39]
  wire [1:0] array_1_io_r; // @[SWChisel.scala 171:39]
  wire [15:0] array_1_io_e_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_1_io_f_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_1_io_ve_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_1_io_vf_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_1_io_vv_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_1_io_e_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_1_io_f_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_1_io_v_o; // @[SWChisel.scala 171:39]
  wire [1:0] array_2_io_q; // @[SWChisel.scala 171:39]
  wire [1:0] array_2_io_r; // @[SWChisel.scala 171:39]
  wire [15:0] array_2_io_e_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_2_io_f_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_2_io_ve_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_2_io_vf_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_2_io_vv_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_2_io_e_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_2_io_f_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_2_io_v_o; // @[SWChisel.scala 171:39]
  wire [1:0] array_3_io_q; // @[SWChisel.scala 171:39]
  wire [1:0] array_3_io_r; // @[SWChisel.scala 171:39]
  wire [15:0] array_3_io_e_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_3_io_f_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_3_io_ve_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_3_io_vf_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_3_io_vv_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_3_io_e_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_3_io_f_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_3_io_v_o; // @[SWChisel.scala 171:39]
  wire [1:0] array_4_io_q; // @[SWChisel.scala 171:39]
  wire [1:0] array_4_io_r; // @[SWChisel.scala 171:39]
  wire [15:0] array_4_io_e_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_4_io_f_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_4_io_ve_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_4_io_vf_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_4_io_vv_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_4_io_e_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_4_io_f_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_4_io_v_o; // @[SWChisel.scala 171:39]
  wire [1:0] array_5_io_q; // @[SWChisel.scala 171:39]
  wire [1:0] array_5_io_r; // @[SWChisel.scala 171:39]
  wire [15:0] array_5_io_e_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_5_io_f_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_5_io_ve_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_5_io_vf_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_5_io_vv_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_5_io_e_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_5_io_f_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_5_io_v_o; // @[SWChisel.scala 171:39]
  wire [1:0] array_6_io_q; // @[SWChisel.scala 171:39]
  wire [1:0] array_6_io_r; // @[SWChisel.scala 171:39]
  wire [15:0] array_6_io_e_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_6_io_f_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_6_io_ve_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_6_io_vf_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_6_io_vv_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_6_io_e_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_6_io_f_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_6_io_v_o; // @[SWChisel.scala 171:39]
  wire [1:0] array_7_io_q; // @[SWChisel.scala 171:39]
  wire [1:0] array_7_io_r; // @[SWChisel.scala 171:39]
  wire [15:0] array_7_io_e_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_7_io_f_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_7_io_ve_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_7_io_vf_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_7_io_vv_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_7_io_e_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_7_io_f_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_7_io_v_o; // @[SWChisel.scala 171:39]
  wire [1:0] array_8_io_q; // @[SWChisel.scala 171:39]
  wire [1:0] array_8_io_r; // @[SWChisel.scala 171:39]
  wire [15:0] array_8_io_e_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_8_io_f_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_8_io_ve_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_8_io_vf_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_8_io_vv_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_8_io_e_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_8_io_f_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_8_io_v_o; // @[SWChisel.scala 171:39]
  wire [1:0] array_9_io_q; // @[SWChisel.scala 171:39]
  wire [1:0] array_9_io_r; // @[SWChisel.scala 171:39]
  wire [15:0] array_9_io_e_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_9_io_f_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_9_io_ve_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_9_io_vf_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_9_io_vv_i; // @[SWChisel.scala 171:39]
  wire [15:0] array_9_io_e_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_9_io_f_o; // @[SWChisel.scala 171:39]
  wire [15:0] array_9_io_v_o; // @[SWChisel.scala 171:39]
  wire  r_count_0_clock; // @[SWChisel.scala 172:41]
  wire  r_count_0_reset; // @[SWChisel.scala 172:41]
  wire  r_count_0_io_en; // @[SWChisel.scala 172:41]
  wire [4:0] r_count_0_io_out; // @[SWChisel.scala 172:41]
  wire  r_count_1_clock; // @[SWChisel.scala 172:41]
  wire  r_count_1_reset; // @[SWChisel.scala 172:41]
  wire  r_count_1_io_en; // @[SWChisel.scala 172:41]
  wire [4:0] r_count_1_io_out; // @[SWChisel.scala 172:41]
  wire  r_count_2_clock; // @[SWChisel.scala 172:41]
  wire  r_count_2_reset; // @[SWChisel.scala 172:41]
  wire  r_count_2_io_en; // @[SWChisel.scala 172:41]
  wire [4:0] r_count_2_io_out; // @[SWChisel.scala 172:41]
  wire  r_count_3_clock; // @[SWChisel.scala 172:41]
  wire  r_count_3_reset; // @[SWChisel.scala 172:41]
  wire  r_count_3_io_en; // @[SWChisel.scala 172:41]
  wire [4:0] r_count_3_io_out; // @[SWChisel.scala 172:41]
  wire  r_count_4_clock; // @[SWChisel.scala 172:41]
  wire  r_count_4_reset; // @[SWChisel.scala 172:41]
  wire  r_count_4_io_en; // @[SWChisel.scala 172:41]
  wire [4:0] r_count_4_io_out; // @[SWChisel.scala 172:41]
  wire  r_count_5_clock; // @[SWChisel.scala 172:41]
  wire  r_count_5_reset; // @[SWChisel.scala 172:41]
  wire  r_count_5_io_en; // @[SWChisel.scala 172:41]
  wire [4:0] r_count_5_io_out; // @[SWChisel.scala 172:41]
  wire  r_count_6_clock; // @[SWChisel.scala 172:41]
  wire  r_count_6_reset; // @[SWChisel.scala 172:41]
  wire  r_count_6_io_en; // @[SWChisel.scala 172:41]
  wire [4:0] r_count_6_io_out; // @[SWChisel.scala 172:41]
  wire  r_count_7_clock; // @[SWChisel.scala 172:41]
  wire  r_count_7_reset; // @[SWChisel.scala 172:41]
  wire  r_count_7_io_en; // @[SWChisel.scala 172:41]
  wire [4:0] r_count_7_io_out; // @[SWChisel.scala 172:41]
  wire  r_count_8_clock; // @[SWChisel.scala 172:41]
  wire  r_count_8_reset; // @[SWChisel.scala 172:41]
  wire  r_count_8_io_en; // @[SWChisel.scala 172:41]
  wire [4:0] r_count_8_io_out; // @[SWChisel.scala 172:41]
  wire  r_count_9_clock; // @[SWChisel.scala 172:41]
  wire  r_count_9_reset; // @[SWChisel.scala 172:41]
  wire  r_count_9_io_en; // @[SWChisel.scala 172:41]
  wire [4:0] r_count_9_io_out; // @[SWChisel.scala 172:41]
  wire  max_clock; // @[SWChisel.scala 175:19]
  wire  max_reset; // @[SWChisel.scala 175:19]
  wire  max_io_start; // @[SWChisel.scala 175:19]
  wire [15:0] max_io_in; // @[SWChisel.scala 175:19]
  wire  max_io_done; // @[SWChisel.scala 175:19]
  wire [15:0] max_io_out; // @[SWChisel.scala 175:19]
  reg [15:0] E_0; // @[SWChisel.scala 162:18]
  reg [15:0] E_1; // @[SWChisel.scala 162:18]
  reg [15:0] E_2; // @[SWChisel.scala 162:18]
  reg [15:0] E_3; // @[SWChisel.scala 162:18]
  reg [15:0] E_4; // @[SWChisel.scala 162:18]
  reg [15:0] E_5; // @[SWChisel.scala 162:18]
  reg [15:0] E_6; // @[SWChisel.scala 162:18]
  reg [15:0] E_7; // @[SWChisel.scala 162:18]
  reg [15:0] E_8; // @[SWChisel.scala 162:18]
  reg [15:0] E_9; // @[SWChisel.scala 162:18]
  reg [15:0] F_1; // @[SWChisel.scala 163:18]
  reg [15:0] F_2; // @[SWChisel.scala 163:18]
  reg [15:0] F_3; // @[SWChisel.scala 163:18]
  reg [15:0] F_4; // @[SWChisel.scala 163:18]
  reg [15:0] F_5; // @[SWChisel.scala 163:18]
  reg [15:0] F_6; // @[SWChisel.scala 163:18]
  reg [15:0] F_7; // @[SWChisel.scala 163:18]
  reg [15:0] F_8; // @[SWChisel.scala 163:18]
  reg [15:0] F_9; // @[SWChisel.scala 163:18]
  reg [15:0] F_10; // @[SWChisel.scala 163:18]
  reg [15:0] V1_1; // @[SWChisel.scala 164:19]
  reg [15:0] V1_2; // @[SWChisel.scala 164:19]
  reg [15:0] V1_3; // @[SWChisel.scala 164:19]
  reg [15:0] V1_4; // @[SWChisel.scala 164:19]
  reg [15:0] V1_5; // @[SWChisel.scala 164:19]
  reg [15:0] V1_6; // @[SWChisel.scala 164:19]
  reg [15:0] V1_7; // @[SWChisel.scala 164:19]
  reg [15:0] V1_8; // @[SWChisel.scala 164:19]
  reg [15:0] V1_9; // @[SWChisel.scala 164:19]
  reg [15:0] V1_10; // @[SWChisel.scala 164:19]
  reg [15:0] V2_1; // @[SWChisel.scala 167:19]
  reg [15:0] V2_2; // @[SWChisel.scala 167:19]
  reg [15:0] V2_3; // @[SWChisel.scala 167:19]
  reg [15:0] V2_4; // @[SWChisel.scala 167:19]
  reg [15:0] V2_5; // @[SWChisel.scala 167:19]
  reg [15:0] V2_6; // @[SWChisel.scala 167:19]
  reg [15:0] V2_7; // @[SWChisel.scala 167:19]
  reg [15:0] V2_8; // @[SWChisel.scala 167:19]
  reg [15:0] V2_9; // @[SWChisel.scala 167:19]
  reg [15:0] V2_10; // @[SWChisel.scala 167:19]
  reg  start_reg_0; // @[SWChisel.scala 168:26]
  reg  start_reg_1; // @[SWChisel.scala 168:26]
  reg  start_reg_2; // @[SWChisel.scala 168:26]
  reg  start_reg_3; // @[SWChisel.scala 168:26]
  reg  start_reg_4; // @[SWChisel.scala 168:26]
  reg  start_reg_5; // @[SWChisel.scala 168:26]
  reg  start_reg_6; // @[SWChisel.scala 168:26]
  reg  start_reg_7; // @[SWChisel.scala 168:26]
  reg  start_reg_8; // @[SWChisel.scala 168:26]
  reg  start_reg_9; // @[SWChisel.scala 168:26]
  wire [1:0] _GEN_31 = 5'h1 == r_count_0_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_32 = 5'h2 == r_count_0_io_out ? io_r_2_b : _GEN_31; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_33 = 5'h3 == r_count_0_io_out ? io_r_3_b : _GEN_32; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_34 = 5'h4 == r_count_0_io_out ? io_r_4_b : _GEN_33; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_35 = 5'h5 == r_count_0_io_out ? io_r_5_b : _GEN_34; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_36 = 5'h6 == r_count_0_io_out ? io_r_6_b : _GEN_35; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_37 = 5'h7 == r_count_0_io_out ? io_r_7_b : _GEN_36; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_38 = 5'h8 == r_count_0_io_out ? io_r_8_b : _GEN_37; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_39 = 5'h9 == r_count_0_io_out ? io_r_9_b : _GEN_38; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_40 = 5'ha == r_count_0_io_out ? io_r_10_b : _GEN_39; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_41 = 5'hb == r_count_0_io_out ? io_r_11_b : _GEN_40; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_42 = 5'hc == r_count_0_io_out ? io_r_12_b : _GEN_41; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_43 = 5'hd == r_count_0_io_out ? io_r_13_b : _GEN_42; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_44 = 5'he == r_count_0_io_out ? io_r_14_b : _GEN_43; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_45 = 5'hf == r_count_0_io_out ? io_r_15_b : _GEN_44; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_48 = 5'h1 == r_count_1_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_49 = 5'h2 == r_count_1_io_out ? io_r_2_b : _GEN_48; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_50 = 5'h3 == r_count_1_io_out ? io_r_3_b : _GEN_49; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_51 = 5'h4 == r_count_1_io_out ? io_r_4_b : _GEN_50; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_52 = 5'h5 == r_count_1_io_out ? io_r_5_b : _GEN_51; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_53 = 5'h6 == r_count_1_io_out ? io_r_6_b : _GEN_52; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_54 = 5'h7 == r_count_1_io_out ? io_r_7_b : _GEN_53; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_55 = 5'h8 == r_count_1_io_out ? io_r_8_b : _GEN_54; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_56 = 5'h9 == r_count_1_io_out ? io_r_9_b : _GEN_55; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_57 = 5'ha == r_count_1_io_out ? io_r_10_b : _GEN_56; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_58 = 5'hb == r_count_1_io_out ? io_r_11_b : _GEN_57; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_59 = 5'hc == r_count_1_io_out ? io_r_12_b : _GEN_58; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_60 = 5'hd == r_count_1_io_out ? io_r_13_b : _GEN_59; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_61 = 5'he == r_count_1_io_out ? io_r_14_b : _GEN_60; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_62 = 5'hf == r_count_1_io_out ? io_r_15_b : _GEN_61; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_65 = 5'h1 == r_count_2_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_66 = 5'h2 == r_count_2_io_out ? io_r_2_b : _GEN_65; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_67 = 5'h3 == r_count_2_io_out ? io_r_3_b : _GEN_66; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_68 = 5'h4 == r_count_2_io_out ? io_r_4_b : _GEN_67; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_69 = 5'h5 == r_count_2_io_out ? io_r_5_b : _GEN_68; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_70 = 5'h6 == r_count_2_io_out ? io_r_6_b : _GEN_69; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_71 = 5'h7 == r_count_2_io_out ? io_r_7_b : _GEN_70; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_72 = 5'h8 == r_count_2_io_out ? io_r_8_b : _GEN_71; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_73 = 5'h9 == r_count_2_io_out ? io_r_9_b : _GEN_72; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_74 = 5'ha == r_count_2_io_out ? io_r_10_b : _GEN_73; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_75 = 5'hb == r_count_2_io_out ? io_r_11_b : _GEN_74; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_76 = 5'hc == r_count_2_io_out ? io_r_12_b : _GEN_75; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_77 = 5'hd == r_count_2_io_out ? io_r_13_b : _GEN_76; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_78 = 5'he == r_count_2_io_out ? io_r_14_b : _GEN_77; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_79 = 5'hf == r_count_2_io_out ? io_r_15_b : _GEN_78; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_82 = 5'h1 == r_count_3_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_83 = 5'h2 == r_count_3_io_out ? io_r_2_b : _GEN_82; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_84 = 5'h3 == r_count_3_io_out ? io_r_3_b : _GEN_83; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_85 = 5'h4 == r_count_3_io_out ? io_r_4_b : _GEN_84; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_86 = 5'h5 == r_count_3_io_out ? io_r_5_b : _GEN_85; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_87 = 5'h6 == r_count_3_io_out ? io_r_6_b : _GEN_86; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_88 = 5'h7 == r_count_3_io_out ? io_r_7_b : _GEN_87; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_89 = 5'h8 == r_count_3_io_out ? io_r_8_b : _GEN_88; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_90 = 5'h9 == r_count_3_io_out ? io_r_9_b : _GEN_89; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_91 = 5'ha == r_count_3_io_out ? io_r_10_b : _GEN_90; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_92 = 5'hb == r_count_3_io_out ? io_r_11_b : _GEN_91; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_93 = 5'hc == r_count_3_io_out ? io_r_12_b : _GEN_92; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_94 = 5'hd == r_count_3_io_out ? io_r_13_b : _GEN_93; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_95 = 5'he == r_count_3_io_out ? io_r_14_b : _GEN_94; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_96 = 5'hf == r_count_3_io_out ? io_r_15_b : _GEN_95; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_99 = 5'h1 == r_count_4_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_100 = 5'h2 == r_count_4_io_out ? io_r_2_b : _GEN_99; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_101 = 5'h3 == r_count_4_io_out ? io_r_3_b : _GEN_100; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_102 = 5'h4 == r_count_4_io_out ? io_r_4_b : _GEN_101; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_103 = 5'h5 == r_count_4_io_out ? io_r_5_b : _GEN_102; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_104 = 5'h6 == r_count_4_io_out ? io_r_6_b : _GEN_103; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_105 = 5'h7 == r_count_4_io_out ? io_r_7_b : _GEN_104; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_106 = 5'h8 == r_count_4_io_out ? io_r_8_b : _GEN_105; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_107 = 5'h9 == r_count_4_io_out ? io_r_9_b : _GEN_106; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_108 = 5'ha == r_count_4_io_out ? io_r_10_b : _GEN_107; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_109 = 5'hb == r_count_4_io_out ? io_r_11_b : _GEN_108; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_110 = 5'hc == r_count_4_io_out ? io_r_12_b : _GEN_109; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_111 = 5'hd == r_count_4_io_out ? io_r_13_b : _GEN_110; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_112 = 5'he == r_count_4_io_out ? io_r_14_b : _GEN_111; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_113 = 5'hf == r_count_4_io_out ? io_r_15_b : _GEN_112; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_116 = 5'h1 == r_count_5_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_117 = 5'h2 == r_count_5_io_out ? io_r_2_b : _GEN_116; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_118 = 5'h3 == r_count_5_io_out ? io_r_3_b : _GEN_117; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_119 = 5'h4 == r_count_5_io_out ? io_r_4_b : _GEN_118; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_120 = 5'h5 == r_count_5_io_out ? io_r_5_b : _GEN_119; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_121 = 5'h6 == r_count_5_io_out ? io_r_6_b : _GEN_120; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_122 = 5'h7 == r_count_5_io_out ? io_r_7_b : _GEN_121; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_123 = 5'h8 == r_count_5_io_out ? io_r_8_b : _GEN_122; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_124 = 5'h9 == r_count_5_io_out ? io_r_9_b : _GEN_123; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_125 = 5'ha == r_count_5_io_out ? io_r_10_b : _GEN_124; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_126 = 5'hb == r_count_5_io_out ? io_r_11_b : _GEN_125; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_127 = 5'hc == r_count_5_io_out ? io_r_12_b : _GEN_126; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_128 = 5'hd == r_count_5_io_out ? io_r_13_b : _GEN_127; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_129 = 5'he == r_count_5_io_out ? io_r_14_b : _GEN_128; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_130 = 5'hf == r_count_5_io_out ? io_r_15_b : _GEN_129; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_133 = 5'h1 == r_count_6_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_134 = 5'h2 == r_count_6_io_out ? io_r_2_b : _GEN_133; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_135 = 5'h3 == r_count_6_io_out ? io_r_3_b : _GEN_134; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_136 = 5'h4 == r_count_6_io_out ? io_r_4_b : _GEN_135; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_137 = 5'h5 == r_count_6_io_out ? io_r_5_b : _GEN_136; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_138 = 5'h6 == r_count_6_io_out ? io_r_6_b : _GEN_137; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_139 = 5'h7 == r_count_6_io_out ? io_r_7_b : _GEN_138; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_140 = 5'h8 == r_count_6_io_out ? io_r_8_b : _GEN_139; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_141 = 5'h9 == r_count_6_io_out ? io_r_9_b : _GEN_140; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_142 = 5'ha == r_count_6_io_out ? io_r_10_b : _GEN_141; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_143 = 5'hb == r_count_6_io_out ? io_r_11_b : _GEN_142; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_144 = 5'hc == r_count_6_io_out ? io_r_12_b : _GEN_143; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_145 = 5'hd == r_count_6_io_out ? io_r_13_b : _GEN_144; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_146 = 5'he == r_count_6_io_out ? io_r_14_b : _GEN_145; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_147 = 5'hf == r_count_6_io_out ? io_r_15_b : _GEN_146; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_150 = 5'h1 == r_count_7_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_151 = 5'h2 == r_count_7_io_out ? io_r_2_b : _GEN_150; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_152 = 5'h3 == r_count_7_io_out ? io_r_3_b : _GEN_151; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_153 = 5'h4 == r_count_7_io_out ? io_r_4_b : _GEN_152; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_154 = 5'h5 == r_count_7_io_out ? io_r_5_b : _GEN_153; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_155 = 5'h6 == r_count_7_io_out ? io_r_6_b : _GEN_154; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_156 = 5'h7 == r_count_7_io_out ? io_r_7_b : _GEN_155; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_157 = 5'h8 == r_count_7_io_out ? io_r_8_b : _GEN_156; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_158 = 5'h9 == r_count_7_io_out ? io_r_9_b : _GEN_157; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_159 = 5'ha == r_count_7_io_out ? io_r_10_b : _GEN_158; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_160 = 5'hb == r_count_7_io_out ? io_r_11_b : _GEN_159; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_161 = 5'hc == r_count_7_io_out ? io_r_12_b : _GEN_160; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_162 = 5'hd == r_count_7_io_out ? io_r_13_b : _GEN_161; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_163 = 5'he == r_count_7_io_out ? io_r_14_b : _GEN_162; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_164 = 5'hf == r_count_7_io_out ? io_r_15_b : _GEN_163; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_167 = 5'h1 == r_count_8_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_168 = 5'h2 == r_count_8_io_out ? io_r_2_b : _GEN_167; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_169 = 5'h3 == r_count_8_io_out ? io_r_3_b : _GEN_168; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_170 = 5'h4 == r_count_8_io_out ? io_r_4_b : _GEN_169; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_171 = 5'h5 == r_count_8_io_out ? io_r_5_b : _GEN_170; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_172 = 5'h6 == r_count_8_io_out ? io_r_6_b : _GEN_171; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_173 = 5'h7 == r_count_8_io_out ? io_r_7_b : _GEN_172; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_174 = 5'h8 == r_count_8_io_out ? io_r_8_b : _GEN_173; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_175 = 5'h9 == r_count_8_io_out ? io_r_9_b : _GEN_174; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_176 = 5'ha == r_count_8_io_out ? io_r_10_b : _GEN_175; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_177 = 5'hb == r_count_8_io_out ? io_r_11_b : _GEN_176; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_178 = 5'hc == r_count_8_io_out ? io_r_12_b : _GEN_177; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_179 = 5'hd == r_count_8_io_out ? io_r_13_b : _GEN_178; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_180 = 5'he == r_count_8_io_out ? io_r_14_b : _GEN_179; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_181 = 5'hf == r_count_8_io_out ? io_r_15_b : _GEN_180; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_184 = 5'h1 == r_count_9_io_out ? io_r_1_b : io_r_0_b; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_185 = 5'h2 == r_count_9_io_out ? io_r_2_b : _GEN_184; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_186 = 5'h3 == r_count_9_io_out ? io_r_3_b : _GEN_185; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_187 = 5'h4 == r_count_9_io_out ? io_r_4_b : _GEN_186; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_188 = 5'h5 == r_count_9_io_out ? io_r_5_b : _GEN_187; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_189 = 5'h6 == r_count_9_io_out ? io_r_6_b : _GEN_188; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_190 = 5'h7 == r_count_9_io_out ? io_r_7_b : _GEN_189; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_191 = 5'h8 == r_count_9_io_out ? io_r_8_b : _GEN_190; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_192 = 5'h9 == r_count_9_io_out ? io_r_9_b : _GEN_191; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_193 = 5'ha == r_count_9_io_out ? io_r_10_b : _GEN_192; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_194 = 5'hb == r_count_9_io_out ? io_r_11_b : _GEN_193; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_195 = 5'hc == r_count_9_io_out ? io_r_12_b : _GEN_194; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_196 = 5'hd == r_count_9_io_out ? io_r_13_b : _GEN_195; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_197 = 5'he == r_count_9_io_out ? io_r_14_b : _GEN_196; // @[SWChisel.scala 222:{19,19}]
  wire [1:0] _GEN_198 = 5'hf == r_count_9_io_out ? io_r_15_b : _GEN_197; // @[SWChisel.scala 222:{19,19}]
  SWCell array_0 ( // @[SWChisel.scala 171:39]
    .io_q(array_0_io_q),
    .io_r(array_0_io_r),
    .io_e_i(array_0_io_e_i),
    .io_f_i(array_0_io_f_i),
    .io_ve_i(array_0_io_ve_i),
    .io_vf_i(array_0_io_vf_i),
    .io_vv_i(array_0_io_vv_i),
    .io_e_o(array_0_io_e_o),
    .io_f_o(array_0_io_f_o),
    .io_v_o(array_0_io_v_o)
  );
  SWCell array_1 ( // @[SWChisel.scala 171:39]
    .io_q(array_1_io_q),
    .io_r(array_1_io_r),
    .io_e_i(array_1_io_e_i),
    .io_f_i(array_1_io_f_i),
    .io_ve_i(array_1_io_ve_i),
    .io_vf_i(array_1_io_vf_i),
    .io_vv_i(array_1_io_vv_i),
    .io_e_o(array_1_io_e_o),
    .io_f_o(array_1_io_f_o),
    .io_v_o(array_1_io_v_o)
  );
  SWCell array_2 ( // @[SWChisel.scala 171:39]
    .io_q(array_2_io_q),
    .io_r(array_2_io_r),
    .io_e_i(array_2_io_e_i),
    .io_f_i(array_2_io_f_i),
    .io_ve_i(array_2_io_ve_i),
    .io_vf_i(array_2_io_vf_i),
    .io_vv_i(array_2_io_vv_i),
    .io_e_o(array_2_io_e_o),
    .io_f_o(array_2_io_f_o),
    .io_v_o(array_2_io_v_o)
  );
  SWCell array_3 ( // @[SWChisel.scala 171:39]
    .io_q(array_3_io_q),
    .io_r(array_3_io_r),
    .io_e_i(array_3_io_e_i),
    .io_f_i(array_3_io_f_i),
    .io_ve_i(array_3_io_ve_i),
    .io_vf_i(array_3_io_vf_i),
    .io_vv_i(array_3_io_vv_i),
    .io_e_o(array_3_io_e_o),
    .io_f_o(array_3_io_f_o),
    .io_v_o(array_3_io_v_o)
  );
  SWCell array_4 ( // @[SWChisel.scala 171:39]
    .io_q(array_4_io_q),
    .io_r(array_4_io_r),
    .io_e_i(array_4_io_e_i),
    .io_f_i(array_4_io_f_i),
    .io_ve_i(array_4_io_ve_i),
    .io_vf_i(array_4_io_vf_i),
    .io_vv_i(array_4_io_vv_i),
    .io_e_o(array_4_io_e_o),
    .io_f_o(array_4_io_f_o),
    .io_v_o(array_4_io_v_o)
  );
  SWCell array_5 ( // @[SWChisel.scala 171:39]
    .io_q(array_5_io_q),
    .io_r(array_5_io_r),
    .io_e_i(array_5_io_e_i),
    .io_f_i(array_5_io_f_i),
    .io_ve_i(array_5_io_ve_i),
    .io_vf_i(array_5_io_vf_i),
    .io_vv_i(array_5_io_vv_i),
    .io_e_o(array_5_io_e_o),
    .io_f_o(array_5_io_f_o),
    .io_v_o(array_5_io_v_o)
  );
  SWCell array_6 ( // @[SWChisel.scala 171:39]
    .io_q(array_6_io_q),
    .io_r(array_6_io_r),
    .io_e_i(array_6_io_e_i),
    .io_f_i(array_6_io_f_i),
    .io_ve_i(array_6_io_ve_i),
    .io_vf_i(array_6_io_vf_i),
    .io_vv_i(array_6_io_vv_i),
    .io_e_o(array_6_io_e_o),
    .io_f_o(array_6_io_f_o),
    .io_v_o(array_6_io_v_o)
  );
  SWCell array_7 ( // @[SWChisel.scala 171:39]
    .io_q(array_7_io_q),
    .io_r(array_7_io_r),
    .io_e_i(array_7_io_e_i),
    .io_f_i(array_7_io_f_i),
    .io_ve_i(array_7_io_ve_i),
    .io_vf_i(array_7_io_vf_i),
    .io_vv_i(array_7_io_vv_i),
    .io_e_o(array_7_io_e_o),
    .io_f_o(array_7_io_f_o),
    .io_v_o(array_7_io_v_o)
  );
  SWCell array_8 ( // @[SWChisel.scala 171:39]
    .io_q(array_8_io_q),
    .io_r(array_8_io_r),
    .io_e_i(array_8_io_e_i),
    .io_f_i(array_8_io_f_i),
    .io_ve_i(array_8_io_ve_i),
    .io_vf_i(array_8_io_vf_i),
    .io_vv_i(array_8_io_vv_i),
    .io_e_o(array_8_io_e_o),
    .io_f_o(array_8_io_f_o),
    .io_v_o(array_8_io_v_o)
  );
  SWCell array_9 ( // @[SWChisel.scala 171:39]
    .io_q(array_9_io_q),
    .io_r(array_9_io_r),
    .io_e_i(array_9_io_e_i),
    .io_f_i(array_9_io_f_i),
    .io_ve_i(array_9_io_ve_i),
    .io_vf_i(array_9_io_vf_i),
    .io_vv_i(array_9_io_vv_i),
    .io_e_o(array_9_io_e_o),
    .io_f_o(array_9_io_f_o),
    .io_v_o(array_9_io_v_o)
  );
  MyCounter r_count_0 ( // @[SWChisel.scala 172:41]
    .clock(r_count_0_clock),
    .reset(r_count_0_reset),
    .io_en(r_count_0_io_en),
    .io_out(r_count_0_io_out)
  );
  MyCounter r_count_1 ( // @[SWChisel.scala 172:41]
    .clock(r_count_1_clock),
    .reset(r_count_1_reset),
    .io_en(r_count_1_io_en),
    .io_out(r_count_1_io_out)
  );
  MyCounter r_count_2 ( // @[SWChisel.scala 172:41]
    .clock(r_count_2_clock),
    .reset(r_count_2_reset),
    .io_en(r_count_2_io_en),
    .io_out(r_count_2_io_out)
  );
  MyCounter r_count_3 ( // @[SWChisel.scala 172:41]
    .clock(r_count_3_clock),
    .reset(r_count_3_reset),
    .io_en(r_count_3_io_en),
    .io_out(r_count_3_io_out)
  );
  MyCounter r_count_4 ( // @[SWChisel.scala 172:41]
    .clock(r_count_4_clock),
    .reset(r_count_4_reset),
    .io_en(r_count_4_io_en),
    .io_out(r_count_4_io_out)
  );
  MyCounter r_count_5 ( // @[SWChisel.scala 172:41]
    .clock(r_count_5_clock),
    .reset(r_count_5_reset),
    .io_en(r_count_5_io_en),
    .io_out(r_count_5_io_out)
  );
  MyCounter r_count_6 ( // @[SWChisel.scala 172:41]
    .clock(r_count_6_clock),
    .reset(r_count_6_reset),
    .io_en(r_count_6_io_en),
    .io_out(r_count_6_io_out)
  );
  MyCounter r_count_7 ( // @[SWChisel.scala 172:41]
    .clock(r_count_7_clock),
    .reset(r_count_7_reset),
    .io_en(r_count_7_io_en),
    .io_out(r_count_7_io_out)
  );
  MyCounter r_count_8 ( // @[SWChisel.scala 172:41]
    .clock(r_count_8_clock),
    .reset(r_count_8_reset),
    .io_en(r_count_8_io_en),
    .io_out(r_count_8_io_out)
  );
  MyCounter r_count_9 ( // @[SWChisel.scala 172:41]
    .clock(r_count_9_clock),
    .reset(r_count_9_reset),
    .io_en(r_count_9_io_en),
    .io_out(r_count_9_io_out)
  );
  MAX max ( // @[SWChisel.scala 175:19]
    .clock(max_clock),
    .reset(max_reset),
    .io_start(max_io_start),
    .io_in(max_io_in),
    .io_done(max_io_done),
    .io_out(max_io_out)
  );
  assign io_result = max_io_out; // @[SWChisel.scala 182:13]
  assign io_done = max_io_done; // @[SWChisel.scala 183:11]
  assign io_v1_out_0 = 16'sh0; // @[SWChisel.scala 242:24]
  assign io_v1_out_1 = V1_1; // @[SWChisel.scala 242:24]
  assign io_v1_out_2 = V1_2; // @[SWChisel.scala 242:24]
  assign io_v1_out_3 = V1_3; // @[SWChisel.scala 242:24]
  assign io_v1_out_4 = V1_4; // @[SWChisel.scala 242:24]
  assign io_v1_out_5 = V1_5; // @[SWChisel.scala 242:24]
  assign io_v1_out_6 = V1_6; // @[SWChisel.scala 242:24]
  assign io_v1_out_7 = V1_7; // @[SWChisel.scala 242:24]
  assign io_v1_out_8 = V1_8; // @[SWChisel.scala 242:24]
  assign io_v1_out_9 = V1_9; // @[SWChisel.scala 242:24]
  assign io_v1_out_10 = V1_10; // @[SWChisel.scala 242:24]
  assign io_v2_out_0 = 16'sh0; // @[SWChisel.scala 245:24]
  assign io_v2_out_1 = V2_1; // @[SWChisel.scala 245:24]
  assign io_v2_out_2 = V2_2; // @[SWChisel.scala 245:24]
  assign io_v2_out_3 = V2_3; // @[SWChisel.scala 245:24]
  assign io_v2_out_4 = V2_4; // @[SWChisel.scala 245:24]
  assign io_v2_out_5 = V2_5; // @[SWChisel.scala 245:24]
  assign io_v2_out_6 = V2_6; // @[SWChisel.scala 245:24]
  assign io_v2_out_7 = V2_7; // @[SWChisel.scala 245:24]
  assign io_v2_out_8 = V2_8; // @[SWChisel.scala 245:24]
  assign io_v2_out_9 = V2_9; // @[SWChisel.scala 245:24]
  assign io_v2_out_10 = V2_10; // @[SWChisel.scala 245:24]
  assign io_e_out_0 = E_0; // @[SWChisel.scala 233:23]
  assign io_e_out_1 = E_1; // @[SWChisel.scala 233:23]
  assign io_e_out_2 = E_2; // @[SWChisel.scala 233:23]
  assign io_e_out_3 = E_3; // @[SWChisel.scala 233:23]
  assign io_e_out_4 = E_4; // @[SWChisel.scala 233:23]
  assign io_e_out_5 = E_5; // @[SWChisel.scala 233:23]
  assign io_e_out_6 = E_6; // @[SWChisel.scala 233:23]
  assign io_e_out_7 = E_7; // @[SWChisel.scala 233:23]
  assign io_e_out_8 = E_8; // @[SWChisel.scala 233:23]
  assign io_e_out_9 = E_9; // @[SWChisel.scala 233:23]
  assign io_f_out_0 = 16'sh0; // @[SWChisel.scala 239:23]
  assign io_f_out_1 = F_1; // @[SWChisel.scala 239:23]
  assign io_f_out_2 = F_2; // @[SWChisel.scala 239:23]
  assign io_f_out_3 = F_3; // @[SWChisel.scala 239:23]
  assign io_f_out_4 = F_4; // @[SWChisel.scala 239:23]
  assign io_f_out_5 = F_5; // @[SWChisel.scala 239:23]
  assign io_f_out_6 = F_6; // @[SWChisel.scala 239:23]
  assign io_f_out_7 = F_7; // @[SWChisel.scala 239:23]
  assign io_f_out_8 = F_8; // @[SWChisel.scala 239:23]
  assign io_f_out_9 = F_9; // @[SWChisel.scala 239:23]
  assign io_f_out_10 = F_10; // @[SWChisel.scala 239:23]
  assign array_0_io_q = io_q_0_b; // @[SWChisel.scala 221:19]
  assign array_0_io_r = 5'h10 == r_count_0_io_out ? io_r_16_b : _GEN_45; // @[SWChisel.scala 222:{19,19}]
  assign array_0_io_e_i = E_0; // @[SWChisel.scala 197:21]
  assign array_0_io_f_i = 16'sh0; // @[SWChisel.scala 199:21]
  assign array_0_io_ve_i = V1_1; // @[SWChisel.scala 198:22]
  assign array_0_io_vf_i = 16'sh0; // @[SWChisel.scala 200:22]
  assign array_0_io_vv_i = 16'sh0; // @[SWChisel.scala 201:22]
  assign array_1_io_q = io_q_1_b; // @[SWChisel.scala 221:19]
  assign array_1_io_r = 5'h10 == r_count_1_io_out ? io_r_16_b : _GEN_62; // @[SWChisel.scala 222:{19,19}]
  assign array_1_io_e_i = E_1; // @[SWChisel.scala 197:21]
  assign array_1_io_f_i = F_1; // @[SWChisel.scala 199:21]
  assign array_1_io_ve_i = V1_2; // @[SWChisel.scala 198:22]
  assign array_1_io_vf_i = V1_1; // @[SWChisel.scala 200:22]
  assign array_1_io_vv_i = V2_1; // @[SWChisel.scala 201:22]
  assign array_2_io_q = io_q_2_b; // @[SWChisel.scala 221:19]
  assign array_2_io_r = 5'h10 == r_count_2_io_out ? io_r_16_b : _GEN_79; // @[SWChisel.scala 222:{19,19}]
  assign array_2_io_e_i = E_2; // @[SWChisel.scala 197:21]
  assign array_2_io_f_i = F_2; // @[SWChisel.scala 199:21]
  assign array_2_io_ve_i = V1_3; // @[SWChisel.scala 198:22]
  assign array_2_io_vf_i = V1_2; // @[SWChisel.scala 200:22]
  assign array_2_io_vv_i = V2_2; // @[SWChisel.scala 201:22]
  assign array_3_io_q = io_q_3_b; // @[SWChisel.scala 221:19]
  assign array_3_io_r = 5'h10 == r_count_3_io_out ? io_r_16_b : _GEN_96; // @[SWChisel.scala 222:{19,19}]
  assign array_3_io_e_i = E_3; // @[SWChisel.scala 197:21]
  assign array_3_io_f_i = F_3; // @[SWChisel.scala 199:21]
  assign array_3_io_ve_i = V1_4; // @[SWChisel.scala 198:22]
  assign array_3_io_vf_i = V1_3; // @[SWChisel.scala 200:22]
  assign array_3_io_vv_i = V2_3; // @[SWChisel.scala 201:22]
  assign array_4_io_q = io_q_4_b; // @[SWChisel.scala 221:19]
  assign array_4_io_r = 5'h10 == r_count_4_io_out ? io_r_16_b : _GEN_113; // @[SWChisel.scala 222:{19,19}]
  assign array_4_io_e_i = E_4; // @[SWChisel.scala 197:21]
  assign array_4_io_f_i = F_4; // @[SWChisel.scala 199:21]
  assign array_4_io_ve_i = V1_5; // @[SWChisel.scala 198:22]
  assign array_4_io_vf_i = V1_4; // @[SWChisel.scala 200:22]
  assign array_4_io_vv_i = V2_4; // @[SWChisel.scala 201:22]
  assign array_5_io_q = io_q_5_b; // @[SWChisel.scala 221:19]
  assign array_5_io_r = 5'h10 == r_count_5_io_out ? io_r_16_b : _GEN_130; // @[SWChisel.scala 222:{19,19}]
  assign array_5_io_e_i = E_5; // @[SWChisel.scala 197:21]
  assign array_5_io_f_i = F_5; // @[SWChisel.scala 199:21]
  assign array_5_io_ve_i = V1_6; // @[SWChisel.scala 198:22]
  assign array_5_io_vf_i = V1_5; // @[SWChisel.scala 200:22]
  assign array_5_io_vv_i = V2_5; // @[SWChisel.scala 201:22]
  assign array_6_io_q = io_q_6_b; // @[SWChisel.scala 221:19]
  assign array_6_io_r = 5'h10 == r_count_6_io_out ? io_r_16_b : _GEN_147; // @[SWChisel.scala 222:{19,19}]
  assign array_6_io_e_i = E_6; // @[SWChisel.scala 197:21]
  assign array_6_io_f_i = F_6; // @[SWChisel.scala 199:21]
  assign array_6_io_ve_i = V1_7; // @[SWChisel.scala 198:22]
  assign array_6_io_vf_i = V1_6; // @[SWChisel.scala 200:22]
  assign array_6_io_vv_i = V2_6; // @[SWChisel.scala 201:22]
  assign array_7_io_q = io_q_7_b; // @[SWChisel.scala 221:19]
  assign array_7_io_r = 5'h10 == r_count_7_io_out ? io_r_16_b : _GEN_164; // @[SWChisel.scala 222:{19,19}]
  assign array_7_io_e_i = E_7; // @[SWChisel.scala 197:21]
  assign array_7_io_f_i = F_7; // @[SWChisel.scala 199:21]
  assign array_7_io_ve_i = V1_8; // @[SWChisel.scala 198:22]
  assign array_7_io_vf_i = V1_7; // @[SWChisel.scala 200:22]
  assign array_7_io_vv_i = V2_7; // @[SWChisel.scala 201:22]
  assign array_8_io_q = io_q_8_b; // @[SWChisel.scala 221:19]
  assign array_8_io_r = 5'h10 == r_count_8_io_out ? io_r_16_b : _GEN_181; // @[SWChisel.scala 222:{19,19}]
  assign array_8_io_e_i = E_8; // @[SWChisel.scala 197:21]
  assign array_8_io_f_i = F_8; // @[SWChisel.scala 199:21]
  assign array_8_io_ve_i = V1_9; // @[SWChisel.scala 198:22]
  assign array_8_io_vf_i = V1_8; // @[SWChisel.scala 200:22]
  assign array_8_io_vv_i = V2_8; // @[SWChisel.scala 201:22]
  assign array_9_io_q = io_q_9_b; // @[SWChisel.scala 221:19]
  assign array_9_io_r = 5'h10 == r_count_9_io_out ? io_r_16_b : _GEN_198; // @[SWChisel.scala 222:{19,19}]
  assign array_9_io_e_i = E_9; // @[SWChisel.scala 197:21]
  assign array_9_io_f_i = F_9; // @[SWChisel.scala 199:21]
  assign array_9_io_ve_i = V1_10; // @[SWChisel.scala 198:22]
  assign array_9_io_vf_i = V1_9; // @[SWChisel.scala 200:22]
  assign array_9_io_vv_i = V2_9; // @[SWChisel.scala 201:22]
  assign r_count_0_clock = clock;
  assign r_count_0_reset = reset;
  assign r_count_0_io_en = start_reg_0; // @[SWChisel.scala 193:22]
  assign r_count_1_clock = clock;
  assign r_count_1_reset = reset;
  assign r_count_1_io_en = start_reg_1; // @[SWChisel.scala 193:22]
  assign r_count_2_clock = clock;
  assign r_count_2_reset = reset;
  assign r_count_2_io_en = start_reg_2; // @[SWChisel.scala 193:22]
  assign r_count_3_clock = clock;
  assign r_count_3_reset = reset;
  assign r_count_3_io_en = start_reg_3; // @[SWChisel.scala 193:22]
  assign r_count_4_clock = clock;
  assign r_count_4_reset = reset;
  assign r_count_4_io_en = start_reg_4; // @[SWChisel.scala 193:22]
  assign r_count_5_clock = clock;
  assign r_count_5_reset = reset;
  assign r_count_5_io_en = start_reg_5; // @[SWChisel.scala 193:22]
  assign r_count_6_clock = clock;
  assign r_count_6_reset = reset;
  assign r_count_6_io_en = start_reg_6; // @[SWChisel.scala 193:22]
  assign r_count_7_clock = clock;
  assign r_count_7_reset = reset;
  assign r_count_7_io_en = start_reg_7; // @[SWChisel.scala 193:22]
  assign r_count_8_clock = clock;
  assign r_count_8_reset = reset;
  assign r_count_8_io_en = start_reg_8; // @[SWChisel.scala 193:22]
  assign r_count_9_clock = clock;
  assign r_count_9_reset = reset;
  assign r_count_9_io_en = start_reg_9; // @[SWChisel.scala 193:22]
  assign max_clock = clock;
  assign max_reset = reset;
  assign max_io_start = start_reg_9; // @[SWChisel.scala 179:16]
  assign max_io_in = V1_10; // @[SWChisel.scala 178:13]
  always @(posedge clock) begin
    if (reset) begin // @[SWChisel.scala 162:18]
      E_0 <= -16'sh2; // @[SWChisel.scala 162:18]
    end else if (start_reg_0) begin // @[SWChisel.scala 208:25]
      E_0 <= array_0_io_e_o; // @[SWChisel.scala 209:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_1 <= -16'sh3; // @[SWChisel.scala 162:18]
    end else if (start_reg_1) begin // @[SWChisel.scala 208:25]
      E_1 <= array_1_io_e_o; // @[SWChisel.scala 209:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_2 <= -16'sh4; // @[SWChisel.scala 162:18]
    end else if (start_reg_2) begin // @[SWChisel.scala 208:25]
      E_2 <= array_2_io_e_o; // @[SWChisel.scala 209:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_3 <= -16'sh5; // @[SWChisel.scala 162:18]
    end else if (start_reg_3) begin // @[SWChisel.scala 208:25]
      E_3 <= array_3_io_e_o; // @[SWChisel.scala 209:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_4 <= -16'sh6; // @[SWChisel.scala 162:18]
    end else if (start_reg_4) begin // @[SWChisel.scala 208:25]
      E_4 <= array_4_io_e_o; // @[SWChisel.scala 209:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_5 <= -16'sh7; // @[SWChisel.scala 162:18]
    end else if (start_reg_5) begin // @[SWChisel.scala 208:25]
      E_5 <= array_5_io_e_o; // @[SWChisel.scala 209:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_6 <= -16'sh8; // @[SWChisel.scala 162:18]
    end else if (start_reg_6) begin // @[SWChisel.scala 208:25]
      E_6 <= array_6_io_e_o; // @[SWChisel.scala 209:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_7 <= -16'sh9; // @[SWChisel.scala 162:18]
    end else if (start_reg_7) begin // @[SWChisel.scala 208:25]
      E_7 <= array_7_io_e_o; // @[SWChisel.scala 209:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_8 <= -16'sha; // @[SWChisel.scala 162:18]
    end else if (start_reg_8) begin // @[SWChisel.scala 208:25]
      E_8 <= array_8_io_e_o; // @[SWChisel.scala 209:12]
    end
    if (reset) begin // @[SWChisel.scala 162:18]
      E_9 <= -16'shb; // @[SWChisel.scala 162:18]
    end else if (start_reg_9) begin // @[SWChisel.scala 208:25]
      E_9 <= array_9_io_e_o; // @[SWChisel.scala 209:12]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_1 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_0) begin // @[SWChisel.scala 208:25]
      F_1 <= array_0_io_f_o; // @[SWChisel.scala 210:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_2 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_1) begin // @[SWChisel.scala 208:25]
      F_2 <= array_1_io_f_o; // @[SWChisel.scala 210:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_3 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_2) begin // @[SWChisel.scala 208:25]
      F_3 <= array_2_io_f_o; // @[SWChisel.scala 210:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_4 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_3) begin // @[SWChisel.scala 208:25]
      F_4 <= array_3_io_f_o; // @[SWChisel.scala 210:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_5 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_4) begin // @[SWChisel.scala 208:25]
      F_5 <= array_4_io_f_o; // @[SWChisel.scala 210:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_6 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_5) begin // @[SWChisel.scala 208:25]
      F_6 <= array_5_io_f_o; // @[SWChisel.scala 210:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_7 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_6) begin // @[SWChisel.scala 208:25]
      F_7 <= array_6_io_f_o; // @[SWChisel.scala 210:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_8 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_7) begin // @[SWChisel.scala 208:25]
      F_8 <= array_7_io_f_o; // @[SWChisel.scala 210:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_9 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_8) begin // @[SWChisel.scala 208:25]
      F_9 <= array_8_io_f_o; // @[SWChisel.scala 210:14]
    end
    if (reset) begin // @[SWChisel.scala 163:18]
      F_10 <= 16'sh0; // @[SWChisel.scala 163:18]
    end else if (start_reg_9) begin // @[SWChisel.scala 208:25]
      F_10 <= array_9_io_f_o; // @[SWChisel.scala 210:14]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_1 <= -16'sh2; // @[SWChisel.scala 164:19]
    end else if (start_reg_0) begin // @[SWChisel.scala 208:25]
      V1_1 <= array_0_io_v_o; // @[SWChisel.scala 211:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_2 <= -16'sh3; // @[SWChisel.scala 164:19]
    end else if (start_reg_1) begin // @[SWChisel.scala 208:25]
      V1_2 <= array_1_io_v_o; // @[SWChisel.scala 211:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_3 <= -16'sh4; // @[SWChisel.scala 164:19]
    end else if (start_reg_2) begin // @[SWChisel.scala 208:25]
      V1_3 <= array_2_io_v_o; // @[SWChisel.scala 211:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_4 <= -16'sh5; // @[SWChisel.scala 164:19]
    end else if (start_reg_3) begin // @[SWChisel.scala 208:25]
      V1_4 <= array_3_io_v_o; // @[SWChisel.scala 211:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_5 <= -16'sh6; // @[SWChisel.scala 164:19]
    end else if (start_reg_4) begin // @[SWChisel.scala 208:25]
      V1_5 <= array_4_io_v_o; // @[SWChisel.scala 211:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_6 <= -16'sh7; // @[SWChisel.scala 164:19]
    end else if (start_reg_5) begin // @[SWChisel.scala 208:25]
      V1_6 <= array_5_io_v_o; // @[SWChisel.scala 211:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_7 <= -16'sh8; // @[SWChisel.scala 164:19]
    end else if (start_reg_6) begin // @[SWChisel.scala 208:25]
      V1_7 <= array_6_io_v_o; // @[SWChisel.scala 211:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_8 <= -16'sh9; // @[SWChisel.scala 164:19]
    end else if (start_reg_7) begin // @[SWChisel.scala 208:25]
      V1_8 <= array_7_io_v_o; // @[SWChisel.scala 211:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_9 <= -16'sha; // @[SWChisel.scala 164:19]
    end else if (start_reg_8) begin // @[SWChisel.scala 208:25]
      V1_9 <= array_8_io_v_o; // @[SWChisel.scala 211:15]
    end
    if (reset) begin // @[SWChisel.scala 164:19]
      V1_10 <= -16'shb; // @[SWChisel.scala 164:19]
    end else if (start_reg_9) begin // @[SWChisel.scala 208:25]
      V1_10 <= array_9_io_v_o; // @[SWChisel.scala 211:15]
    end
    if (reset) begin // @[SWChisel.scala 167:19]
      V2_1 <= 16'sh0; // @[SWChisel.scala 167:19]
    end else begin
      V2_1 <= V1_1; // @[SWChisel.scala 227:11]
    end
    if (reset) begin // @[SWChisel.scala 167:19]
      V2_2 <= 16'sh0; // @[SWChisel.scala 167:19]
    end else begin
      V2_2 <= V1_2; // @[SWChisel.scala 227:11]
    end
    if (reset) begin // @[SWChisel.scala 167:19]
      V2_3 <= 16'sh0; // @[SWChisel.scala 167:19]
    end else begin
      V2_3 <= V1_3; // @[SWChisel.scala 227:11]
    end
    if (reset) begin // @[SWChisel.scala 167:19]
      V2_4 <= 16'sh0; // @[SWChisel.scala 167:19]
    end else begin
      V2_4 <= V1_4; // @[SWChisel.scala 227:11]
    end
    if (reset) begin // @[SWChisel.scala 167:19]
      V2_5 <= 16'sh0; // @[SWChisel.scala 167:19]
    end else begin
      V2_5 <= V1_5; // @[SWChisel.scala 227:11]
    end
    if (reset) begin // @[SWChisel.scala 167:19]
      V2_6 <= 16'sh0; // @[SWChisel.scala 167:19]
    end else begin
      V2_6 <= V1_6; // @[SWChisel.scala 227:11]
    end
    if (reset) begin // @[SWChisel.scala 167:19]
      V2_7 <= 16'sh0; // @[SWChisel.scala 167:19]
    end else begin
      V2_7 <= V1_7; // @[SWChisel.scala 227:11]
    end
    if (reset) begin // @[SWChisel.scala 167:19]
      V2_8 <= 16'sh0; // @[SWChisel.scala 167:19]
    end else begin
      V2_8 <= V1_8; // @[SWChisel.scala 227:11]
    end
    if (reset) begin // @[SWChisel.scala 167:19]
      V2_9 <= 16'sh0; // @[SWChisel.scala 167:19]
    end else begin
      V2_9 <= V1_9; // @[SWChisel.scala 227:11]
    end
    if (reset) begin // @[SWChisel.scala 167:19]
      V2_10 <= 16'sh0; // @[SWChisel.scala 167:19]
    end else begin
      V2_10 <= V1_10; // @[SWChisel.scala 227:11]
    end
    if (reset) begin // @[SWChisel.scala 168:26]
      start_reg_0 <= 1'h0; // @[SWChisel.scala 168:26]
    end else begin
      start_reg_0 <= io_start; // @[SWChisel.scala 186:16]
    end
    if (reset) begin // @[SWChisel.scala 168:26]
      start_reg_1 <= 1'h0; // @[SWChisel.scala 168:26]
    end else begin
      start_reg_1 <= start_reg_0; // @[SWChisel.scala 188:18]
    end
    if (reset) begin // @[SWChisel.scala 168:26]
      start_reg_2 <= 1'h0; // @[SWChisel.scala 168:26]
    end else begin
      start_reg_2 <= start_reg_1; // @[SWChisel.scala 188:18]
    end
    if (reset) begin // @[SWChisel.scala 168:26]
      start_reg_3 <= 1'h0; // @[SWChisel.scala 168:26]
    end else begin
      start_reg_3 <= start_reg_2; // @[SWChisel.scala 188:18]
    end
    if (reset) begin // @[SWChisel.scala 168:26]
      start_reg_4 <= 1'h0; // @[SWChisel.scala 168:26]
    end else begin
      start_reg_4 <= start_reg_3; // @[SWChisel.scala 188:18]
    end
    if (reset) begin // @[SWChisel.scala 168:26]
      start_reg_5 <= 1'h0; // @[SWChisel.scala 168:26]
    end else begin
      start_reg_5 <= start_reg_4; // @[SWChisel.scala 188:18]
    end
    if (reset) begin // @[SWChisel.scala 168:26]
      start_reg_6 <= 1'h0; // @[SWChisel.scala 168:26]
    end else begin
      start_reg_6 <= start_reg_5; // @[SWChisel.scala 188:18]
    end
    if (reset) begin // @[SWChisel.scala 168:26]
      start_reg_7 <= 1'h0; // @[SWChisel.scala 168:26]
    end else begin
      start_reg_7 <= start_reg_6; // @[SWChisel.scala 188:18]
    end
    if (reset) begin // @[SWChisel.scala 168:26]
      start_reg_8 <= 1'h0; // @[SWChisel.scala 168:26]
    end else begin
      start_reg_8 <= start_reg_7; // @[SWChisel.scala 188:18]
    end
    if (reset) begin // @[SWChisel.scala 168:26]
      start_reg_9 <= 1'h0; // @[SWChisel.scala 168:26]
    end else begin
      start_reg_9 <= start_reg_8; // @[SWChisel.scala 188:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  E_0 = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  E_1 = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  E_2 = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  E_3 = _RAND_3[15:0];
  _RAND_4 = {1{`RANDOM}};
  E_4 = _RAND_4[15:0];
  _RAND_5 = {1{`RANDOM}};
  E_5 = _RAND_5[15:0];
  _RAND_6 = {1{`RANDOM}};
  E_6 = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  E_7 = _RAND_7[15:0];
  _RAND_8 = {1{`RANDOM}};
  E_8 = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  E_9 = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  F_1 = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  F_2 = _RAND_11[15:0];
  _RAND_12 = {1{`RANDOM}};
  F_3 = _RAND_12[15:0];
  _RAND_13 = {1{`RANDOM}};
  F_4 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  F_5 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  F_6 = _RAND_15[15:0];
  _RAND_16 = {1{`RANDOM}};
  F_7 = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  F_8 = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  F_9 = _RAND_18[15:0];
  _RAND_19 = {1{`RANDOM}};
  F_10 = _RAND_19[15:0];
  _RAND_20 = {1{`RANDOM}};
  V1_1 = _RAND_20[15:0];
  _RAND_21 = {1{`RANDOM}};
  V1_2 = _RAND_21[15:0];
  _RAND_22 = {1{`RANDOM}};
  V1_3 = _RAND_22[15:0];
  _RAND_23 = {1{`RANDOM}};
  V1_4 = _RAND_23[15:0];
  _RAND_24 = {1{`RANDOM}};
  V1_5 = _RAND_24[15:0];
  _RAND_25 = {1{`RANDOM}};
  V1_6 = _RAND_25[15:0];
  _RAND_26 = {1{`RANDOM}};
  V1_7 = _RAND_26[15:0];
  _RAND_27 = {1{`RANDOM}};
  V1_8 = _RAND_27[15:0];
  _RAND_28 = {1{`RANDOM}};
  V1_9 = _RAND_28[15:0];
  _RAND_29 = {1{`RANDOM}};
  V1_10 = _RAND_29[15:0];
  _RAND_30 = {1{`RANDOM}};
  V2_1 = _RAND_30[15:0];
  _RAND_31 = {1{`RANDOM}};
  V2_2 = _RAND_31[15:0];
  _RAND_32 = {1{`RANDOM}};
  V2_3 = _RAND_32[15:0];
  _RAND_33 = {1{`RANDOM}};
  V2_4 = _RAND_33[15:0];
  _RAND_34 = {1{`RANDOM}};
  V2_5 = _RAND_34[15:0];
  _RAND_35 = {1{`RANDOM}};
  V2_6 = _RAND_35[15:0];
  _RAND_36 = {1{`RANDOM}};
  V2_7 = _RAND_36[15:0];
  _RAND_37 = {1{`RANDOM}};
  V2_8 = _RAND_37[15:0];
  _RAND_38 = {1{`RANDOM}};
  V2_9 = _RAND_38[15:0];
  _RAND_39 = {1{`RANDOM}};
  V2_10 = _RAND_39[15:0];
  _RAND_40 = {1{`RANDOM}};
  start_reg_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  start_reg_1 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  start_reg_2 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  start_reg_3 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  start_reg_4 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  start_reg_5 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  start_reg_6 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  start_reg_7 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  start_reg_8 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  start_reg_9 = _RAND_49[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
